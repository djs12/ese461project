
module Top ( clk, reset, inputSramWe, pixels, weight1, w2SramWeOffChip, 
        weight2, weight2AddrOffChip, weight2_loadNextRow, rdata );
  input [89:0] pixels;
  input [8:0] weight1;
  input [15:0] weight2;
  input [3:0] weight2AddrOffChip;
  output [15:0] rdata;
  input clk, reset, inputSramWe, w2SramWeOffChip;
  output weight2_loadNextRow;
  wire   \sig_in[15] , \INPUTSRAM/mem_i[9][8] , \INPUTSRAM/mem_i[9][7] ,
         \INPUTSRAM/mem_i[9][6] , \INPUTSRAM/mem_i[9][5] ,
         \INPUTSRAM/mem_i[9][4] , \INPUTSRAM/mem_i[9][3] ,
         \INPUTSRAM/mem_i[9][2] , \INPUTSRAM/mem_i[9][1] ,
         \INPUTSRAM/mem_i[9][0] , \INPUTSRAM/mem_i[8][8] ,
         \INPUTSRAM/mem_i[8][7] , \INPUTSRAM/mem_i[8][6] ,
         \INPUTSRAM/mem_i[8][5] , \INPUTSRAM/mem_i[8][4] ,
         \INPUTSRAM/mem_i[8][3] , \INPUTSRAM/mem_i[8][2] ,
         \INPUTSRAM/mem_i[8][1] , \INPUTSRAM/mem_i[8][0] ,
         \INPUTSRAM/mem_i[7][8] , \INPUTSRAM/mem_i[7][7] ,
         \INPUTSRAM/mem_i[7][6] , \INPUTSRAM/mem_i[7][5] ,
         \INPUTSRAM/mem_i[7][4] , \INPUTSRAM/mem_i[7][3] ,
         \INPUTSRAM/mem_i[7][2] , \INPUTSRAM/mem_i[7][1] ,
         \INPUTSRAM/mem_i[7][0] , \INPUTSRAM/mem_i[6][8] ,
         \INPUTSRAM/mem_i[6][7] , \INPUTSRAM/mem_i[6][6] ,
         \INPUTSRAM/mem_i[6][5] , \INPUTSRAM/mem_i[6][4] ,
         \INPUTSRAM/mem_i[6][3] , \INPUTSRAM/mem_i[6][2] ,
         \INPUTSRAM/mem_i[6][1] , \INPUTSRAM/mem_i[6][0] ,
         \INPUTSRAM/mem_i[5][8] , \INPUTSRAM/mem_i[5][7] ,
         \INPUTSRAM/mem_i[5][6] , \INPUTSRAM/mem_i[5][5] ,
         \INPUTSRAM/mem_i[5][4] , \INPUTSRAM/mem_i[5][3] ,
         \INPUTSRAM/mem_i[5][2] , \INPUTSRAM/mem_i[5][1] ,
         \INPUTSRAM/mem_i[5][0] , \INPUTSRAM/mem_i[4][8] ,
         \INPUTSRAM/mem_i[4][7] , \INPUTSRAM/mem_i[4][6] ,
         \INPUTSRAM/mem_i[4][5] , \INPUTSRAM/mem_i[4][4] ,
         \INPUTSRAM/mem_i[4][3] , \INPUTSRAM/mem_i[4][2] ,
         \INPUTSRAM/mem_i[4][1] , \INPUTSRAM/mem_i[4][0] ,
         \INPUTSRAM/mem_i[3][8] , \INPUTSRAM/mem_i[3][7] ,
         \INPUTSRAM/mem_i[3][6] , \INPUTSRAM/mem_i[3][5] ,
         \INPUTSRAM/mem_i[3][4] , \INPUTSRAM/mem_i[3][3] ,
         \INPUTSRAM/mem_i[3][2] , \INPUTSRAM/mem_i[3][1] ,
         \INPUTSRAM/mem_i[3][0] , \INPUTSRAM/mem_i[2][8] ,
         \INPUTSRAM/mem_i[2][7] , \INPUTSRAM/mem_i[2][6] ,
         \INPUTSRAM/mem_i[2][5] , \INPUTSRAM/mem_i[2][4] ,
         \INPUTSRAM/mem_i[2][3] , \INPUTSRAM/mem_i[2][2] ,
         \INPUTSRAM/mem_i[2][1] , \INPUTSRAM/mem_i[2][0] ,
         \INPUTSRAM/mem_i[1][8] , \INPUTSRAM/mem_i[1][7] ,
         \INPUTSRAM/mem_i[1][6] , \INPUTSRAM/mem_i[1][5] ,
         \INPUTSRAM/mem_i[1][4] , \INPUTSRAM/mem_i[1][3] ,
         \INPUTSRAM/mem_i[1][2] , \INPUTSRAM/mem_i[1][1] ,
         \INPUTSRAM/mem_i[1][0] , \INPUTSRAM/mem_i[0][8] ,
         \INPUTSRAM/mem_i[0][7] , \INPUTSRAM/mem_i[0][6] ,
         \INPUTSRAM/mem_i[0][5] , \INPUTSRAM/mem_i[0][4] ,
         \INPUTSRAM/mem_i[0][3] , \INPUTSRAM/mem_i[0][2] ,
         \INPUTSRAM/mem_i[0][1] , \INPUTSRAM/mem_i[0][0] , \CNTRL/N242 ,
         \CNTRL/N241 , \CNTRL/N240 , \CNTRL/N239 , \CNTRL/N238 , \CNTRL/N237 ,
         \CNTRL/N236 , \CNTRL/N235 , \CNTRL/N234 , \CNTRL/N233 ,
         \WEIGHT_2/mem_w2[9][15] , \WEIGHT_2/mem_w2[9][14] ,
         \WEIGHT_2/mem_w2[9][13] , \WEIGHT_2/mem_w2[9][12] ,
         \WEIGHT_2/mem_w2[9][11] , \WEIGHT_2/mem_w2[9][10] ,
         \WEIGHT_2/mem_w2[9][9] , \WEIGHT_2/mem_w2[9][8] ,
         \WEIGHT_2/mem_w2[9][7] , \WEIGHT_2/mem_w2[9][6] ,
         \WEIGHT_2/mem_w2[9][5] , \WEIGHT_2/mem_w2[9][4] ,
         \WEIGHT_2/mem_w2[9][3] , \WEIGHT_2/mem_w2[9][2] ,
         \WEIGHT_2/mem_w2[9][1] , \WEIGHT_2/mem_w2[9][0] ,
         \WEIGHT_2/mem_w2[8][15] , \WEIGHT_2/mem_w2[8][14] ,
         \WEIGHT_2/mem_w2[8][13] , \WEIGHT_2/mem_w2[8][12] ,
         \WEIGHT_2/mem_w2[8][11] , \WEIGHT_2/mem_w2[8][10] ,
         \WEIGHT_2/mem_w2[8][9] , \WEIGHT_2/mem_w2[8][8] ,
         \WEIGHT_2/mem_w2[8][7] , \WEIGHT_2/mem_w2[8][6] ,
         \WEIGHT_2/mem_w2[8][5] , \WEIGHT_2/mem_w2[8][4] ,
         \WEIGHT_2/mem_w2[8][3] , \WEIGHT_2/mem_w2[8][2] ,
         \WEIGHT_2/mem_w2[8][1] , \WEIGHT_2/mem_w2[8][0] ,
         \WEIGHT_2/mem_w2[7][15] , \WEIGHT_2/mem_w2[7][14] ,
         \WEIGHT_2/mem_w2[7][13] , \WEIGHT_2/mem_w2[7][12] ,
         \WEIGHT_2/mem_w2[7][11] , \WEIGHT_2/mem_w2[7][10] ,
         \WEIGHT_2/mem_w2[7][9] , \WEIGHT_2/mem_w2[7][8] ,
         \WEIGHT_2/mem_w2[7][7] , \WEIGHT_2/mem_w2[7][6] ,
         \WEIGHT_2/mem_w2[7][5] , \WEIGHT_2/mem_w2[7][4] ,
         \WEIGHT_2/mem_w2[7][3] , \WEIGHT_2/mem_w2[7][2] ,
         \WEIGHT_2/mem_w2[7][1] , \WEIGHT_2/mem_w2[7][0] ,
         \WEIGHT_2/mem_w2[6][15] , \WEIGHT_2/mem_w2[6][14] ,
         \WEIGHT_2/mem_w2[6][13] , \WEIGHT_2/mem_w2[6][12] ,
         \WEIGHT_2/mem_w2[6][11] , \WEIGHT_2/mem_w2[6][10] ,
         \WEIGHT_2/mem_w2[6][9] , \WEIGHT_2/mem_w2[6][8] ,
         \WEIGHT_2/mem_w2[6][7] , \WEIGHT_2/mem_w2[6][6] ,
         \WEIGHT_2/mem_w2[6][5] , \WEIGHT_2/mem_w2[6][4] ,
         \WEIGHT_2/mem_w2[6][3] , \WEIGHT_2/mem_w2[6][2] ,
         \WEIGHT_2/mem_w2[6][1] , \WEIGHT_2/mem_w2[6][0] ,
         \WEIGHT_2/mem_w2[5][15] , \WEIGHT_2/mem_w2[5][14] ,
         \WEIGHT_2/mem_w2[5][13] , \WEIGHT_2/mem_w2[5][12] ,
         \WEIGHT_2/mem_w2[5][11] , \WEIGHT_2/mem_w2[5][10] ,
         \WEIGHT_2/mem_w2[5][9] , \WEIGHT_2/mem_w2[5][8] ,
         \WEIGHT_2/mem_w2[5][7] , \WEIGHT_2/mem_w2[5][6] ,
         \WEIGHT_2/mem_w2[5][5] , \WEIGHT_2/mem_w2[5][4] ,
         \WEIGHT_2/mem_w2[5][3] , \WEIGHT_2/mem_w2[5][2] ,
         \WEIGHT_2/mem_w2[5][1] , \WEIGHT_2/mem_w2[5][0] ,
         \WEIGHT_2/mem_w2[4][15] , \WEIGHT_2/mem_w2[4][14] ,
         \WEIGHT_2/mem_w2[4][13] , \WEIGHT_2/mem_w2[4][12] ,
         \WEIGHT_2/mem_w2[4][11] , \WEIGHT_2/mem_w2[4][10] ,
         \WEIGHT_2/mem_w2[4][9] , \WEIGHT_2/mem_w2[4][8] ,
         \WEIGHT_2/mem_w2[4][7] , \WEIGHT_2/mem_w2[4][6] ,
         \WEIGHT_2/mem_w2[4][5] , \WEIGHT_2/mem_w2[4][4] ,
         \WEIGHT_2/mem_w2[4][3] , \WEIGHT_2/mem_w2[4][2] ,
         \WEIGHT_2/mem_w2[4][1] , \WEIGHT_2/mem_w2[4][0] ,
         \WEIGHT_2/mem_w2[3][15] , \WEIGHT_2/mem_w2[3][14] ,
         \WEIGHT_2/mem_w2[3][13] , \WEIGHT_2/mem_w2[3][12] ,
         \WEIGHT_2/mem_w2[3][11] , \WEIGHT_2/mem_w2[3][10] ,
         \WEIGHT_2/mem_w2[3][9] , \WEIGHT_2/mem_w2[3][8] ,
         \WEIGHT_2/mem_w2[3][7] , \WEIGHT_2/mem_w2[3][6] ,
         \WEIGHT_2/mem_w2[3][5] , \WEIGHT_2/mem_w2[3][4] ,
         \WEIGHT_2/mem_w2[3][3] , \WEIGHT_2/mem_w2[3][2] ,
         \WEIGHT_2/mem_w2[3][1] , \WEIGHT_2/mem_w2[3][0] ,
         \WEIGHT_2/mem_w2[2][15] , \WEIGHT_2/mem_w2[2][14] ,
         \WEIGHT_2/mem_w2[2][13] , \WEIGHT_2/mem_w2[2][12] ,
         \WEIGHT_2/mem_w2[2][11] , \WEIGHT_2/mem_w2[2][10] ,
         \WEIGHT_2/mem_w2[2][9] , \WEIGHT_2/mem_w2[2][8] ,
         \WEIGHT_2/mem_w2[2][7] , \WEIGHT_2/mem_w2[2][6] ,
         \WEIGHT_2/mem_w2[2][5] , \WEIGHT_2/mem_w2[2][4] ,
         \WEIGHT_2/mem_w2[2][3] , \WEIGHT_2/mem_w2[2][2] ,
         \WEIGHT_2/mem_w2[2][1] , \WEIGHT_2/mem_w2[2][0] ,
         \WEIGHT_2/mem_w2[1][15] , \WEIGHT_2/mem_w2[1][14] ,
         \WEIGHT_2/mem_w2[1][13] , \WEIGHT_2/mem_w2[1][12] ,
         \WEIGHT_2/mem_w2[1][11] , \WEIGHT_2/mem_w2[1][10] ,
         \WEIGHT_2/mem_w2[1][9] , \WEIGHT_2/mem_w2[1][8] ,
         \WEIGHT_2/mem_w2[1][7] , \WEIGHT_2/mem_w2[1][6] ,
         \WEIGHT_2/mem_w2[1][5] , \WEIGHT_2/mem_w2[1][4] ,
         \WEIGHT_2/mem_w2[1][3] , \WEIGHT_2/mem_w2[1][2] ,
         \WEIGHT_2/mem_w2[1][1] , \WEIGHT_2/mem_w2[1][0] ,
         \WEIGHT_2/mem_w2[0][15] , \WEIGHT_2/mem_w2[0][14] ,
         \WEIGHT_2/mem_w2[0][13] , \WEIGHT_2/mem_w2[0][12] ,
         \WEIGHT_2/mem_w2[0][11] , \WEIGHT_2/mem_w2[0][10] ,
         \WEIGHT_2/mem_w2[0][9] , \WEIGHT_2/mem_w2[0][8] ,
         \WEIGHT_2/mem_w2[0][7] , \WEIGHT_2/mem_w2[0][6] ,
         \WEIGHT_2/mem_w2[0][5] , \WEIGHT_2/mem_w2[0][4] ,
         \WEIGHT_2/mem_w2[0][3] , \WEIGHT_2/mem_w2[0][2] ,
         \WEIGHT_2/mem_w2[0][1] , \WEIGHT_2/mem_w2[0][0] , \ANSWER/N487 ,
         \ANSWER/N486 , \ANSWER/N485 , \ANSWER/N484 , \ANSWER/N483 ,
         \ANSWER/N482 , \ANSWER/N481 , \ANSWER/N480 , \ANSWER/N479 ,
         \ANSWER/N478 , \ANSWER/N477 , \ANSWER/N476 , \ANSWER/N475 ,
         \ANSWER/N474 , \ANSWER/N473 , \ANSWER/N472 , \ANSWER/mem[9][9][15] ,
         \ANSWER/mem[9][9][14] , \ANSWER/mem[9][9][13] ,
         \ANSWER/mem[9][9][12] , \ANSWER/mem[9][9][11] ,
         \ANSWER/mem[9][9][10] , \ANSWER/mem[9][9][9] , \ANSWER/mem[9][9][8] ,
         \ANSWER/mem[9][9][7] , \ANSWER/mem[9][9][6] , \ANSWER/mem[9][9][5] ,
         \ANSWER/mem[9][9][4] , \ANSWER/mem[9][9][3] , \ANSWER/mem[9][9][2] ,
         \ANSWER/mem[9][9][1] , \ANSWER/mem[9][9][0] , \ANSWER/mem[9][8][15] ,
         \ANSWER/mem[9][8][14] , \ANSWER/mem[9][8][13] ,
         \ANSWER/mem[9][8][12] , \ANSWER/mem[9][8][11] ,
         \ANSWER/mem[9][8][10] , \ANSWER/mem[9][8][9] , \ANSWER/mem[9][8][8] ,
         \ANSWER/mem[9][8][7] , \ANSWER/mem[9][8][6] , \ANSWER/mem[9][8][5] ,
         \ANSWER/mem[9][8][4] , \ANSWER/mem[9][8][3] , \ANSWER/mem[9][8][2] ,
         \ANSWER/mem[9][8][1] , \ANSWER/mem[9][8][0] , \ANSWER/mem[9][7][15] ,
         \ANSWER/mem[9][7][14] , \ANSWER/mem[9][7][13] ,
         \ANSWER/mem[9][7][12] , \ANSWER/mem[9][7][11] ,
         \ANSWER/mem[9][7][10] , \ANSWER/mem[9][7][9] , \ANSWER/mem[9][7][8] ,
         \ANSWER/mem[9][7][7] , \ANSWER/mem[9][7][6] , \ANSWER/mem[9][7][5] ,
         \ANSWER/mem[9][7][4] , \ANSWER/mem[9][7][3] , \ANSWER/mem[9][7][2] ,
         \ANSWER/mem[9][7][1] , \ANSWER/mem[9][7][0] , \ANSWER/mem[9][6][15] ,
         \ANSWER/mem[9][6][14] , \ANSWER/mem[9][6][13] ,
         \ANSWER/mem[9][6][12] , \ANSWER/mem[9][6][11] ,
         \ANSWER/mem[9][6][10] , \ANSWER/mem[9][6][9] , \ANSWER/mem[9][6][8] ,
         \ANSWER/mem[9][6][7] , \ANSWER/mem[9][6][6] , \ANSWER/mem[9][6][5] ,
         \ANSWER/mem[9][6][4] , \ANSWER/mem[9][6][3] , \ANSWER/mem[9][6][2] ,
         \ANSWER/mem[9][6][1] , \ANSWER/mem[9][6][0] , \ANSWER/mem[9][5][15] ,
         \ANSWER/mem[9][5][14] , \ANSWER/mem[9][5][13] ,
         \ANSWER/mem[9][5][12] , \ANSWER/mem[9][5][11] ,
         \ANSWER/mem[9][5][10] , \ANSWER/mem[9][5][9] , \ANSWER/mem[9][5][8] ,
         \ANSWER/mem[9][5][7] , \ANSWER/mem[9][5][6] , \ANSWER/mem[9][5][5] ,
         \ANSWER/mem[9][5][4] , \ANSWER/mem[9][5][3] , \ANSWER/mem[9][5][2] ,
         \ANSWER/mem[9][5][1] , \ANSWER/mem[9][5][0] , \ANSWER/mem[9][4][15] ,
         \ANSWER/mem[9][4][14] , \ANSWER/mem[9][4][13] ,
         \ANSWER/mem[9][4][12] , \ANSWER/mem[9][4][11] ,
         \ANSWER/mem[9][4][10] , \ANSWER/mem[9][4][9] , \ANSWER/mem[9][4][8] ,
         \ANSWER/mem[9][4][7] , \ANSWER/mem[9][4][6] , \ANSWER/mem[9][4][5] ,
         \ANSWER/mem[9][4][4] , \ANSWER/mem[9][4][3] , \ANSWER/mem[9][4][2] ,
         \ANSWER/mem[9][4][1] , \ANSWER/mem[9][4][0] , \ANSWER/mem[9][3][15] ,
         \ANSWER/mem[9][3][14] , \ANSWER/mem[9][3][13] ,
         \ANSWER/mem[9][3][12] , \ANSWER/mem[9][3][11] ,
         \ANSWER/mem[9][3][10] , \ANSWER/mem[9][3][9] , \ANSWER/mem[9][3][8] ,
         \ANSWER/mem[9][3][7] , \ANSWER/mem[9][3][6] , \ANSWER/mem[9][3][5] ,
         \ANSWER/mem[9][3][4] , \ANSWER/mem[9][3][3] , \ANSWER/mem[9][3][2] ,
         \ANSWER/mem[9][3][1] , \ANSWER/mem[9][3][0] , \ANSWER/mem[9][2][15] ,
         \ANSWER/mem[9][2][14] , \ANSWER/mem[9][2][13] ,
         \ANSWER/mem[9][2][12] , \ANSWER/mem[9][2][11] ,
         \ANSWER/mem[9][2][10] , \ANSWER/mem[9][2][9] , \ANSWER/mem[9][2][8] ,
         \ANSWER/mem[9][2][7] , \ANSWER/mem[9][2][6] , \ANSWER/mem[9][2][5] ,
         \ANSWER/mem[9][2][4] , \ANSWER/mem[9][2][3] , \ANSWER/mem[9][2][2] ,
         \ANSWER/mem[9][2][1] , \ANSWER/mem[9][2][0] , \ANSWER/mem[9][1][15] ,
         \ANSWER/mem[9][1][14] , \ANSWER/mem[9][1][13] ,
         \ANSWER/mem[9][1][12] , \ANSWER/mem[9][1][11] ,
         \ANSWER/mem[9][1][10] , \ANSWER/mem[9][1][9] , \ANSWER/mem[9][1][8] ,
         \ANSWER/mem[9][1][7] , \ANSWER/mem[9][1][6] , \ANSWER/mem[9][1][5] ,
         \ANSWER/mem[9][1][4] , \ANSWER/mem[9][1][3] , \ANSWER/mem[9][1][2] ,
         \ANSWER/mem[9][1][1] , \ANSWER/mem[9][1][0] , \ANSWER/mem[9][0][15] ,
         \ANSWER/mem[9][0][14] , \ANSWER/mem[9][0][13] ,
         \ANSWER/mem[9][0][12] , \ANSWER/mem[9][0][11] ,
         \ANSWER/mem[9][0][10] , \ANSWER/mem[9][0][9] , \ANSWER/mem[9][0][8] ,
         \ANSWER/mem[9][0][7] , \ANSWER/mem[9][0][6] , \ANSWER/mem[9][0][5] ,
         \ANSWER/mem[9][0][4] , \ANSWER/mem[9][0][3] , \ANSWER/mem[9][0][2] ,
         \ANSWER/mem[9][0][1] , \ANSWER/mem[9][0][0] , \ANSWER/mem[8][9][15] ,
         \ANSWER/mem[8][9][14] , \ANSWER/mem[8][9][13] ,
         \ANSWER/mem[8][9][12] , \ANSWER/mem[8][9][11] ,
         \ANSWER/mem[8][9][10] , \ANSWER/mem[8][9][9] , \ANSWER/mem[8][9][8] ,
         \ANSWER/mem[8][9][7] , \ANSWER/mem[8][9][6] , \ANSWER/mem[8][9][5] ,
         \ANSWER/mem[8][9][4] , \ANSWER/mem[8][9][3] , \ANSWER/mem[8][9][2] ,
         \ANSWER/mem[8][9][1] , \ANSWER/mem[8][9][0] , \ANSWER/mem[8][8][15] ,
         \ANSWER/mem[8][8][14] , \ANSWER/mem[8][8][13] ,
         \ANSWER/mem[8][8][12] , \ANSWER/mem[8][8][11] ,
         \ANSWER/mem[8][8][10] , \ANSWER/mem[8][8][9] , \ANSWER/mem[8][8][8] ,
         \ANSWER/mem[8][8][7] , \ANSWER/mem[8][8][6] , \ANSWER/mem[8][8][5] ,
         \ANSWER/mem[8][8][4] , \ANSWER/mem[8][8][3] , \ANSWER/mem[8][8][2] ,
         \ANSWER/mem[8][8][1] , \ANSWER/mem[8][8][0] , \ANSWER/mem[8][7][15] ,
         \ANSWER/mem[8][7][14] , \ANSWER/mem[8][7][13] ,
         \ANSWER/mem[8][7][12] , \ANSWER/mem[8][7][11] ,
         \ANSWER/mem[8][7][10] , \ANSWER/mem[8][7][9] , \ANSWER/mem[8][7][8] ,
         \ANSWER/mem[8][7][7] , \ANSWER/mem[8][7][6] , \ANSWER/mem[8][7][5] ,
         \ANSWER/mem[8][7][4] , \ANSWER/mem[8][7][3] , \ANSWER/mem[8][7][2] ,
         \ANSWER/mem[8][7][1] , \ANSWER/mem[8][7][0] , \ANSWER/mem[8][6][15] ,
         \ANSWER/mem[8][6][14] , \ANSWER/mem[8][6][13] ,
         \ANSWER/mem[8][6][12] , \ANSWER/mem[8][6][11] ,
         \ANSWER/mem[8][6][10] , \ANSWER/mem[8][6][9] , \ANSWER/mem[8][6][8] ,
         \ANSWER/mem[8][6][7] , \ANSWER/mem[8][6][6] , \ANSWER/mem[8][6][5] ,
         \ANSWER/mem[8][6][4] , \ANSWER/mem[8][6][3] , \ANSWER/mem[8][6][2] ,
         \ANSWER/mem[8][6][1] , \ANSWER/mem[8][6][0] , \ANSWER/mem[8][5][15] ,
         \ANSWER/mem[8][5][14] , \ANSWER/mem[8][5][13] ,
         \ANSWER/mem[8][5][12] , \ANSWER/mem[8][5][11] ,
         \ANSWER/mem[8][5][10] , \ANSWER/mem[8][5][9] , \ANSWER/mem[8][5][8] ,
         \ANSWER/mem[8][5][7] , \ANSWER/mem[8][5][6] , \ANSWER/mem[8][5][5] ,
         \ANSWER/mem[8][5][4] , \ANSWER/mem[8][5][3] , \ANSWER/mem[8][5][2] ,
         \ANSWER/mem[8][5][1] , \ANSWER/mem[8][5][0] , \ANSWER/mem[8][4][15] ,
         \ANSWER/mem[8][4][14] , \ANSWER/mem[8][4][13] ,
         \ANSWER/mem[8][4][12] , \ANSWER/mem[8][4][11] ,
         \ANSWER/mem[8][4][10] , \ANSWER/mem[8][4][9] , \ANSWER/mem[8][4][8] ,
         \ANSWER/mem[8][4][7] , \ANSWER/mem[8][4][6] , \ANSWER/mem[8][4][5] ,
         \ANSWER/mem[8][4][4] , \ANSWER/mem[8][4][3] , \ANSWER/mem[8][4][2] ,
         \ANSWER/mem[8][4][1] , \ANSWER/mem[8][4][0] , \ANSWER/mem[8][3][15] ,
         \ANSWER/mem[8][3][14] , \ANSWER/mem[8][3][13] ,
         \ANSWER/mem[8][3][12] , \ANSWER/mem[8][3][11] ,
         \ANSWER/mem[8][3][10] , \ANSWER/mem[8][3][9] , \ANSWER/mem[8][3][8] ,
         \ANSWER/mem[8][3][7] , \ANSWER/mem[8][3][6] , \ANSWER/mem[8][3][5] ,
         \ANSWER/mem[8][3][4] , \ANSWER/mem[8][3][3] , \ANSWER/mem[8][3][2] ,
         \ANSWER/mem[8][3][1] , \ANSWER/mem[8][3][0] , \ANSWER/mem[8][2][15] ,
         \ANSWER/mem[8][2][14] , \ANSWER/mem[8][2][13] ,
         \ANSWER/mem[8][2][12] , \ANSWER/mem[8][2][11] ,
         \ANSWER/mem[8][2][10] , \ANSWER/mem[8][2][9] , \ANSWER/mem[8][2][8] ,
         \ANSWER/mem[8][2][7] , \ANSWER/mem[8][2][6] , \ANSWER/mem[8][2][5] ,
         \ANSWER/mem[8][2][4] , \ANSWER/mem[8][2][3] , \ANSWER/mem[8][2][2] ,
         \ANSWER/mem[8][2][1] , \ANSWER/mem[8][2][0] , \ANSWER/mem[8][1][15] ,
         \ANSWER/mem[8][1][14] , \ANSWER/mem[8][1][13] ,
         \ANSWER/mem[8][1][12] , \ANSWER/mem[8][1][11] ,
         \ANSWER/mem[8][1][10] , \ANSWER/mem[8][1][9] , \ANSWER/mem[8][1][8] ,
         \ANSWER/mem[8][1][7] , \ANSWER/mem[8][1][6] , \ANSWER/mem[8][1][5] ,
         \ANSWER/mem[8][1][4] , \ANSWER/mem[8][1][3] , \ANSWER/mem[8][1][2] ,
         \ANSWER/mem[8][1][1] , \ANSWER/mem[8][1][0] , \ANSWER/mem[8][0][15] ,
         \ANSWER/mem[8][0][14] , \ANSWER/mem[8][0][13] ,
         \ANSWER/mem[8][0][12] , \ANSWER/mem[8][0][11] ,
         \ANSWER/mem[8][0][10] , \ANSWER/mem[8][0][9] , \ANSWER/mem[8][0][8] ,
         \ANSWER/mem[8][0][7] , \ANSWER/mem[8][0][6] , \ANSWER/mem[8][0][5] ,
         \ANSWER/mem[8][0][4] , \ANSWER/mem[8][0][3] , \ANSWER/mem[8][0][2] ,
         \ANSWER/mem[8][0][1] , \ANSWER/mem[8][0][0] , \ANSWER/mem[7][9][15] ,
         \ANSWER/mem[7][9][14] , \ANSWER/mem[7][9][13] ,
         \ANSWER/mem[7][9][12] , \ANSWER/mem[7][9][11] ,
         \ANSWER/mem[7][9][10] , \ANSWER/mem[7][9][9] , \ANSWER/mem[7][9][8] ,
         \ANSWER/mem[7][9][7] , \ANSWER/mem[7][9][6] , \ANSWER/mem[7][9][5] ,
         \ANSWER/mem[7][9][4] , \ANSWER/mem[7][9][3] , \ANSWER/mem[7][9][2] ,
         \ANSWER/mem[7][9][1] , \ANSWER/mem[7][9][0] , \ANSWER/mem[7][8][15] ,
         \ANSWER/mem[7][8][14] , \ANSWER/mem[7][8][13] ,
         \ANSWER/mem[7][8][12] , \ANSWER/mem[7][8][11] ,
         \ANSWER/mem[7][8][10] , \ANSWER/mem[7][8][9] , \ANSWER/mem[7][8][8] ,
         \ANSWER/mem[7][8][7] , \ANSWER/mem[7][8][6] , \ANSWER/mem[7][8][5] ,
         \ANSWER/mem[7][8][4] , \ANSWER/mem[7][8][3] , \ANSWER/mem[7][8][2] ,
         \ANSWER/mem[7][8][1] , \ANSWER/mem[7][8][0] , \ANSWER/mem[7][7][15] ,
         \ANSWER/mem[7][7][14] , \ANSWER/mem[7][7][13] ,
         \ANSWER/mem[7][7][12] , \ANSWER/mem[7][7][11] ,
         \ANSWER/mem[7][7][10] , \ANSWER/mem[7][7][9] , \ANSWER/mem[7][7][8] ,
         \ANSWER/mem[7][7][7] , \ANSWER/mem[7][7][6] , \ANSWER/mem[7][7][5] ,
         \ANSWER/mem[7][7][4] , \ANSWER/mem[7][7][3] , \ANSWER/mem[7][7][2] ,
         \ANSWER/mem[7][7][1] , \ANSWER/mem[7][7][0] , \ANSWER/mem[7][6][15] ,
         \ANSWER/mem[7][6][14] , \ANSWER/mem[7][6][13] ,
         \ANSWER/mem[7][6][12] , \ANSWER/mem[7][6][11] ,
         \ANSWER/mem[7][6][10] , \ANSWER/mem[7][6][9] , \ANSWER/mem[7][6][8] ,
         \ANSWER/mem[7][6][7] , \ANSWER/mem[7][6][6] , \ANSWER/mem[7][6][5] ,
         \ANSWER/mem[7][6][4] , \ANSWER/mem[7][6][3] , \ANSWER/mem[7][6][2] ,
         \ANSWER/mem[7][6][1] , \ANSWER/mem[7][6][0] , \ANSWER/mem[7][5][15] ,
         \ANSWER/mem[7][5][14] , \ANSWER/mem[7][5][13] ,
         \ANSWER/mem[7][5][12] , \ANSWER/mem[7][5][11] ,
         \ANSWER/mem[7][5][10] , \ANSWER/mem[7][5][9] , \ANSWER/mem[7][5][8] ,
         \ANSWER/mem[7][5][7] , \ANSWER/mem[7][5][6] , \ANSWER/mem[7][5][5] ,
         \ANSWER/mem[7][5][4] , \ANSWER/mem[7][5][3] , \ANSWER/mem[7][5][2] ,
         \ANSWER/mem[7][5][1] , \ANSWER/mem[7][5][0] , \ANSWER/mem[7][4][15] ,
         \ANSWER/mem[7][4][14] , \ANSWER/mem[7][4][13] ,
         \ANSWER/mem[7][4][12] , \ANSWER/mem[7][4][11] ,
         \ANSWER/mem[7][4][10] , \ANSWER/mem[7][4][9] , \ANSWER/mem[7][4][8] ,
         \ANSWER/mem[7][4][7] , \ANSWER/mem[7][4][6] , \ANSWER/mem[7][4][5] ,
         \ANSWER/mem[7][4][4] , \ANSWER/mem[7][4][3] , \ANSWER/mem[7][4][2] ,
         \ANSWER/mem[7][4][1] , \ANSWER/mem[7][4][0] , \ANSWER/mem[7][3][15] ,
         \ANSWER/mem[7][3][14] , \ANSWER/mem[7][3][13] ,
         \ANSWER/mem[7][3][12] , \ANSWER/mem[7][3][11] ,
         \ANSWER/mem[7][3][10] , \ANSWER/mem[7][3][9] , \ANSWER/mem[7][3][8] ,
         \ANSWER/mem[7][3][7] , \ANSWER/mem[7][3][6] , \ANSWER/mem[7][3][5] ,
         \ANSWER/mem[7][3][4] , \ANSWER/mem[7][3][3] , \ANSWER/mem[7][3][2] ,
         \ANSWER/mem[7][3][1] , \ANSWER/mem[7][3][0] , \ANSWER/mem[7][2][15] ,
         \ANSWER/mem[7][2][14] , \ANSWER/mem[7][2][13] ,
         \ANSWER/mem[7][2][12] , \ANSWER/mem[7][2][11] ,
         \ANSWER/mem[7][2][10] , \ANSWER/mem[7][2][9] , \ANSWER/mem[7][2][8] ,
         \ANSWER/mem[7][2][7] , \ANSWER/mem[7][2][6] , \ANSWER/mem[7][2][5] ,
         \ANSWER/mem[7][2][4] , \ANSWER/mem[7][2][3] , \ANSWER/mem[7][2][2] ,
         \ANSWER/mem[7][2][1] , \ANSWER/mem[7][2][0] , \ANSWER/mem[7][1][15] ,
         \ANSWER/mem[7][1][14] , \ANSWER/mem[7][1][13] ,
         \ANSWER/mem[7][1][12] , \ANSWER/mem[7][1][11] ,
         \ANSWER/mem[7][1][10] , \ANSWER/mem[7][1][9] , \ANSWER/mem[7][1][8] ,
         \ANSWER/mem[7][1][7] , \ANSWER/mem[7][1][6] , \ANSWER/mem[7][1][5] ,
         \ANSWER/mem[7][1][4] , \ANSWER/mem[7][1][3] , \ANSWER/mem[7][1][2] ,
         \ANSWER/mem[7][1][1] , \ANSWER/mem[7][1][0] , \ANSWER/mem[7][0][15] ,
         \ANSWER/mem[7][0][14] , \ANSWER/mem[7][0][13] ,
         \ANSWER/mem[7][0][12] , \ANSWER/mem[7][0][11] ,
         \ANSWER/mem[7][0][10] , \ANSWER/mem[7][0][9] , \ANSWER/mem[7][0][8] ,
         \ANSWER/mem[7][0][7] , \ANSWER/mem[7][0][6] , \ANSWER/mem[7][0][5] ,
         \ANSWER/mem[7][0][4] , \ANSWER/mem[7][0][3] , \ANSWER/mem[7][0][2] ,
         \ANSWER/mem[7][0][1] , \ANSWER/mem[7][0][0] , \ANSWER/mem[6][9][15] ,
         \ANSWER/mem[6][9][14] , \ANSWER/mem[6][9][13] ,
         \ANSWER/mem[6][9][12] , \ANSWER/mem[6][9][11] ,
         \ANSWER/mem[6][9][10] , \ANSWER/mem[6][9][9] , \ANSWER/mem[6][9][8] ,
         \ANSWER/mem[6][9][7] , \ANSWER/mem[6][9][6] , \ANSWER/mem[6][9][5] ,
         \ANSWER/mem[6][9][4] , \ANSWER/mem[6][9][3] , \ANSWER/mem[6][9][2] ,
         \ANSWER/mem[6][9][1] , \ANSWER/mem[6][9][0] , \ANSWER/mem[6][8][15] ,
         \ANSWER/mem[6][8][14] , \ANSWER/mem[6][8][13] ,
         \ANSWER/mem[6][8][12] , \ANSWER/mem[6][8][11] ,
         \ANSWER/mem[6][8][10] , \ANSWER/mem[6][8][9] , \ANSWER/mem[6][8][8] ,
         \ANSWER/mem[6][8][7] , \ANSWER/mem[6][8][6] , \ANSWER/mem[6][8][5] ,
         \ANSWER/mem[6][8][4] , \ANSWER/mem[6][8][3] , \ANSWER/mem[6][8][2] ,
         \ANSWER/mem[6][8][1] , \ANSWER/mem[6][8][0] , \ANSWER/mem[6][7][15] ,
         \ANSWER/mem[6][7][14] , \ANSWER/mem[6][7][13] ,
         \ANSWER/mem[6][7][12] , \ANSWER/mem[6][7][11] ,
         \ANSWER/mem[6][7][10] , \ANSWER/mem[6][7][9] , \ANSWER/mem[6][7][8] ,
         \ANSWER/mem[6][7][7] , \ANSWER/mem[6][7][6] , \ANSWER/mem[6][7][5] ,
         \ANSWER/mem[6][7][4] , \ANSWER/mem[6][7][3] , \ANSWER/mem[6][7][2] ,
         \ANSWER/mem[6][7][1] , \ANSWER/mem[6][7][0] , \ANSWER/mem[6][6][15] ,
         \ANSWER/mem[6][6][14] , \ANSWER/mem[6][6][13] ,
         \ANSWER/mem[6][6][12] , \ANSWER/mem[6][6][11] ,
         \ANSWER/mem[6][6][10] , \ANSWER/mem[6][6][9] , \ANSWER/mem[6][6][8] ,
         \ANSWER/mem[6][6][7] , \ANSWER/mem[6][6][6] , \ANSWER/mem[6][6][5] ,
         \ANSWER/mem[6][6][4] , \ANSWER/mem[6][6][3] , \ANSWER/mem[6][6][2] ,
         \ANSWER/mem[6][6][1] , \ANSWER/mem[6][6][0] , \ANSWER/mem[6][5][15] ,
         \ANSWER/mem[6][5][14] , \ANSWER/mem[6][5][13] ,
         \ANSWER/mem[6][5][12] , \ANSWER/mem[6][5][11] ,
         \ANSWER/mem[6][5][10] , \ANSWER/mem[6][5][9] , \ANSWER/mem[6][5][8] ,
         \ANSWER/mem[6][5][7] , \ANSWER/mem[6][5][6] , \ANSWER/mem[6][5][5] ,
         \ANSWER/mem[6][5][4] , \ANSWER/mem[6][5][3] , \ANSWER/mem[6][5][2] ,
         \ANSWER/mem[6][5][1] , \ANSWER/mem[6][5][0] , \ANSWER/mem[6][4][15] ,
         \ANSWER/mem[6][4][14] , \ANSWER/mem[6][4][13] ,
         \ANSWER/mem[6][4][12] , \ANSWER/mem[6][4][11] ,
         \ANSWER/mem[6][4][10] , \ANSWER/mem[6][4][9] , \ANSWER/mem[6][4][8] ,
         \ANSWER/mem[6][4][7] , \ANSWER/mem[6][4][6] , \ANSWER/mem[6][4][5] ,
         \ANSWER/mem[6][4][4] , \ANSWER/mem[6][4][3] , \ANSWER/mem[6][4][2] ,
         \ANSWER/mem[6][4][1] , \ANSWER/mem[6][4][0] , \ANSWER/mem[6][3][15] ,
         \ANSWER/mem[6][3][14] , \ANSWER/mem[6][3][13] ,
         \ANSWER/mem[6][3][12] , \ANSWER/mem[6][3][11] ,
         \ANSWER/mem[6][3][10] , \ANSWER/mem[6][3][9] , \ANSWER/mem[6][3][8] ,
         \ANSWER/mem[6][3][7] , \ANSWER/mem[6][3][6] , \ANSWER/mem[6][3][5] ,
         \ANSWER/mem[6][3][4] , \ANSWER/mem[6][3][3] , \ANSWER/mem[6][3][2] ,
         \ANSWER/mem[6][3][1] , \ANSWER/mem[6][3][0] , \ANSWER/mem[6][2][15] ,
         \ANSWER/mem[6][2][14] , \ANSWER/mem[6][2][13] ,
         \ANSWER/mem[6][2][12] , \ANSWER/mem[6][2][11] ,
         \ANSWER/mem[6][2][10] , \ANSWER/mem[6][2][9] , \ANSWER/mem[6][2][8] ,
         \ANSWER/mem[6][2][7] , \ANSWER/mem[6][2][6] , \ANSWER/mem[6][2][5] ,
         \ANSWER/mem[6][2][4] , \ANSWER/mem[6][2][3] , \ANSWER/mem[6][2][2] ,
         \ANSWER/mem[6][2][1] , \ANSWER/mem[6][2][0] , \ANSWER/mem[6][1][15] ,
         \ANSWER/mem[6][1][14] , \ANSWER/mem[6][1][13] ,
         \ANSWER/mem[6][1][12] , \ANSWER/mem[6][1][11] ,
         \ANSWER/mem[6][1][10] , \ANSWER/mem[6][1][9] , \ANSWER/mem[6][1][8] ,
         \ANSWER/mem[6][1][7] , \ANSWER/mem[6][1][6] , \ANSWER/mem[6][1][5] ,
         \ANSWER/mem[6][1][4] , \ANSWER/mem[6][1][3] , \ANSWER/mem[6][1][2] ,
         \ANSWER/mem[6][1][1] , \ANSWER/mem[6][1][0] , \ANSWER/mem[6][0][15] ,
         \ANSWER/mem[6][0][14] , \ANSWER/mem[6][0][13] ,
         \ANSWER/mem[6][0][12] , \ANSWER/mem[6][0][11] ,
         \ANSWER/mem[6][0][10] , \ANSWER/mem[6][0][9] , \ANSWER/mem[6][0][8] ,
         \ANSWER/mem[6][0][7] , \ANSWER/mem[6][0][6] , \ANSWER/mem[6][0][5] ,
         \ANSWER/mem[6][0][4] , \ANSWER/mem[6][0][3] , \ANSWER/mem[6][0][2] ,
         \ANSWER/mem[6][0][1] , \ANSWER/mem[6][0][0] , \ANSWER/mem[5][9][15] ,
         \ANSWER/mem[5][9][14] , \ANSWER/mem[5][9][13] ,
         \ANSWER/mem[5][9][12] , \ANSWER/mem[5][9][11] ,
         \ANSWER/mem[5][9][10] , \ANSWER/mem[5][9][9] , \ANSWER/mem[5][9][8] ,
         \ANSWER/mem[5][9][7] , \ANSWER/mem[5][9][6] , \ANSWER/mem[5][9][5] ,
         \ANSWER/mem[5][9][4] , \ANSWER/mem[5][9][3] , \ANSWER/mem[5][9][2] ,
         \ANSWER/mem[5][9][1] , \ANSWER/mem[5][9][0] , \ANSWER/mem[5][8][15] ,
         \ANSWER/mem[5][8][14] , \ANSWER/mem[5][8][13] ,
         \ANSWER/mem[5][8][12] , \ANSWER/mem[5][8][11] ,
         \ANSWER/mem[5][8][10] , \ANSWER/mem[5][8][9] , \ANSWER/mem[5][8][8] ,
         \ANSWER/mem[5][8][7] , \ANSWER/mem[5][8][6] , \ANSWER/mem[5][8][5] ,
         \ANSWER/mem[5][8][4] , \ANSWER/mem[5][8][3] , \ANSWER/mem[5][8][2] ,
         \ANSWER/mem[5][8][1] , \ANSWER/mem[5][8][0] , \ANSWER/mem[5][7][15] ,
         \ANSWER/mem[5][7][14] , \ANSWER/mem[5][7][13] ,
         \ANSWER/mem[5][7][12] , \ANSWER/mem[5][7][11] ,
         \ANSWER/mem[5][7][10] , \ANSWER/mem[5][7][9] , \ANSWER/mem[5][7][8] ,
         \ANSWER/mem[5][7][7] , \ANSWER/mem[5][7][6] , \ANSWER/mem[5][7][5] ,
         \ANSWER/mem[5][7][4] , \ANSWER/mem[5][7][3] , \ANSWER/mem[5][7][2] ,
         \ANSWER/mem[5][7][1] , \ANSWER/mem[5][7][0] , \ANSWER/mem[5][6][15] ,
         \ANSWER/mem[5][6][14] , \ANSWER/mem[5][6][13] ,
         \ANSWER/mem[5][6][12] , \ANSWER/mem[5][6][11] ,
         \ANSWER/mem[5][6][10] , \ANSWER/mem[5][6][9] , \ANSWER/mem[5][6][8] ,
         \ANSWER/mem[5][6][7] , \ANSWER/mem[5][6][6] , \ANSWER/mem[5][6][5] ,
         \ANSWER/mem[5][6][4] , \ANSWER/mem[5][6][3] , \ANSWER/mem[5][6][2] ,
         \ANSWER/mem[5][6][1] , \ANSWER/mem[5][6][0] , \ANSWER/mem[5][5][15] ,
         \ANSWER/mem[5][5][14] , \ANSWER/mem[5][5][13] ,
         \ANSWER/mem[5][5][12] , \ANSWER/mem[5][5][11] ,
         \ANSWER/mem[5][5][10] , \ANSWER/mem[5][5][9] , \ANSWER/mem[5][5][8] ,
         \ANSWER/mem[5][5][7] , \ANSWER/mem[5][5][6] , \ANSWER/mem[5][5][5] ,
         \ANSWER/mem[5][5][4] , \ANSWER/mem[5][5][3] , \ANSWER/mem[5][5][2] ,
         \ANSWER/mem[5][5][1] , \ANSWER/mem[5][5][0] , \ANSWER/mem[5][4][15] ,
         \ANSWER/mem[5][4][14] , \ANSWER/mem[5][4][13] ,
         \ANSWER/mem[5][4][12] , \ANSWER/mem[5][4][11] ,
         \ANSWER/mem[5][4][10] , \ANSWER/mem[5][4][9] , \ANSWER/mem[5][4][8] ,
         \ANSWER/mem[5][4][7] , \ANSWER/mem[5][4][6] , \ANSWER/mem[5][4][5] ,
         \ANSWER/mem[5][4][4] , \ANSWER/mem[5][4][3] , \ANSWER/mem[5][4][2] ,
         \ANSWER/mem[5][4][1] , \ANSWER/mem[5][4][0] , \ANSWER/mem[5][3][15] ,
         \ANSWER/mem[5][3][14] , \ANSWER/mem[5][3][13] ,
         \ANSWER/mem[5][3][12] , \ANSWER/mem[5][3][11] ,
         \ANSWER/mem[5][3][10] , \ANSWER/mem[5][3][9] , \ANSWER/mem[5][3][8] ,
         \ANSWER/mem[5][3][7] , \ANSWER/mem[5][3][6] , \ANSWER/mem[5][3][5] ,
         \ANSWER/mem[5][3][4] , \ANSWER/mem[5][3][3] , \ANSWER/mem[5][3][2] ,
         \ANSWER/mem[5][3][1] , \ANSWER/mem[5][3][0] , \ANSWER/mem[5][2][15] ,
         \ANSWER/mem[5][2][14] , \ANSWER/mem[5][2][13] ,
         \ANSWER/mem[5][2][12] , \ANSWER/mem[5][2][11] ,
         \ANSWER/mem[5][2][10] , \ANSWER/mem[5][2][9] , \ANSWER/mem[5][2][8] ,
         \ANSWER/mem[5][2][7] , \ANSWER/mem[5][2][6] , \ANSWER/mem[5][2][5] ,
         \ANSWER/mem[5][2][4] , \ANSWER/mem[5][2][3] , \ANSWER/mem[5][2][2] ,
         \ANSWER/mem[5][2][1] , \ANSWER/mem[5][2][0] , \ANSWER/mem[5][1][15] ,
         \ANSWER/mem[5][1][14] , \ANSWER/mem[5][1][13] ,
         \ANSWER/mem[5][1][12] , \ANSWER/mem[5][1][11] ,
         \ANSWER/mem[5][1][10] , \ANSWER/mem[5][1][9] , \ANSWER/mem[5][1][8] ,
         \ANSWER/mem[5][1][7] , \ANSWER/mem[5][1][6] , \ANSWER/mem[5][1][5] ,
         \ANSWER/mem[5][1][4] , \ANSWER/mem[5][1][3] , \ANSWER/mem[5][1][2] ,
         \ANSWER/mem[5][1][1] , \ANSWER/mem[5][1][0] , \ANSWER/mem[5][0][15] ,
         \ANSWER/mem[5][0][14] , \ANSWER/mem[5][0][13] ,
         \ANSWER/mem[5][0][12] , \ANSWER/mem[5][0][11] ,
         \ANSWER/mem[5][0][10] , \ANSWER/mem[5][0][9] , \ANSWER/mem[5][0][8] ,
         \ANSWER/mem[5][0][7] , \ANSWER/mem[5][0][6] , \ANSWER/mem[5][0][5] ,
         \ANSWER/mem[5][0][4] , \ANSWER/mem[5][0][3] , \ANSWER/mem[5][0][2] ,
         \ANSWER/mem[5][0][1] , \ANSWER/mem[5][0][0] , \ANSWER/mem[4][9][15] ,
         \ANSWER/mem[4][9][14] , \ANSWER/mem[4][9][13] ,
         \ANSWER/mem[4][9][12] , \ANSWER/mem[4][9][11] ,
         \ANSWER/mem[4][9][10] , \ANSWER/mem[4][9][9] , \ANSWER/mem[4][9][8] ,
         \ANSWER/mem[4][9][7] , \ANSWER/mem[4][9][6] , \ANSWER/mem[4][9][5] ,
         \ANSWER/mem[4][9][4] , \ANSWER/mem[4][9][3] , \ANSWER/mem[4][9][2] ,
         \ANSWER/mem[4][9][1] , \ANSWER/mem[4][9][0] , \ANSWER/mem[4][8][15] ,
         \ANSWER/mem[4][8][14] , \ANSWER/mem[4][8][13] ,
         \ANSWER/mem[4][8][12] , \ANSWER/mem[4][8][11] ,
         \ANSWER/mem[4][8][10] , \ANSWER/mem[4][8][9] , \ANSWER/mem[4][8][8] ,
         \ANSWER/mem[4][8][7] , \ANSWER/mem[4][8][6] , \ANSWER/mem[4][8][5] ,
         \ANSWER/mem[4][8][4] , \ANSWER/mem[4][8][3] , \ANSWER/mem[4][8][2] ,
         \ANSWER/mem[4][8][1] , \ANSWER/mem[4][8][0] , \ANSWER/mem[4][7][15] ,
         \ANSWER/mem[4][7][14] , \ANSWER/mem[4][7][13] ,
         \ANSWER/mem[4][7][12] , \ANSWER/mem[4][7][11] ,
         \ANSWER/mem[4][7][10] , \ANSWER/mem[4][7][9] , \ANSWER/mem[4][7][8] ,
         \ANSWER/mem[4][7][7] , \ANSWER/mem[4][7][6] , \ANSWER/mem[4][7][5] ,
         \ANSWER/mem[4][7][4] , \ANSWER/mem[4][7][3] , \ANSWER/mem[4][7][2] ,
         \ANSWER/mem[4][7][1] , \ANSWER/mem[4][7][0] , \ANSWER/mem[4][6][15] ,
         \ANSWER/mem[4][6][14] , \ANSWER/mem[4][6][13] ,
         \ANSWER/mem[4][6][12] , \ANSWER/mem[4][6][11] ,
         \ANSWER/mem[4][6][10] , \ANSWER/mem[4][6][9] , \ANSWER/mem[4][6][8] ,
         \ANSWER/mem[4][6][7] , \ANSWER/mem[4][6][6] , \ANSWER/mem[4][6][5] ,
         \ANSWER/mem[4][6][4] , \ANSWER/mem[4][6][3] , \ANSWER/mem[4][6][2] ,
         \ANSWER/mem[4][6][1] , \ANSWER/mem[4][6][0] , \ANSWER/mem[4][5][15] ,
         \ANSWER/mem[4][5][14] , \ANSWER/mem[4][5][13] ,
         \ANSWER/mem[4][5][12] , \ANSWER/mem[4][5][11] ,
         \ANSWER/mem[4][5][10] , \ANSWER/mem[4][5][9] , \ANSWER/mem[4][5][8] ,
         \ANSWER/mem[4][5][7] , \ANSWER/mem[4][5][6] , \ANSWER/mem[4][5][5] ,
         \ANSWER/mem[4][5][4] , \ANSWER/mem[4][5][3] , \ANSWER/mem[4][5][2] ,
         \ANSWER/mem[4][5][1] , \ANSWER/mem[4][5][0] , \ANSWER/mem[4][4][15] ,
         \ANSWER/mem[4][4][14] , \ANSWER/mem[4][4][13] ,
         \ANSWER/mem[4][4][12] , \ANSWER/mem[4][4][11] ,
         \ANSWER/mem[4][4][10] , \ANSWER/mem[4][4][9] , \ANSWER/mem[4][4][8] ,
         \ANSWER/mem[4][4][7] , \ANSWER/mem[4][4][6] , \ANSWER/mem[4][4][5] ,
         \ANSWER/mem[4][4][4] , \ANSWER/mem[4][4][3] , \ANSWER/mem[4][4][2] ,
         \ANSWER/mem[4][4][1] , \ANSWER/mem[4][4][0] , \ANSWER/mem[4][3][15] ,
         \ANSWER/mem[4][3][14] , \ANSWER/mem[4][3][13] ,
         \ANSWER/mem[4][3][12] , \ANSWER/mem[4][3][11] ,
         \ANSWER/mem[4][3][10] , \ANSWER/mem[4][3][9] , \ANSWER/mem[4][3][8] ,
         \ANSWER/mem[4][3][7] , \ANSWER/mem[4][3][6] , \ANSWER/mem[4][3][5] ,
         \ANSWER/mem[4][3][4] , \ANSWER/mem[4][3][3] , \ANSWER/mem[4][3][2] ,
         \ANSWER/mem[4][3][1] , \ANSWER/mem[4][3][0] , \ANSWER/mem[4][2][15] ,
         \ANSWER/mem[4][2][14] , \ANSWER/mem[4][2][13] ,
         \ANSWER/mem[4][2][12] , \ANSWER/mem[4][2][11] ,
         \ANSWER/mem[4][2][10] , \ANSWER/mem[4][2][9] , \ANSWER/mem[4][2][8] ,
         \ANSWER/mem[4][2][7] , \ANSWER/mem[4][2][6] , \ANSWER/mem[4][2][5] ,
         \ANSWER/mem[4][2][4] , \ANSWER/mem[4][2][3] , \ANSWER/mem[4][2][2] ,
         \ANSWER/mem[4][2][1] , \ANSWER/mem[4][2][0] , \ANSWER/mem[4][1][15] ,
         \ANSWER/mem[4][1][14] , \ANSWER/mem[4][1][13] ,
         \ANSWER/mem[4][1][12] , \ANSWER/mem[4][1][11] ,
         \ANSWER/mem[4][1][10] , \ANSWER/mem[4][1][9] , \ANSWER/mem[4][1][8] ,
         \ANSWER/mem[4][1][7] , \ANSWER/mem[4][1][6] , \ANSWER/mem[4][1][5] ,
         \ANSWER/mem[4][1][4] , \ANSWER/mem[4][1][3] , \ANSWER/mem[4][1][2] ,
         \ANSWER/mem[4][1][1] , \ANSWER/mem[4][1][0] , \ANSWER/mem[4][0][15] ,
         \ANSWER/mem[4][0][14] , \ANSWER/mem[4][0][13] ,
         \ANSWER/mem[4][0][12] , \ANSWER/mem[4][0][11] ,
         \ANSWER/mem[4][0][10] , \ANSWER/mem[4][0][9] , \ANSWER/mem[4][0][8] ,
         \ANSWER/mem[4][0][7] , \ANSWER/mem[4][0][6] , \ANSWER/mem[4][0][5] ,
         \ANSWER/mem[4][0][4] , \ANSWER/mem[4][0][3] , \ANSWER/mem[4][0][2] ,
         \ANSWER/mem[4][0][1] , \ANSWER/mem[4][0][0] , \ANSWER/mem[3][9][15] ,
         \ANSWER/mem[3][9][14] , \ANSWER/mem[3][9][13] ,
         \ANSWER/mem[3][9][12] , \ANSWER/mem[3][9][11] ,
         \ANSWER/mem[3][9][10] , \ANSWER/mem[3][9][9] , \ANSWER/mem[3][9][8] ,
         \ANSWER/mem[3][9][7] , \ANSWER/mem[3][9][6] , \ANSWER/mem[3][9][5] ,
         \ANSWER/mem[3][9][4] , \ANSWER/mem[3][9][3] , \ANSWER/mem[3][9][2] ,
         \ANSWER/mem[3][9][1] , \ANSWER/mem[3][9][0] , \ANSWER/mem[3][8][15] ,
         \ANSWER/mem[3][8][14] , \ANSWER/mem[3][8][13] ,
         \ANSWER/mem[3][8][12] , \ANSWER/mem[3][8][11] ,
         \ANSWER/mem[3][8][10] , \ANSWER/mem[3][8][9] , \ANSWER/mem[3][8][8] ,
         \ANSWER/mem[3][8][7] , \ANSWER/mem[3][8][6] , \ANSWER/mem[3][8][5] ,
         \ANSWER/mem[3][8][4] , \ANSWER/mem[3][8][3] , \ANSWER/mem[3][8][2] ,
         \ANSWER/mem[3][8][1] , \ANSWER/mem[3][8][0] , \ANSWER/mem[3][7][15] ,
         \ANSWER/mem[3][7][14] , \ANSWER/mem[3][7][13] ,
         \ANSWER/mem[3][7][12] , \ANSWER/mem[3][7][11] ,
         \ANSWER/mem[3][7][10] , \ANSWER/mem[3][7][9] , \ANSWER/mem[3][7][8] ,
         \ANSWER/mem[3][7][7] , \ANSWER/mem[3][7][6] , \ANSWER/mem[3][7][5] ,
         \ANSWER/mem[3][7][4] , \ANSWER/mem[3][7][3] , \ANSWER/mem[3][7][2] ,
         \ANSWER/mem[3][7][1] , \ANSWER/mem[3][7][0] , \ANSWER/mem[3][6][15] ,
         \ANSWER/mem[3][6][14] , \ANSWER/mem[3][6][13] ,
         \ANSWER/mem[3][6][12] , \ANSWER/mem[3][6][11] ,
         \ANSWER/mem[3][6][10] , \ANSWER/mem[3][6][9] , \ANSWER/mem[3][6][8] ,
         \ANSWER/mem[3][6][7] , \ANSWER/mem[3][6][6] , \ANSWER/mem[3][6][5] ,
         \ANSWER/mem[3][6][4] , \ANSWER/mem[3][6][3] , \ANSWER/mem[3][6][2] ,
         \ANSWER/mem[3][6][1] , \ANSWER/mem[3][6][0] , \ANSWER/mem[3][5][15] ,
         \ANSWER/mem[3][5][14] , \ANSWER/mem[3][5][13] ,
         \ANSWER/mem[3][5][12] , \ANSWER/mem[3][5][11] ,
         \ANSWER/mem[3][5][10] , \ANSWER/mem[3][5][9] , \ANSWER/mem[3][5][8] ,
         \ANSWER/mem[3][5][7] , \ANSWER/mem[3][5][6] , \ANSWER/mem[3][5][5] ,
         \ANSWER/mem[3][5][4] , \ANSWER/mem[3][5][3] , \ANSWER/mem[3][5][2] ,
         \ANSWER/mem[3][5][1] , \ANSWER/mem[3][5][0] , \ANSWER/mem[3][4][15] ,
         \ANSWER/mem[3][4][14] , \ANSWER/mem[3][4][13] ,
         \ANSWER/mem[3][4][12] , \ANSWER/mem[3][4][11] ,
         \ANSWER/mem[3][4][10] , \ANSWER/mem[3][4][9] , \ANSWER/mem[3][4][8] ,
         \ANSWER/mem[3][4][7] , \ANSWER/mem[3][4][6] , \ANSWER/mem[3][4][5] ,
         \ANSWER/mem[3][4][4] , \ANSWER/mem[3][4][3] , \ANSWER/mem[3][4][2] ,
         \ANSWER/mem[3][4][1] , \ANSWER/mem[3][4][0] , \ANSWER/mem[3][3][15] ,
         \ANSWER/mem[3][3][14] , \ANSWER/mem[3][3][13] ,
         \ANSWER/mem[3][3][12] , \ANSWER/mem[3][3][11] ,
         \ANSWER/mem[3][3][10] , \ANSWER/mem[3][3][9] , \ANSWER/mem[3][3][8] ,
         \ANSWER/mem[3][3][7] , \ANSWER/mem[3][3][6] , \ANSWER/mem[3][3][5] ,
         \ANSWER/mem[3][3][4] , \ANSWER/mem[3][3][3] , \ANSWER/mem[3][3][2] ,
         \ANSWER/mem[3][3][1] , \ANSWER/mem[3][3][0] , \ANSWER/mem[3][2][15] ,
         \ANSWER/mem[3][2][14] , \ANSWER/mem[3][2][13] ,
         \ANSWER/mem[3][2][12] , \ANSWER/mem[3][2][11] ,
         \ANSWER/mem[3][2][10] , \ANSWER/mem[3][2][9] , \ANSWER/mem[3][2][8] ,
         \ANSWER/mem[3][2][7] , \ANSWER/mem[3][2][6] , \ANSWER/mem[3][2][5] ,
         \ANSWER/mem[3][2][4] , \ANSWER/mem[3][2][3] , \ANSWER/mem[3][2][2] ,
         \ANSWER/mem[3][2][1] , \ANSWER/mem[3][2][0] , \ANSWER/mem[3][1][15] ,
         \ANSWER/mem[3][1][14] , \ANSWER/mem[3][1][13] ,
         \ANSWER/mem[3][1][12] , \ANSWER/mem[3][1][11] ,
         \ANSWER/mem[3][1][10] , \ANSWER/mem[3][1][9] , \ANSWER/mem[3][1][8] ,
         \ANSWER/mem[3][1][7] , \ANSWER/mem[3][1][6] , \ANSWER/mem[3][1][5] ,
         \ANSWER/mem[3][1][4] , \ANSWER/mem[3][1][3] , \ANSWER/mem[3][1][2] ,
         \ANSWER/mem[3][1][1] , \ANSWER/mem[3][1][0] , \ANSWER/mem[3][0][15] ,
         \ANSWER/mem[3][0][14] , \ANSWER/mem[3][0][13] ,
         \ANSWER/mem[3][0][12] , \ANSWER/mem[3][0][11] ,
         \ANSWER/mem[3][0][10] , \ANSWER/mem[3][0][9] , \ANSWER/mem[3][0][8] ,
         \ANSWER/mem[3][0][7] , \ANSWER/mem[3][0][6] , \ANSWER/mem[3][0][5] ,
         \ANSWER/mem[3][0][4] , \ANSWER/mem[3][0][3] , \ANSWER/mem[3][0][2] ,
         \ANSWER/mem[3][0][1] , \ANSWER/mem[3][0][0] , \ANSWER/mem[2][9][15] ,
         \ANSWER/mem[2][9][14] , \ANSWER/mem[2][9][13] ,
         \ANSWER/mem[2][9][12] , \ANSWER/mem[2][9][11] ,
         \ANSWER/mem[2][9][10] , \ANSWER/mem[2][9][9] , \ANSWER/mem[2][9][8] ,
         \ANSWER/mem[2][9][7] , \ANSWER/mem[2][9][6] , \ANSWER/mem[2][9][5] ,
         \ANSWER/mem[2][9][4] , \ANSWER/mem[2][9][3] , \ANSWER/mem[2][9][2] ,
         \ANSWER/mem[2][9][1] , \ANSWER/mem[2][9][0] , \ANSWER/mem[2][8][15] ,
         \ANSWER/mem[2][8][14] , \ANSWER/mem[2][8][13] ,
         \ANSWER/mem[2][8][12] , \ANSWER/mem[2][8][11] ,
         \ANSWER/mem[2][8][10] , \ANSWER/mem[2][8][9] , \ANSWER/mem[2][8][8] ,
         \ANSWER/mem[2][8][7] , \ANSWER/mem[2][8][6] , \ANSWER/mem[2][8][5] ,
         \ANSWER/mem[2][8][4] , \ANSWER/mem[2][8][3] , \ANSWER/mem[2][8][2] ,
         \ANSWER/mem[2][8][1] , \ANSWER/mem[2][8][0] , \ANSWER/mem[2][7][15] ,
         \ANSWER/mem[2][7][14] , \ANSWER/mem[2][7][13] ,
         \ANSWER/mem[2][7][12] , \ANSWER/mem[2][7][11] ,
         \ANSWER/mem[2][7][10] , \ANSWER/mem[2][7][9] , \ANSWER/mem[2][7][8] ,
         \ANSWER/mem[2][7][7] , \ANSWER/mem[2][7][6] , \ANSWER/mem[2][7][5] ,
         \ANSWER/mem[2][7][4] , \ANSWER/mem[2][7][3] , \ANSWER/mem[2][7][2] ,
         \ANSWER/mem[2][7][1] , \ANSWER/mem[2][7][0] , \ANSWER/mem[2][6][15] ,
         \ANSWER/mem[2][6][14] , \ANSWER/mem[2][6][13] ,
         \ANSWER/mem[2][6][12] , \ANSWER/mem[2][6][11] ,
         \ANSWER/mem[2][6][10] , \ANSWER/mem[2][6][9] , \ANSWER/mem[2][6][8] ,
         \ANSWER/mem[2][6][7] , \ANSWER/mem[2][6][6] , \ANSWER/mem[2][6][5] ,
         \ANSWER/mem[2][6][4] , \ANSWER/mem[2][6][3] , \ANSWER/mem[2][6][2] ,
         \ANSWER/mem[2][6][1] , \ANSWER/mem[2][6][0] , \ANSWER/mem[2][5][15] ,
         \ANSWER/mem[2][5][14] , \ANSWER/mem[2][5][13] ,
         \ANSWER/mem[2][5][12] , \ANSWER/mem[2][5][11] ,
         \ANSWER/mem[2][5][10] , \ANSWER/mem[2][5][9] , \ANSWER/mem[2][5][8] ,
         \ANSWER/mem[2][5][7] , \ANSWER/mem[2][5][6] , \ANSWER/mem[2][5][5] ,
         \ANSWER/mem[2][5][4] , \ANSWER/mem[2][5][3] , \ANSWER/mem[2][5][2] ,
         \ANSWER/mem[2][5][1] , \ANSWER/mem[2][5][0] , \ANSWER/mem[2][4][15] ,
         \ANSWER/mem[2][4][14] , \ANSWER/mem[2][4][13] ,
         \ANSWER/mem[2][4][12] , \ANSWER/mem[2][4][11] ,
         \ANSWER/mem[2][4][10] , \ANSWER/mem[2][4][9] , \ANSWER/mem[2][4][8] ,
         \ANSWER/mem[2][4][7] , \ANSWER/mem[2][4][6] , \ANSWER/mem[2][4][5] ,
         \ANSWER/mem[2][4][4] , \ANSWER/mem[2][4][3] , \ANSWER/mem[2][4][2] ,
         \ANSWER/mem[2][4][1] , \ANSWER/mem[2][4][0] , \ANSWER/mem[2][3][15] ,
         \ANSWER/mem[2][3][14] , \ANSWER/mem[2][3][13] ,
         \ANSWER/mem[2][3][12] , \ANSWER/mem[2][3][11] ,
         \ANSWER/mem[2][3][10] , \ANSWER/mem[2][3][9] , \ANSWER/mem[2][3][8] ,
         \ANSWER/mem[2][3][7] , \ANSWER/mem[2][3][6] , \ANSWER/mem[2][3][5] ,
         \ANSWER/mem[2][3][4] , \ANSWER/mem[2][3][3] , \ANSWER/mem[2][3][2] ,
         \ANSWER/mem[2][3][1] , \ANSWER/mem[2][3][0] , \ANSWER/mem[2][2][15] ,
         \ANSWER/mem[2][2][14] , \ANSWER/mem[2][2][13] ,
         \ANSWER/mem[2][2][12] , \ANSWER/mem[2][2][11] ,
         \ANSWER/mem[2][2][10] , \ANSWER/mem[2][2][9] , \ANSWER/mem[2][2][8] ,
         \ANSWER/mem[2][2][7] , \ANSWER/mem[2][2][6] , \ANSWER/mem[2][2][5] ,
         \ANSWER/mem[2][2][4] , \ANSWER/mem[2][2][3] , \ANSWER/mem[2][2][2] ,
         \ANSWER/mem[2][2][1] , \ANSWER/mem[2][2][0] , \ANSWER/mem[2][1][15] ,
         \ANSWER/mem[2][1][14] , \ANSWER/mem[2][1][13] ,
         \ANSWER/mem[2][1][12] , \ANSWER/mem[2][1][11] ,
         \ANSWER/mem[2][1][10] , \ANSWER/mem[2][1][9] , \ANSWER/mem[2][1][8] ,
         \ANSWER/mem[2][1][7] , \ANSWER/mem[2][1][6] , \ANSWER/mem[2][1][5] ,
         \ANSWER/mem[2][1][4] , \ANSWER/mem[2][1][3] , \ANSWER/mem[2][1][2] ,
         \ANSWER/mem[2][1][1] , \ANSWER/mem[2][1][0] , \ANSWER/mem[2][0][15] ,
         \ANSWER/mem[2][0][14] , \ANSWER/mem[2][0][13] ,
         \ANSWER/mem[2][0][12] , \ANSWER/mem[2][0][11] ,
         \ANSWER/mem[2][0][10] , \ANSWER/mem[2][0][9] , \ANSWER/mem[2][0][8] ,
         \ANSWER/mem[2][0][7] , \ANSWER/mem[2][0][6] , \ANSWER/mem[2][0][5] ,
         \ANSWER/mem[2][0][4] , \ANSWER/mem[2][0][3] , \ANSWER/mem[2][0][2] ,
         \ANSWER/mem[2][0][1] , \ANSWER/mem[2][0][0] , \ANSWER/mem[1][9][15] ,
         \ANSWER/mem[1][9][14] , \ANSWER/mem[1][9][13] ,
         \ANSWER/mem[1][9][12] , \ANSWER/mem[1][9][11] ,
         \ANSWER/mem[1][9][10] , \ANSWER/mem[1][9][9] , \ANSWER/mem[1][9][8] ,
         \ANSWER/mem[1][9][7] , \ANSWER/mem[1][9][6] , \ANSWER/mem[1][9][5] ,
         \ANSWER/mem[1][9][4] , \ANSWER/mem[1][9][3] , \ANSWER/mem[1][9][2] ,
         \ANSWER/mem[1][9][1] , \ANSWER/mem[1][9][0] , \ANSWER/mem[1][8][15] ,
         \ANSWER/mem[1][8][14] , \ANSWER/mem[1][8][13] ,
         \ANSWER/mem[1][8][12] , \ANSWER/mem[1][8][11] ,
         \ANSWER/mem[1][8][10] , \ANSWER/mem[1][8][9] , \ANSWER/mem[1][8][8] ,
         \ANSWER/mem[1][8][7] , \ANSWER/mem[1][8][6] , \ANSWER/mem[1][8][5] ,
         \ANSWER/mem[1][8][4] , \ANSWER/mem[1][8][3] , \ANSWER/mem[1][8][2] ,
         \ANSWER/mem[1][8][1] , \ANSWER/mem[1][8][0] , \ANSWER/mem[1][7][15] ,
         \ANSWER/mem[1][7][14] , \ANSWER/mem[1][7][13] ,
         \ANSWER/mem[1][7][12] , \ANSWER/mem[1][7][11] ,
         \ANSWER/mem[1][7][10] , \ANSWER/mem[1][7][9] , \ANSWER/mem[1][7][8] ,
         \ANSWER/mem[1][7][7] , \ANSWER/mem[1][7][6] , \ANSWER/mem[1][7][5] ,
         \ANSWER/mem[1][7][4] , \ANSWER/mem[1][7][3] , \ANSWER/mem[1][7][2] ,
         \ANSWER/mem[1][7][1] , \ANSWER/mem[1][7][0] , \ANSWER/mem[1][6][15] ,
         \ANSWER/mem[1][6][14] , \ANSWER/mem[1][6][13] ,
         \ANSWER/mem[1][6][12] , \ANSWER/mem[1][6][11] ,
         \ANSWER/mem[1][6][10] , \ANSWER/mem[1][6][9] , \ANSWER/mem[1][6][8] ,
         \ANSWER/mem[1][6][7] , \ANSWER/mem[1][6][6] , \ANSWER/mem[1][6][5] ,
         \ANSWER/mem[1][6][4] , \ANSWER/mem[1][6][3] , \ANSWER/mem[1][6][2] ,
         \ANSWER/mem[1][6][1] , \ANSWER/mem[1][6][0] , \ANSWER/mem[1][5][15] ,
         \ANSWER/mem[1][5][14] , \ANSWER/mem[1][5][13] ,
         \ANSWER/mem[1][5][12] , \ANSWER/mem[1][5][11] ,
         \ANSWER/mem[1][5][10] , \ANSWER/mem[1][5][9] , \ANSWER/mem[1][5][8] ,
         \ANSWER/mem[1][5][7] , \ANSWER/mem[1][5][6] , \ANSWER/mem[1][5][5] ,
         \ANSWER/mem[1][5][4] , \ANSWER/mem[1][5][3] , \ANSWER/mem[1][5][2] ,
         \ANSWER/mem[1][5][1] , \ANSWER/mem[1][5][0] , \ANSWER/mem[1][4][15] ,
         \ANSWER/mem[1][4][14] , \ANSWER/mem[1][4][13] ,
         \ANSWER/mem[1][4][12] , \ANSWER/mem[1][4][11] ,
         \ANSWER/mem[1][4][10] , \ANSWER/mem[1][4][9] , \ANSWER/mem[1][4][8] ,
         \ANSWER/mem[1][4][7] , \ANSWER/mem[1][4][6] , \ANSWER/mem[1][4][5] ,
         \ANSWER/mem[1][4][4] , \ANSWER/mem[1][4][3] , \ANSWER/mem[1][4][2] ,
         \ANSWER/mem[1][4][1] , \ANSWER/mem[1][4][0] , \ANSWER/mem[1][3][15] ,
         \ANSWER/mem[1][3][14] , \ANSWER/mem[1][3][13] ,
         \ANSWER/mem[1][3][12] , \ANSWER/mem[1][3][11] ,
         \ANSWER/mem[1][3][10] , \ANSWER/mem[1][3][9] , \ANSWER/mem[1][3][8] ,
         \ANSWER/mem[1][3][7] , \ANSWER/mem[1][3][6] , \ANSWER/mem[1][3][5] ,
         \ANSWER/mem[1][3][4] , \ANSWER/mem[1][3][3] , \ANSWER/mem[1][3][2] ,
         \ANSWER/mem[1][3][1] , \ANSWER/mem[1][3][0] , \ANSWER/mem[1][2][15] ,
         \ANSWER/mem[1][2][14] , \ANSWER/mem[1][2][13] ,
         \ANSWER/mem[1][2][12] , \ANSWER/mem[1][2][11] ,
         \ANSWER/mem[1][2][10] , \ANSWER/mem[1][2][9] , \ANSWER/mem[1][2][8] ,
         \ANSWER/mem[1][2][7] , \ANSWER/mem[1][2][6] , \ANSWER/mem[1][2][5] ,
         \ANSWER/mem[1][2][4] , \ANSWER/mem[1][2][3] , \ANSWER/mem[1][2][2] ,
         \ANSWER/mem[1][2][1] , \ANSWER/mem[1][2][0] , \ANSWER/mem[1][1][15] ,
         \ANSWER/mem[1][1][14] , \ANSWER/mem[1][1][13] ,
         \ANSWER/mem[1][1][12] , \ANSWER/mem[1][1][11] ,
         \ANSWER/mem[1][1][10] , \ANSWER/mem[1][1][9] , \ANSWER/mem[1][1][8] ,
         \ANSWER/mem[1][1][7] , \ANSWER/mem[1][1][6] , \ANSWER/mem[1][1][5] ,
         \ANSWER/mem[1][1][4] , \ANSWER/mem[1][1][3] , \ANSWER/mem[1][1][2] ,
         \ANSWER/mem[1][1][1] , \ANSWER/mem[1][1][0] , \ANSWER/mem[1][0][15] ,
         \ANSWER/mem[1][0][14] , \ANSWER/mem[1][0][13] ,
         \ANSWER/mem[1][0][12] , \ANSWER/mem[1][0][11] ,
         \ANSWER/mem[1][0][10] , \ANSWER/mem[1][0][9] , \ANSWER/mem[1][0][8] ,
         \ANSWER/mem[1][0][7] , \ANSWER/mem[1][0][6] , \ANSWER/mem[1][0][5] ,
         \ANSWER/mem[1][0][4] , \ANSWER/mem[1][0][3] , \ANSWER/mem[1][0][2] ,
         \ANSWER/mem[1][0][1] , \ANSWER/mem[1][0][0] , \ANSWER/mem[0][9][15] ,
         \ANSWER/mem[0][9][14] , \ANSWER/mem[0][9][13] ,
         \ANSWER/mem[0][9][12] , \ANSWER/mem[0][9][11] ,
         \ANSWER/mem[0][9][10] , \ANSWER/mem[0][9][9] , \ANSWER/mem[0][9][8] ,
         \ANSWER/mem[0][9][7] , \ANSWER/mem[0][9][6] , \ANSWER/mem[0][9][5] ,
         \ANSWER/mem[0][9][4] , \ANSWER/mem[0][9][3] , \ANSWER/mem[0][9][2] ,
         \ANSWER/mem[0][9][1] , \ANSWER/mem[0][9][0] , \ANSWER/mem[0][8][15] ,
         \ANSWER/mem[0][8][14] , \ANSWER/mem[0][8][13] ,
         \ANSWER/mem[0][8][12] , \ANSWER/mem[0][8][11] ,
         \ANSWER/mem[0][8][10] , \ANSWER/mem[0][8][9] , \ANSWER/mem[0][8][8] ,
         \ANSWER/mem[0][8][7] , \ANSWER/mem[0][8][6] , \ANSWER/mem[0][8][5] ,
         \ANSWER/mem[0][8][4] , \ANSWER/mem[0][8][3] , \ANSWER/mem[0][8][2] ,
         \ANSWER/mem[0][8][1] , \ANSWER/mem[0][8][0] , \ANSWER/mem[0][7][15] ,
         \ANSWER/mem[0][7][14] , \ANSWER/mem[0][7][13] ,
         \ANSWER/mem[0][7][12] , \ANSWER/mem[0][7][11] ,
         \ANSWER/mem[0][7][10] , \ANSWER/mem[0][7][9] , \ANSWER/mem[0][7][8] ,
         \ANSWER/mem[0][7][7] , \ANSWER/mem[0][7][6] , \ANSWER/mem[0][7][5] ,
         \ANSWER/mem[0][7][4] , \ANSWER/mem[0][7][3] , \ANSWER/mem[0][7][2] ,
         \ANSWER/mem[0][7][1] , \ANSWER/mem[0][7][0] , \ANSWER/mem[0][6][15] ,
         \ANSWER/mem[0][6][14] , \ANSWER/mem[0][6][13] ,
         \ANSWER/mem[0][6][12] , \ANSWER/mem[0][6][11] ,
         \ANSWER/mem[0][6][10] , \ANSWER/mem[0][6][9] , \ANSWER/mem[0][6][8] ,
         \ANSWER/mem[0][6][7] , \ANSWER/mem[0][6][6] , \ANSWER/mem[0][6][5] ,
         \ANSWER/mem[0][6][4] , \ANSWER/mem[0][6][3] , \ANSWER/mem[0][6][2] ,
         \ANSWER/mem[0][6][1] , \ANSWER/mem[0][6][0] , \ANSWER/mem[0][5][15] ,
         \ANSWER/mem[0][5][14] , \ANSWER/mem[0][5][13] ,
         \ANSWER/mem[0][5][12] , \ANSWER/mem[0][5][11] ,
         \ANSWER/mem[0][5][10] , \ANSWER/mem[0][5][9] , \ANSWER/mem[0][5][8] ,
         \ANSWER/mem[0][5][7] , \ANSWER/mem[0][5][6] , \ANSWER/mem[0][5][5] ,
         \ANSWER/mem[0][5][4] , \ANSWER/mem[0][5][3] , \ANSWER/mem[0][5][2] ,
         \ANSWER/mem[0][5][1] , \ANSWER/mem[0][5][0] , \ANSWER/mem[0][4][15] ,
         \ANSWER/mem[0][4][14] , \ANSWER/mem[0][4][13] ,
         \ANSWER/mem[0][4][12] , \ANSWER/mem[0][4][11] ,
         \ANSWER/mem[0][4][10] , \ANSWER/mem[0][4][9] , \ANSWER/mem[0][4][8] ,
         \ANSWER/mem[0][4][7] , \ANSWER/mem[0][4][6] , \ANSWER/mem[0][4][5] ,
         \ANSWER/mem[0][4][4] , \ANSWER/mem[0][4][3] , \ANSWER/mem[0][4][2] ,
         \ANSWER/mem[0][4][1] , \ANSWER/mem[0][4][0] , \ANSWER/mem[0][3][15] ,
         \ANSWER/mem[0][3][14] , \ANSWER/mem[0][3][13] ,
         \ANSWER/mem[0][3][12] , \ANSWER/mem[0][3][11] ,
         \ANSWER/mem[0][3][10] , \ANSWER/mem[0][3][9] , \ANSWER/mem[0][3][8] ,
         \ANSWER/mem[0][3][7] , \ANSWER/mem[0][3][6] , \ANSWER/mem[0][3][5] ,
         \ANSWER/mem[0][3][4] , \ANSWER/mem[0][3][3] , \ANSWER/mem[0][3][2] ,
         \ANSWER/mem[0][3][1] , \ANSWER/mem[0][3][0] , \ANSWER/mem[0][2][15] ,
         \ANSWER/mem[0][2][14] , \ANSWER/mem[0][2][13] ,
         \ANSWER/mem[0][2][12] , \ANSWER/mem[0][2][11] ,
         \ANSWER/mem[0][2][10] , \ANSWER/mem[0][2][9] , \ANSWER/mem[0][2][8] ,
         \ANSWER/mem[0][2][7] , \ANSWER/mem[0][2][6] , \ANSWER/mem[0][2][5] ,
         \ANSWER/mem[0][2][4] , \ANSWER/mem[0][2][3] , \ANSWER/mem[0][2][2] ,
         \ANSWER/mem[0][2][1] , \ANSWER/mem[0][2][0] , \ANSWER/mem[0][1][15] ,
         \ANSWER/mem[0][1][14] , \ANSWER/mem[0][1][13] ,
         \ANSWER/mem[0][1][12] , \ANSWER/mem[0][1][11] ,
         \ANSWER/mem[0][1][10] , \ANSWER/mem[0][1][9] , \ANSWER/mem[0][1][8] ,
         \ANSWER/mem[0][1][7] , \ANSWER/mem[0][1][6] , \ANSWER/mem[0][1][5] ,
         \ANSWER/mem[0][1][4] , \ANSWER/mem[0][1][3] , \ANSWER/mem[0][1][2] ,
         \ANSWER/mem[0][1][1] , \ANSWER/mem[0][1][0] , \ANSWER/mem[0][0][15] ,
         \ANSWER/mem[0][0][14] , \ANSWER/mem[0][0][13] ,
         \ANSWER/mem[0][0][12] , \ANSWER/mem[0][0][11] ,
         \ANSWER/mem[0][0][10] , \ANSWER/mem[0][0][9] , \ANSWER/mem[0][0][8] ,
         \ANSWER/mem[0][0][7] , \ANSWER/mem[0][0][6] , \ANSWER/mem[0][0][5] ,
         \ANSWER/mem[0][0][4] , \ANSWER/mem[0][0][3] , \ANSWER/mem[0][0][2] ,
         \ANSWER/mem[0][0][1] , \ANSWER/mem[0][0][0] , \SIGMOID/N64 ,
         \SIGMOID/sign_bit , n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218;
  wire   [159:0] m1Inputs;
  wire   [159:0] column;
  wire   [15:0] m2DataIn;
  wire   [15:0] q_w2;
  wire   [15:0] \STAGE_1/weightReg ;
  wire   [15:0] \STAGE_1/M1/sum ;
  wire   [15:0] \STAGE_1/M2/sum ;
  wire   [15:0] \STAGE_1/M3/sum ;
  wire   [15:0] \STAGE_1/M4/sum ;
  wire   [15:0] \STAGE_1/M5/sum ;
  wire   [15:0] \STAGE_1/M6/sum ;
  wire   [15:0] \STAGE_1/M7/sum ;
  wire   [15:0] \STAGE_1/M8/sum ;
  wire   [15:0] \STAGE_1/M9/sum ;
  wire   [15:0] \STAGE_1/M10/sum ;
  wire   [4:0] \CNTRL/count_20Q ;
  wire   [3:0] \CNTRL/count_10_2Q ;
  wire   [3:0] \CNTRL/count_10Q ;
  wire   [7:0] \CNTRL/count_layer1_200Q ;
  wire   [9:0] \CNTRL/count_layer1_784Q ;
  wire   [3:0] \CNTRL/currentState ;
  wire   [159:0] \ROUTEDATA/regData ;
  wire   [15:0] \SIGMOID/lut_out ;

  dp_1 \STAGE_1/weightReg_reg[1]  ( .ip(weight1[1]), .ck(clk), .q(
        \STAGE_1/weightReg [1]) );
  dp_1 \STAGE_1/weightReg_reg[2]  ( .ip(weight1[2]), .ck(clk), .q(
        \STAGE_1/weightReg [2]) );
  dp_1 \STAGE_1/weightReg_reg[3]  ( .ip(weight1[3]), .ck(clk), .q(
        \STAGE_1/weightReg [3]) );
  dp_1 \STAGE_1/weightReg_reg[4]  ( .ip(weight1[4]), .ck(clk), .q(
        \STAGE_1/weightReg [4]) );
  dp_1 \STAGE_1/weightReg_reg[5]  ( .ip(weight1[5]), .ck(clk), .q(
        \STAGE_1/weightReg [5]) );
  dp_1 \STAGE_1/weightReg_reg[6]  ( .ip(weight1[6]), .ck(clk), .q(
        \STAGE_1/weightReg [6]) );
  dp_1 \STAGE_1/M1/result_reg[0]  ( .ip(\STAGE_1/M1/sum [0]), .ck(clk), .q(
        column[0]) );
  dp_1 \STAGE_1/M1/result_reg[1]  ( .ip(\STAGE_1/M1/sum [1]), .ck(clk), .q(
        column[1]) );
  dp_1 \STAGE_1/M1/result_reg[2]  ( .ip(\STAGE_1/M1/sum [2]), .ck(clk), .q(
        column[2]) );
  dp_1 \STAGE_1/M1/result_reg[3]  ( .ip(\STAGE_1/M1/sum [3]), .ck(clk), .q(
        column[3]) );
  dp_1 \STAGE_1/M1/result_reg[4]  ( .ip(\STAGE_1/M1/sum [4]), .ck(clk), .q(
        column[4]) );
  dp_1 \STAGE_1/M1/result_reg[5]  ( .ip(\STAGE_1/M1/sum [5]), .ck(clk), .q(
        column[5]) );
  dp_1 \STAGE_1/M1/result_reg[6]  ( .ip(\STAGE_1/M1/sum [6]), .ck(clk), .q(
        column[6]) );
  dp_1 \STAGE_1/M1/result_reg[7]  ( .ip(\STAGE_1/M1/sum [7]), .ck(clk), .q(
        column[7]) );
  dp_1 \STAGE_1/M1/result_reg[8]  ( .ip(\STAGE_1/M1/sum [8]), .ck(clk), .q(
        column[8]) );
  dp_1 \STAGE_1/M1/result_reg[9]  ( .ip(\STAGE_1/M1/sum [9]), .ck(clk), .q(
        column[9]) );
  dp_1 \STAGE_1/M1/result_reg[10]  ( .ip(\STAGE_1/M1/sum [10]), .ck(clk), .q(
        column[10]) );
  dp_1 \STAGE_1/M1/result_reg[11]  ( .ip(\STAGE_1/M1/sum [11]), .ck(clk), .q(
        column[11]) );
  dp_1 \STAGE_1/M1/result_reg[12]  ( .ip(\STAGE_1/M1/sum [12]), .ck(clk), .q(
        column[12]) );
  dp_1 \STAGE_1/M1/result_reg[13]  ( .ip(\STAGE_1/M1/sum [13]), .ck(clk), .q(
        column[13]) );
  dp_1 \STAGE_1/M1/result_reg[14]  ( .ip(\STAGE_1/M1/sum [14]), .ck(clk), .q(
        column[14]) );
  dp_1 \STAGE_1/M1/result_reg[15]  ( .ip(\STAGE_1/M1/sum [15]), .ck(clk), .q(
        column[15]) );
  dp_1 \STAGE_1/M2/result_reg[0]  ( .ip(\STAGE_1/M2/sum [0]), .ck(clk), .q(
        column[16]) );
  dp_1 \STAGE_1/M2/result_reg[1]  ( .ip(\STAGE_1/M2/sum [1]), .ck(clk), .q(
        column[17]) );
  dp_1 \STAGE_1/M2/result_reg[2]  ( .ip(\STAGE_1/M2/sum [2]), .ck(clk), .q(
        column[18]) );
  dp_1 \STAGE_1/M2/result_reg[3]  ( .ip(\STAGE_1/M2/sum [3]), .ck(clk), .q(
        column[19]) );
  dp_1 \STAGE_1/M2/result_reg[4]  ( .ip(\STAGE_1/M2/sum [4]), .ck(clk), .q(
        column[20]) );
  dp_1 \STAGE_1/M2/result_reg[5]  ( .ip(\STAGE_1/M2/sum [5]), .ck(clk), .q(
        column[21]) );
  dp_1 \STAGE_1/M2/result_reg[6]  ( .ip(\STAGE_1/M2/sum [6]), .ck(clk), .q(
        column[22]) );
  dp_1 \STAGE_1/M2/result_reg[7]  ( .ip(\STAGE_1/M2/sum [7]), .ck(clk), .q(
        column[23]) );
  dp_1 \STAGE_1/M2/result_reg[8]  ( .ip(\STAGE_1/M2/sum [8]), .ck(clk), .q(
        column[24]) );
  dp_1 \STAGE_1/M2/result_reg[9]  ( .ip(\STAGE_1/M2/sum [9]), .ck(clk), .q(
        column[25]) );
  dp_1 \STAGE_1/M2/result_reg[10]  ( .ip(\STAGE_1/M2/sum [10]), .ck(clk), .q(
        column[26]) );
  dp_1 \STAGE_1/M2/result_reg[11]  ( .ip(\STAGE_1/M2/sum [11]), .ck(clk), .q(
        column[27]) );
  dp_1 \STAGE_1/M2/result_reg[12]  ( .ip(\STAGE_1/M2/sum [12]), .ck(clk), .q(
        column[28]) );
  dp_1 \STAGE_1/M2/result_reg[13]  ( .ip(\STAGE_1/M2/sum [13]), .ck(clk), .q(
        column[29]) );
  dp_1 \STAGE_1/M2/result_reg[14]  ( .ip(\STAGE_1/M2/sum [14]), .ck(clk), .q(
        column[30]) );
  dp_1 \STAGE_1/M2/result_reg[15]  ( .ip(\STAGE_1/M2/sum [15]), .ck(clk), .q(
        column[31]) );
  dp_1 \STAGE_1/M3/result_reg[0]  ( .ip(\STAGE_1/M3/sum [0]), .ck(clk), .q(
        column[32]) );
  dp_1 \STAGE_1/M3/result_reg[1]  ( .ip(\STAGE_1/M3/sum [1]), .ck(clk), .q(
        column[33]) );
  dp_1 \STAGE_1/M3/result_reg[2]  ( .ip(\STAGE_1/M3/sum [2]), .ck(clk), .q(
        column[34]) );
  dp_1 \STAGE_1/M3/result_reg[3]  ( .ip(\STAGE_1/M3/sum [3]), .ck(clk), .q(
        column[35]) );
  dp_1 \STAGE_1/M3/result_reg[4]  ( .ip(\STAGE_1/M3/sum [4]), .ck(clk), .q(
        column[36]) );
  dp_1 \STAGE_1/M3/result_reg[5]  ( .ip(\STAGE_1/M3/sum [5]), .ck(clk), .q(
        column[37]) );
  dp_1 \STAGE_1/M3/result_reg[6]  ( .ip(\STAGE_1/M3/sum [6]), .ck(clk), .q(
        column[38]) );
  dp_1 \STAGE_1/M3/result_reg[7]  ( .ip(\STAGE_1/M3/sum [7]), .ck(clk), .q(
        column[39]) );
  dp_1 \STAGE_1/M3/result_reg[8]  ( .ip(\STAGE_1/M3/sum [8]), .ck(clk), .q(
        column[40]) );
  dp_1 \STAGE_1/M3/result_reg[9]  ( .ip(\STAGE_1/M3/sum [9]), .ck(clk), .q(
        column[41]) );
  dp_1 \STAGE_1/M3/result_reg[10]  ( .ip(\STAGE_1/M3/sum [10]), .ck(clk), .q(
        column[42]) );
  dp_1 \STAGE_1/M3/result_reg[11]  ( .ip(\STAGE_1/M3/sum [11]), .ck(clk), .q(
        column[43]) );
  dp_1 \STAGE_1/M3/result_reg[12]  ( .ip(\STAGE_1/M3/sum [12]), .ck(clk), .q(
        column[44]) );
  dp_1 \STAGE_1/M3/result_reg[13]  ( .ip(\STAGE_1/M3/sum [13]), .ck(clk), .q(
        column[45]) );
  dp_1 \STAGE_1/M3/result_reg[14]  ( .ip(\STAGE_1/M3/sum [14]), .ck(clk), .q(
        column[46]) );
  dp_1 \STAGE_1/M3/result_reg[15]  ( .ip(\STAGE_1/M3/sum [15]), .ck(clk), .q(
        column[47]) );
  dp_1 \STAGE_1/M4/result_reg[0]  ( .ip(\STAGE_1/M4/sum [0]), .ck(clk), .q(
        column[48]) );
  dp_1 \STAGE_1/M4/result_reg[1]  ( .ip(\STAGE_1/M4/sum [1]), .ck(clk), .q(
        column[49]) );
  dp_1 \STAGE_1/M4/result_reg[2]  ( .ip(\STAGE_1/M4/sum [2]), .ck(clk), .q(
        column[50]) );
  dp_1 \STAGE_1/M4/result_reg[3]  ( .ip(\STAGE_1/M4/sum [3]), .ck(clk), .q(
        column[51]) );
  dp_1 \STAGE_1/M4/result_reg[4]  ( .ip(\STAGE_1/M4/sum [4]), .ck(clk), .q(
        column[52]) );
  dp_1 \STAGE_1/M4/result_reg[5]  ( .ip(\STAGE_1/M4/sum [5]), .ck(clk), .q(
        column[53]) );
  dp_1 \STAGE_1/M4/result_reg[6]  ( .ip(\STAGE_1/M4/sum [6]), .ck(clk), .q(
        column[54]) );
  dp_1 \STAGE_1/M4/result_reg[7]  ( .ip(\STAGE_1/M4/sum [7]), .ck(clk), .q(
        column[55]) );
  dp_1 \STAGE_1/M4/result_reg[8]  ( .ip(\STAGE_1/M4/sum [8]), .ck(clk), .q(
        column[56]) );
  dp_1 \STAGE_1/M4/result_reg[9]  ( .ip(\STAGE_1/M4/sum [9]), .ck(clk), .q(
        column[57]) );
  dp_1 \STAGE_1/M4/result_reg[10]  ( .ip(\STAGE_1/M4/sum [10]), .ck(clk), .q(
        column[58]) );
  dp_1 \STAGE_1/M4/result_reg[11]  ( .ip(\STAGE_1/M4/sum [11]), .ck(clk), .q(
        column[59]) );
  dp_1 \STAGE_1/M4/result_reg[12]  ( .ip(\STAGE_1/M4/sum [12]), .ck(clk), .q(
        column[60]) );
  dp_1 \STAGE_1/M4/result_reg[13]  ( .ip(\STAGE_1/M4/sum [13]), .ck(clk), .q(
        column[61]) );
  dp_1 \STAGE_1/M4/result_reg[14]  ( .ip(\STAGE_1/M4/sum [14]), .ck(clk), .q(
        column[62]) );
  dp_1 \STAGE_1/M4/result_reg[15]  ( .ip(\STAGE_1/M4/sum [15]), .ck(clk), .q(
        column[63]) );
  dp_1 \STAGE_1/M5/result_reg[0]  ( .ip(\STAGE_1/M5/sum [0]), .ck(clk), .q(
        column[64]) );
  dp_1 \STAGE_1/M5/result_reg[1]  ( .ip(\STAGE_1/M5/sum [1]), .ck(clk), .q(
        column[65]) );
  dp_1 \STAGE_1/M5/result_reg[2]  ( .ip(\STAGE_1/M5/sum [2]), .ck(clk), .q(
        column[66]) );
  dp_1 \STAGE_1/M5/result_reg[3]  ( .ip(\STAGE_1/M5/sum [3]), .ck(clk), .q(
        column[67]) );
  dp_1 \STAGE_1/M5/result_reg[4]  ( .ip(\STAGE_1/M5/sum [4]), .ck(clk), .q(
        column[68]) );
  dp_1 \STAGE_1/M5/result_reg[5]  ( .ip(\STAGE_1/M5/sum [5]), .ck(clk), .q(
        column[69]) );
  dp_1 \STAGE_1/M5/result_reg[6]  ( .ip(\STAGE_1/M5/sum [6]), .ck(clk), .q(
        column[70]) );
  dp_1 \STAGE_1/M5/result_reg[7]  ( .ip(\STAGE_1/M5/sum [7]), .ck(clk), .q(
        column[71]) );
  dp_1 \STAGE_1/M5/result_reg[8]  ( .ip(\STAGE_1/M5/sum [8]), .ck(clk), .q(
        column[72]) );
  dp_1 \STAGE_1/M5/result_reg[9]  ( .ip(\STAGE_1/M5/sum [9]), .ck(clk), .q(
        column[73]) );
  dp_1 \STAGE_1/M5/result_reg[10]  ( .ip(\STAGE_1/M5/sum [10]), .ck(clk), .q(
        column[74]) );
  dp_1 \STAGE_1/M5/result_reg[11]  ( .ip(\STAGE_1/M5/sum [11]), .ck(clk), .q(
        column[75]) );
  dp_1 \STAGE_1/M5/result_reg[12]  ( .ip(\STAGE_1/M5/sum [12]), .ck(clk), .q(
        column[76]) );
  dp_1 \STAGE_1/M5/result_reg[13]  ( .ip(\STAGE_1/M5/sum [13]), .ck(clk), .q(
        column[77]) );
  dp_1 \STAGE_1/M5/result_reg[14]  ( .ip(\STAGE_1/M5/sum [14]), .ck(clk), .q(
        column[78]) );
  dp_1 \STAGE_1/M5/result_reg[15]  ( .ip(\STAGE_1/M5/sum [15]), .ck(clk), .q(
        column[79]) );
  dp_1 \STAGE_1/M6/result_reg[0]  ( .ip(\STAGE_1/M6/sum [0]), .ck(clk), .q(
        column[80]) );
  dp_1 \STAGE_1/M6/result_reg[1]  ( .ip(\STAGE_1/M6/sum [1]), .ck(clk), .q(
        column[81]) );
  dp_1 \STAGE_1/M6/result_reg[2]  ( .ip(\STAGE_1/M6/sum [2]), .ck(clk), .q(
        column[82]) );
  dp_1 \STAGE_1/M6/result_reg[3]  ( .ip(\STAGE_1/M6/sum [3]), .ck(clk), .q(
        column[83]) );
  dp_1 \STAGE_1/M6/result_reg[4]  ( .ip(\STAGE_1/M6/sum [4]), .ck(clk), .q(
        column[84]) );
  dp_1 \STAGE_1/M6/result_reg[5]  ( .ip(\STAGE_1/M6/sum [5]), .ck(clk), .q(
        column[85]) );
  dp_1 \STAGE_1/M6/result_reg[6]  ( .ip(\STAGE_1/M6/sum [6]), .ck(clk), .q(
        column[86]) );
  dp_1 \STAGE_1/M6/result_reg[7]  ( .ip(\STAGE_1/M6/sum [7]), .ck(clk), .q(
        column[87]) );
  dp_1 \STAGE_1/M6/result_reg[8]  ( .ip(\STAGE_1/M6/sum [8]), .ck(clk), .q(
        column[88]) );
  dp_1 \STAGE_1/M6/result_reg[9]  ( .ip(\STAGE_1/M6/sum [9]), .ck(clk), .q(
        column[89]) );
  dp_1 \STAGE_1/M6/result_reg[10]  ( .ip(\STAGE_1/M6/sum [10]), .ck(clk), .q(
        column[90]) );
  dp_1 \STAGE_1/M6/result_reg[11]  ( .ip(\STAGE_1/M6/sum [11]), .ck(clk), .q(
        column[91]) );
  dp_1 \STAGE_1/M6/result_reg[12]  ( .ip(\STAGE_1/M6/sum [12]), .ck(clk), .q(
        column[92]) );
  dp_1 \STAGE_1/M6/result_reg[13]  ( .ip(\STAGE_1/M6/sum [13]), .ck(clk), .q(
        column[93]) );
  dp_1 \STAGE_1/M6/result_reg[14]  ( .ip(\STAGE_1/M6/sum [14]), .ck(clk), .q(
        column[94]) );
  dp_1 \STAGE_1/M6/result_reg[15]  ( .ip(\STAGE_1/M6/sum [15]), .ck(clk), .q(
        column[95]) );
  dp_1 \STAGE_1/M7/result_reg[0]  ( .ip(\STAGE_1/M7/sum [0]), .ck(clk), .q(
        column[96]) );
  dp_1 \STAGE_1/M7/result_reg[1]  ( .ip(\STAGE_1/M7/sum [1]), .ck(clk), .q(
        column[97]) );
  dp_1 \STAGE_1/M7/result_reg[2]  ( .ip(\STAGE_1/M7/sum [2]), .ck(clk), .q(
        column[98]) );
  dp_1 \STAGE_1/M7/result_reg[3]  ( .ip(\STAGE_1/M7/sum [3]), .ck(clk), .q(
        column[99]) );
  dp_1 \STAGE_1/M7/result_reg[4]  ( .ip(\STAGE_1/M7/sum [4]), .ck(clk), .q(
        column[100]) );
  dp_1 \STAGE_1/M7/result_reg[5]  ( .ip(\STAGE_1/M7/sum [5]), .ck(clk), .q(
        column[101]) );
  dp_1 \STAGE_1/M7/result_reg[6]  ( .ip(\STAGE_1/M7/sum [6]), .ck(clk), .q(
        column[102]) );
  dp_1 \STAGE_1/M7/result_reg[7]  ( .ip(\STAGE_1/M7/sum [7]), .ck(clk), .q(
        column[103]) );
  dp_1 \STAGE_1/M7/result_reg[8]  ( .ip(\STAGE_1/M7/sum [8]), .ck(clk), .q(
        column[104]) );
  dp_1 \STAGE_1/M7/result_reg[9]  ( .ip(\STAGE_1/M7/sum [9]), .ck(clk), .q(
        column[105]) );
  dp_1 \STAGE_1/M7/result_reg[10]  ( .ip(\STAGE_1/M7/sum [10]), .ck(clk), .q(
        column[106]) );
  dp_1 \STAGE_1/M7/result_reg[11]  ( .ip(\STAGE_1/M7/sum [11]), .ck(clk), .q(
        column[107]) );
  dp_1 \STAGE_1/M7/result_reg[12]  ( .ip(\STAGE_1/M7/sum [12]), .ck(clk), .q(
        column[108]) );
  dp_1 \STAGE_1/M7/result_reg[13]  ( .ip(\STAGE_1/M7/sum [13]), .ck(clk), .q(
        column[109]) );
  dp_1 \STAGE_1/M7/result_reg[14]  ( .ip(\STAGE_1/M7/sum [14]), .ck(clk), .q(
        column[110]) );
  dp_1 \STAGE_1/M7/result_reg[15]  ( .ip(\STAGE_1/M7/sum [15]), .ck(clk), .q(
        column[111]) );
  dp_1 \STAGE_1/M8/result_reg[0]  ( .ip(\STAGE_1/M8/sum [0]), .ck(clk), .q(
        column[112]) );
  dp_1 \STAGE_1/M8/result_reg[1]  ( .ip(\STAGE_1/M8/sum [1]), .ck(clk), .q(
        column[113]) );
  dp_1 \STAGE_1/M8/result_reg[2]  ( .ip(\STAGE_1/M8/sum [2]), .ck(clk), .q(
        column[114]) );
  dp_1 \STAGE_1/M8/result_reg[3]  ( .ip(\STAGE_1/M8/sum [3]), .ck(clk), .q(
        column[115]) );
  dp_1 \STAGE_1/M8/result_reg[4]  ( .ip(\STAGE_1/M8/sum [4]), .ck(clk), .q(
        column[116]) );
  dp_1 \STAGE_1/M8/result_reg[5]  ( .ip(\STAGE_1/M8/sum [5]), .ck(clk), .q(
        column[117]) );
  dp_1 \STAGE_1/M8/result_reg[6]  ( .ip(\STAGE_1/M8/sum [6]), .ck(clk), .q(
        column[118]) );
  dp_1 \STAGE_1/M8/result_reg[7]  ( .ip(\STAGE_1/M8/sum [7]), .ck(clk), .q(
        column[119]) );
  dp_1 \STAGE_1/M8/result_reg[8]  ( .ip(\STAGE_1/M8/sum [8]), .ck(clk), .q(
        column[120]) );
  dp_1 \STAGE_1/M8/result_reg[9]  ( .ip(\STAGE_1/M8/sum [9]), .ck(clk), .q(
        column[121]) );
  dp_1 \STAGE_1/M8/result_reg[10]  ( .ip(\STAGE_1/M8/sum [10]), .ck(clk), .q(
        column[122]) );
  dp_1 \STAGE_1/M8/result_reg[11]  ( .ip(\STAGE_1/M8/sum [11]), .ck(clk), .q(
        column[123]) );
  dp_1 \STAGE_1/M8/result_reg[12]  ( .ip(\STAGE_1/M8/sum [12]), .ck(clk), .q(
        column[124]) );
  dp_1 \STAGE_1/M8/result_reg[13]  ( .ip(\STAGE_1/M8/sum [13]), .ck(clk), .q(
        column[125]) );
  dp_1 \STAGE_1/M8/result_reg[14]  ( .ip(\STAGE_1/M8/sum [14]), .ck(clk), .q(
        column[126]) );
  dp_1 \STAGE_1/M8/result_reg[15]  ( .ip(\STAGE_1/M8/sum [15]), .ck(clk), .q(
        column[127]) );
  dp_1 \STAGE_1/M9/result_reg[0]  ( .ip(\STAGE_1/M9/sum [0]), .ck(clk), .q(
        column[128]) );
  dp_1 \STAGE_1/M9/result_reg[1]  ( .ip(\STAGE_1/M9/sum [1]), .ck(clk), .q(
        column[129]) );
  dp_1 \STAGE_1/M9/result_reg[2]  ( .ip(\STAGE_1/M9/sum [2]), .ck(clk), .q(
        column[130]) );
  dp_1 \STAGE_1/M9/result_reg[3]  ( .ip(\STAGE_1/M9/sum [3]), .ck(clk), .q(
        column[131]) );
  dp_1 \STAGE_1/M9/result_reg[4]  ( .ip(\STAGE_1/M9/sum [4]), .ck(clk), .q(
        column[132]) );
  dp_1 \STAGE_1/M9/result_reg[5]  ( .ip(\STAGE_1/M9/sum [5]), .ck(clk), .q(
        column[133]) );
  dp_1 \STAGE_1/M9/result_reg[6]  ( .ip(\STAGE_1/M9/sum [6]), .ck(clk), .q(
        column[134]) );
  dp_1 \STAGE_1/M9/result_reg[7]  ( .ip(\STAGE_1/M9/sum [7]), .ck(clk), .q(
        column[135]) );
  dp_1 \STAGE_1/M9/result_reg[8]  ( .ip(\STAGE_1/M9/sum [8]), .ck(clk), .q(
        column[136]) );
  dp_1 \STAGE_1/M9/result_reg[9]  ( .ip(\STAGE_1/M9/sum [9]), .ck(clk), .q(
        column[137]) );
  dp_1 \STAGE_1/M9/result_reg[10]  ( .ip(\STAGE_1/M9/sum [10]), .ck(clk), .q(
        column[138]) );
  dp_1 \STAGE_1/M9/result_reg[11]  ( .ip(\STAGE_1/M9/sum [11]), .ck(clk), .q(
        column[139]) );
  dp_1 \STAGE_1/M9/result_reg[12]  ( .ip(\STAGE_1/M9/sum [12]), .ck(clk), .q(
        column[140]) );
  dp_1 \STAGE_1/M9/result_reg[13]  ( .ip(\STAGE_1/M9/sum [13]), .ck(clk), .q(
        column[141]) );
  dp_1 \STAGE_1/M9/result_reg[14]  ( .ip(\STAGE_1/M9/sum [14]), .ck(clk), .q(
        column[142]) );
  dp_1 \STAGE_1/M9/result_reg[15]  ( .ip(\STAGE_1/M9/sum [15]), .ck(clk), .q(
        column[143]) );
  dp_1 \STAGE_1/M10/result_reg[0]  ( .ip(\STAGE_1/M10/sum [0]), .ck(clk), .q(
        column[144]) );
  dp_1 \STAGE_1/M10/result_reg[1]  ( .ip(\STAGE_1/M10/sum [1]), .ck(clk), .q(
        column[145]) );
  dp_1 \STAGE_1/M10/result_reg[2]  ( .ip(\STAGE_1/M10/sum [2]), .ck(clk), .q(
        column[146]) );
  dp_1 \STAGE_1/M10/result_reg[3]  ( .ip(\STAGE_1/M10/sum [3]), .ck(clk), .q(
        column[147]) );
  dp_1 \STAGE_1/M10/result_reg[4]  ( .ip(\STAGE_1/M10/sum [4]), .ck(clk), .q(
        column[148]) );
  dp_1 \STAGE_1/M10/result_reg[5]  ( .ip(\STAGE_1/M10/sum [5]), .ck(clk), .q(
        column[149]) );
  dp_1 \STAGE_1/M10/result_reg[6]  ( .ip(\STAGE_1/M10/sum [6]), .ck(clk), .q(
        column[150]) );
  dp_1 \STAGE_1/M10/result_reg[7]  ( .ip(\STAGE_1/M10/sum [7]), .ck(clk), .q(
        column[151]) );
  dp_1 \STAGE_1/M10/result_reg[8]  ( .ip(\STAGE_1/M10/sum [8]), .ck(clk), .q(
        column[152]) );
  dp_1 \STAGE_1/M10/result_reg[9]  ( .ip(\STAGE_1/M10/sum [9]), .ck(clk), .q(
        column[153]) );
  dp_1 \STAGE_1/M10/result_reg[10]  ( .ip(\STAGE_1/M10/sum [10]), .ck(clk), 
        .q(column[154]) );
  dp_1 \STAGE_1/M10/result_reg[11]  ( .ip(\STAGE_1/M10/sum [11]), .ck(clk), 
        .q(column[155]) );
  dp_1 \STAGE_1/M10/result_reg[12]  ( .ip(\STAGE_1/M10/sum [12]), .ck(clk), 
        .q(column[156]) );
  dp_1 \STAGE_1/M10/result_reg[13]  ( .ip(\STAGE_1/M10/sum [13]), .ck(clk), 
        .q(column[157]) );
  dp_1 \STAGE_1/M10/result_reg[14]  ( .ip(\STAGE_1/M10/sum [14]), .ck(clk), 
        .q(column[158]) );
  dp_1 \STAGE_1/M10/result_reg[15]  ( .ip(\STAGE_1/M10/sum [15]), .ck(clk), 
        .q(column[159]) );
  dp_1 \INPUTSRAM/q_reg[0]  ( .ip(\INPUTSRAM/mem_i[0][0] ), .ck(clk), .q(
        m1Inputs[0]) );
  dp_1 \INPUTSRAM/q_reg[1]  ( .ip(\INPUTSRAM/mem_i[0][1] ), .ck(clk), .q(
        m1Inputs[1]) );
  dp_1 \INPUTSRAM/q_reg[3]  ( .ip(\INPUTSRAM/mem_i[0][3] ), .ck(clk), .q(
        m1Inputs[3]) );
  dp_1 \INPUTSRAM/q_reg[5]  ( .ip(\INPUTSRAM/mem_i[0][5] ), .ck(clk), .q(
        m1Inputs[5]) );
  dp_1 \INPUTSRAM/q_reg[6]  ( .ip(\INPUTSRAM/mem_i[0][6] ), .ck(clk), .q(
        m1Inputs[6]) );
  dp_1 \INPUTSRAM/q_reg[7]  ( .ip(\INPUTSRAM/mem_i[0][7] ), .ck(clk), .q(
        m1Inputs[7]) );
  dp_1 \INPUTSRAM/q_reg[16]  ( .ip(\INPUTSRAM/mem_i[1][0] ), .ck(clk), .q(
        m1Inputs[16]) );
  dp_1 \INPUTSRAM/q_reg[17]  ( .ip(\INPUTSRAM/mem_i[1][1] ), .ck(clk), .q(
        m1Inputs[17]) );
  dp_1 \INPUTSRAM/q_reg[19]  ( .ip(\INPUTSRAM/mem_i[1][3] ), .ck(clk), .q(
        m1Inputs[19]) );
  dp_1 \INPUTSRAM/q_reg[20]  ( .ip(\INPUTSRAM/mem_i[1][4] ), .ck(clk), .q(
        m1Inputs[20]) );
  dp_1 \INPUTSRAM/q_reg[21]  ( .ip(\INPUTSRAM/mem_i[1][5] ), .ck(clk), .q(
        m1Inputs[21]) );
  dp_1 \INPUTSRAM/q_reg[22]  ( .ip(\INPUTSRAM/mem_i[1][6] ), .ck(clk), .q(
        m1Inputs[22]) );
  dp_1 \INPUTSRAM/q_reg[23]  ( .ip(\INPUTSRAM/mem_i[1][7] ), .ck(clk), .q(
        m1Inputs[23]) );
  dp_1 \INPUTSRAM/q_reg[32]  ( .ip(\INPUTSRAM/mem_i[2][0] ), .ck(clk), .q(
        m1Inputs[32]) );
  dp_1 \INPUTSRAM/q_reg[33]  ( .ip(\INPUTSRAM/mem_i[2][1] ), .ck(clk), .q(
        m1Inputs[33]) );
  dp_1 \INPUTSRAM/q_reg[35]  ( .ip(\INPUTSRAM/mem_i[2][3] ), .ck(clk), .q(
        m1Inputs[35]) );
  dp_1 \INPUTSRAM/q_reg[36]  ( .ip(\INPUTSRAM/mem_i[2][4] ), .ck(clk), .q(
        m1Inputs[36]) );
  dp_1 \INPUTSRAM/q_reg[37]  ( .ip(\INPUTSRAM/mem_i[2][5] ), .ck(clk), .q(
        m1Inputs[37]) );
  dp_1 \INPUTSRAM/q_reg[38]  ( .ip(\INPUTSRAM/mem_i[2][6] ), .ck(clk), .q(
        m1Inputs[38]) );
  dp_1 \INPUTSRAM/q_reg[39]  ( .ip(\INPUTSRAM/mem_i[2][7] ), .ck(clk), .q(
        m1Inputs[39]) );
  dp_1 \INPUTSRAM/q_reg[40]  ( .ip(\INPUTSRAM/mem_i[2][8] ), .ck(clk), .q(
        m1Inputs[40]) );
  dp_1 \INPUTSRAM/q_reg[48]  ( .ip(\INPUTSRAM/mem_i[3][0] ), .ck(clk), .q(
        m1Inputs[48]) );
  dp_1 \INPUTSRAM/q_reg[49]  ( .ip(\INPUTSRAM/mem_i[3][1] ), .ck(clk), .q(
        m1Inputs[49]) );
  dp_1 \INPUTSRAM/q_reg[51]  ( .ip(\INPUTSRAM/mem_i[3][3] ), .ck(clk), .q(
        m1Inputs[51]) );
  dp_1 \INPUTSRAM/q_reg[52]  ( .ip(\INPUTSRAM/mem_i[3][4] ), .ck(clk), .q(
        m1Inputs[52]) );
  dp_1 \INPUTSRAM/q_reg[53]  ( .ip(\INPUTSRAM/mem_i[3][5] ), .ck(clk), .q(
        m1Inputs[53]) );
  dp_1 \INPUTSRAM/q_reg[54]  ( .ip(\INPUTSRAM/mem_i[3][6] ), .ck(clk), .q(
        m1Inputs[54]) );
  dp_1 \INPUTSRAM/q_reg[55]  ( .ip(\INPUTSRAM/mem_i[3][7] ), .ck(clk), .q(
        m1Inputs[55]) );
  dp_1 \INPUTSRAM/q_reg[64]  ( .ip(\INPUTSRAM/mem_i[4][0] ), .ck(clk), .q(
        m1Inputs[64]) );
  dp_1 \INPUTSRAM/q_reg[65]  ( .ip(\INPUTSRAM/mem_i[4][1] ), .ck(clk), .q(
        m1Inputs[65]) );
  dp_1 \INPUTSRAM/q_reg[67]  ( .ip(\INPUTSRAM/mem_i[4][3] ), .ck(clk), .q(
        m1Inputs[67]) );
  dp_1 \INPUTSRAM/q_reg[68]  ( .ip(\INPUTSRAM/mem_i[4][4] ), .ck(clk), .q(
        m1Inputs[68]) );
  dp_1 \INPUTSRAM/q_reg[69]  ( .ip(\INPUTSRAM/mem_i[4][5] ), .ck(clk), .q(
        m1Inputs[69]) );
  dp_1 \INPUTSRAM/q_reg[70]  ( .ip(\INPUTSRAM/mem_i[4][6] ), .ck(clk), .q(
        m1Inputs[70]) );
  dp_1 \INPUTSRAM/q_reg[71]  ( .ip(\INPUTSRAM/mem_i[4][7] ), .ck(clk), .q(
        m1Inputs[71]) );
  dp_1 \INPUTSRAM/q_reg[72]  ( .ip(\INPUTSRAM/mem_i[4][8] ), .ck(clk), .q(
        m1Inputs[72]) );
  dp_1 \INPUTSRAM/q_reg[80]  ( .ip(\INPUTSRAM/mem_i[5][0] ), .ck(clk), .q(
        m1Inputs[80]) );
  dp_1 \INPUTSRAM/q_reg[81]  ( .ip(\INPUTSRAM/mem_i[5][1] ), .ck(clk), .q(
        m1Inputs[81]) );
  dp_1 \INPUTSRAM/q_reg[83]  ( .ip(\INPUTSRAM/mem_i[5][3] ), .ck(clk), .q(
        m1Inputs[83]) );
  dp_1 \INPUTSRAM/q_reg[84]  ( .ip(\INPUTSRAM/mem_i[5][4] ), .ck(clk), .q(
        m1Inputs[84]) );
  dp_1 \INPUTSRAM/q_reg[85]  ( .ip(\INPUTSRAM/mem_i[5][5] ), .ck(clk), .q(
        m1Inputs[85]) );
  dp_1 \INPUTSRAM/q_reg[86]  ( .ip(\INPUTSRAM/mem_i[5][6] ), .ck(clk), .q(
        m1Inputs[86]) );
  dp_1 \INPUTSRAM/q_reg[87]  ( .ip(\INPUTSRAM/mem_i[5][7] ), .ck(clk), .q(
        m1Inputs[87]) );
  dp_1 \INPUTSRAM/q_reg[96]  ( .ip(\INPUTSRAM/mem_i[6][0] ), .ck(clk), .q(
        m1Inputs[96]) );
  dp_1 \INPUTSRAM/q_reg[97]  ( .ip(\INPUTSRAM/mem_i[6][1] ), .ck(clk), .q(
        m1Inputs[97]) );
  dp_1 \INPUTSRAM/q_reg[99]  ( .ip(\INPUTSRAM/mem_i[6][3] ), .ck(clk), .q(
        m1Inputs[99]) );
  dp_1 \INPUTSRAM/q_reg[100]  ( .ip(\INPUTSRAM/mem_i[6][4] ), .ck(clk), .q(
        m1Inputs[100]) );
  dp_1 \INPUTSRAM/q_reg[101]  ( .ip(\INPUTSRAM/mem_i[6][5] ), .ck(clk), .q(
        m1Inputs[101]) );
  dp_1 \INPUTSRAM/q_reg[102]  ( .ip(\INPUTSRAM/mem_i[6][6] ), .ck(clk), .q(
        m1Inputs[102]) );
  dp_1 \INPUTSRAM/q_reg[103]  ( .ip(\INPUTSRAM/mem_i[6][7] ), .ck(clk), .q(
        m1Inputs[103]) );
  dp_1 \INPUTSRAM/q_reg[104]  ( .ip(\INPUTSRAM/mem_i[6][8] ), .ck(clk), .q(
        m1Inputs[104]) );
  dp_1 \INPUTSRAM/q_reg[112]  ( .ip(\INPUTSRAM/mem_i[7][0] ), .ck(clk), .q(
        m1Inputs[112]) );
  dp_1 \INPUTSRAM/q_reg[113]  ( .ip(\INPUTSRAM/mem_i[7][1] ), .ck(clk), .q(
        m1Inputs[113]) );
  dp_1 \INPUTSRAM/q_reg[115]  ( .ip(\INPUTSRAM/mem_i[7][3] ), .ck(clk), .q(
        m1Inputs[115]) );
  dp_1 \INPUTSRAM/q_reg[116]  ( .ip(\INPUTSRAM/mem_i[7][4] ), .ck(clk), .q(
        m1Inputs[116]) );
  dp_1 \INPUTSRAM/q_reg[117]  ( .ip(\INPUTSRAM/mem_i[7][5] ), .ck(clk), .q(
        m1Inputs[117]) );
  dp_1 \INPUTSRAM/q_reg[118]  ( .ip(\INPUTSRAM/mem_i[7][6] ), .ck(clk), .q(
        m1Inputs[118]) );
  dp_1 \INPUTSRAM/q_reg[119]  ( .ip(\INPUTSRAM/mem_i[7][7] ), .ck(clk), .q(
        m1Inputs[119]) );
  dp_1 \INPUTSRAM/q_reg[120]  ( .ip(\INPUTSRAM/mem_i[7][8] ), .ck(clk), .q(
        m1Inputs[120]) );
  dp_1 \INPUTSRAM/q_reg[128]  ( .ip(\INPUTSRAM/mem_i[8][0] ), .ck(clk), .q(
        m1Inputs[128]) );
  dp_1 \INPUTSRAM/q_reg[129]  ( .ip(\INPUTSRAM/mem_i[8][1] ), .ck(clk), .q(
        m1Inputs[129]) );
  dp_1 \INPUTSRAM/q_reg[131]  ( .ip(\INPUTSRAM/mem_i[8][3] ), .ck(clk), .q(
        m1Inputs[131]) );
  dp_1 \INPUTSRAM/q_reg[132]  ( .ip(\INPUTSRAM/mem_i[8][4] ), .ck(clk), .q(
        m1Inputs[132]) );
  dp_1 \INPUTSRAM/q_reg[133]  ( .ip(\INPUTSRAM/mem_i[8][5] ), .ck(clk), .q(
        m1Inputs[133]) );
  dp_1 \INPUTSRAM/q_reg[134]  ( .ip(\INPUTSRAM/mem_i[8][6] ), .ck(clk), .q(
        m1Inputs[134]) );
  dp_1 \INPUTSRAM/q_reg[135]  ( .ip(\INPUTSRAM/mem_i[8][7] ), .ck(clk), .q(
        m1Inputs[135]) );
  dp_1 \INPUTSRAM/q_reg[144]  ( .ip(\INPUTSRAM/mem_i[9][0] ), .ck(clk), .q(
        m1Inputs[144]) );
  dp_1 \INPUTSRAM/q_reg[145]  ( .ip(\INPUTSRAM/mem_i[9][1] ), .ck(clk), .q(
        m1Inputs[145]) );
  dp_1 \INPUTSRAM/q_reg[147]  ( .ip(\INPUTSRAM/mem_i[9][3] ), .ck(clk), .q(
        m1Inputs[147]) );
  dp_1 \INPUTSRAM/q_reg[148]  ( .ip(\INPUTSRAM/mem_i[9][4] ), .ck(clk), .q(
        m1Inputs[148]) );
  dp_1 \INPUTSRAM/q_reg[149]  ( .ip(\INPUTSRAM/mem_i[9][5] ), .ck(clk), .q(
        m1Inputs[149]) );
  dp_1 \INPUTSRAM/q_reg[150]  ( .ip(\INPUTSRAM/mem_i[9][6] ), .ck(clk), .q(
        m1Inputs[150]) );
  dp_1 \INPUTSRAM/q_reg[151]  ( .ip(\INPUTSRAM/mem_i[9][7] ), .ck(clk), .q(
        m1Inputs[151]) );
  dp_1 \INPUTSRAM/q_reg[152]  ( .ip(\INPUTSRAM/mem_i[9][8] ), .ck(clk), .q(
        m1Inputs[152]) );
  dp_1 \CNTRL/count_20Q_reg[4]  ( .ip(n4043), .ck(clk), .q(
        \CNTRL/count_20Q [4]) );
  dp_1 \CNTRL/count_10Q_reg[3]  ( .ip(n4027), .ck(clk), .q(
        \CNTRL/count_10Q [3]) );
  dp_1 \CNTRL/currentState_reg[0]  ( .ip(n4039), .ck(clk), .q(
        \CNTRL/currentState [0]) );
  dp_1 \CNTRL/count_layer1_200Q_reg[7]  ( .ip(n4019), .ck(clk), .q(
        \CNTRL/count_layer1_200Q [7]) );
  dp_1 \CNTRL/count_layer1_784Q_reg[9]  ( .ip(\CNTRL/N242 ), .ck(clk), .q(
        \CNTRL/count_layer1_784Q [9]) );
  dp_1 \CNTRL/currentState_reg[1]  ( .ip(n4040), .ck(clk), .q(
        \CNTRL/currentState [1]) );
  dp_1 \CNTRL/currentState_reg[2]  ( .ip(n4041), .ck(clk), .q(
        \CNTRL/currentState [2]) );
  dp_1 \CNTRL/count_20Q_reg[0]  ( .ip(n4038), .ck(clk), .q(
        \CNTRL/count_20Q [0]) );
  dp_1 \CNTRL/count_20Q_reg[1]  ( .ip(n4037), .ck(clk), .q(
        \CNTRL/count_20Q [1]) );
  dp_1 \CNTRL/count_20Q_reg[2]  ( .ip(n4036), .ck(clk), .q(
        \CNTRL/count_20Q [2]) );
  dp_1 \CNTRL/count_20Q_reg[3]  ( .ip(n4035), .ck(clk), .q(
        \CNTRL/count_20Q [3]) );
  dp_1 \CNTRL/count_10Q_reg[0]  ( .ip(n4030), .ck(clk), .q(
        \CNTRL/count_10Q [0]) );
  dp_1 \CNTRL/count_10Q_reg[1]  ( .ip(n4029), .ck(clk), .q(
        \CNTRL/count_10Q [1]) );
  dp_1 \CNTRL/count_10Q_reg[2]  ( .ip(n4028), .ck(clk), .q(
        \CNTRL/count_10Q [2]) );
  dp_1 \CNTRL/count_layer1_784Q_reg[0]  ( .ip(\CNTRL/N233 ), .ck(clk), .q(
        \CNTRL/count_layer1_784Q [0]) );
  dp_1 \CNTRL/count_layer1_784Q_reg[1]  ( .ip(\CNTRL/N234 ), .ck(clk), .q(
        \CNTRL/count_layer1_784Q [1]) );
  dp_1 \CNTRL/count_layer1_784Q_reg[2]  ( .ip(\CNTRL/N235 ), .ck(clk), .q(
        \CNTRL/count_layer1_784Q [2]) );
  dp_1 \CNTRL/count_layer1_784Q_reg[3]  ( .ip(\CNTRL/N236 ), .ck(clk), .q(
        \CNTRL/count_layer1_784Q [3]) );
  dp_1 \CNTRL/count_layer1_784Q_reg[4]  ( .ip(\CNTRL/N237 ), .ck(clk), .q(
        \CNTRL/count_layer1_784Q [4]) );
  dp_1 \CNTRL/count_layer1_784Q_reg[5]  ( .ip(\CNTRL/N238 ), .ck(clk), .q(
        \CNTRL/count_layer1_784Q [5]) );
  dp_1 \CNTRL/count_layer1_784Q_reg[6]  ( .ip(\CNTRL/N239 ), .ck(clk), .q(
        \CNTRL/count_layer1_784Q [6]) );
  dp_1 \CNTRL/count_layer1_784Q_reg[7]  ( .ip(\CNTRL/N240 ), .ck(clk), .q(
        \CNTRL/count_layer1_784Q [7]) );
  dp_1 \CNTRL/count_layer1_784Q_reg[8]  ( .ip(\CNTRL/N241 ), .ck(clk), .q(
        \CNTRL/count_layer1_784Q [8]) );
  dp_1 \CNTRL/count_layer1_200Q_reg[1]  ( .ip(n4026), .ck(clk), .q(
        \CNTRL/count_layer1_200Q [1]) );
  dp_1 \CNTRL/count_layer1_200Q_reg[0]  ( .ip(n4025), .ck(clk), .q(
        \CNTRL/count_layer1_200Q [0]) );
  dp_1 \CNTRL/count_layer1_200Q_reg[2]  ( .ip(n4024), .ck(clk), .q(
        \CNTRL/count_layer1_200Q [2]) );
  dp_1 \CNTRL/count_layer1_200Q_reg[3]  ( .ip(n4023), .ck(clk), .q(
        \CNTRL/count_layer1_200Q [3]) );
  dp_1 \CNTRL/count_layer1_200Q_reg[4]  ( .ip(n4022), .ck(clk), .q(
        \CNTRL/count_layer1_200Q [4]) );
  dp_1 \CNTRL/count_layer1_200Q_reg[5]  ( .ip(n4021), .ck(clk), .q(
        \CNTRL/count_layer1_200Q [5]) );
  dp_1 \CNTRL/count_layer1_200Q_reg[6]  ( .ip(n4020), .ck(clk), .q(
        \CNTRL/count_layer1_200Q [6]) );
  dp_1 \CNTRL/count_10_2Q_reg[0]  ( .ip(n4034), .ck(clk), .q(
        \CNTRL/count_10_2Q [0]) );
  dp_1 \CNTRL/count_10_2Q_reg[1]  ( .ip(n4033), .ck(clk), .q(
        \CNTRL/count_10_2Q [1]) );
  dp_1 \CNTRL/count_10_2Q_reg[2]  ( .ip(n4032), .ck(clk), .q(
        \CNTRL/count_10_2Q [2]) );
  dp_1 \CNTRL/count_10_2Q_reg[3]  ( .ip(n4031), .ck(clk), .q(
        \CNTRL/count_10_2Q [3]) );
  dp_1 \ROUTEDATA/DataToM2_reg[0]  ( .ip(n4018), .ck(clk), .q(m2DataIn[0]) );
  dp_1 \ROUTEDATA/DataToM2_reg[1]  ( .ip(n4017), .ck(clk), .q(m2DataIn[1]) );
  dp_1 \ROUTEDATA/DataToM2_reg[2]  ( .ip(n4016), .ck(clk), .q(m2DataIn[2]) );
  dp_1 \ROUTEDATA/DataToM2_reg[3]  ( .ip(n4015), .ck(clk), .q(m2DataIn[3]) );
  dp_1 \ROUTEDATA/DataToM2_reg[4]  ( .ip(n4014), .ck(clk), .q(m2DataIn[4]) );
  dp_1 \ROUTEDATA/DataToM2_reg[5]  ( .ip(n4013), .ck(clk), .q(m2DataIn[5]) );
  dp_1 \ROUTEDATA/DataToM2_reg[6]  ( .ip(n4012), .ck(clk), .q(m2DataIn[6]) );
  dp_1 \ROUTEDATA/DataToM2_reg[7]  ( .ip(n4011), .ck(clk), .q(m2DataIn[7]) );
  dp_1 \ROUTEDATA/DataToM2_reg[8]  ( .ip(n4010), .ck(clk), .q(m2DataIn[8]) );
  dp_1 \ROUTEDATA/DataToM2_reg[9]  ( .ip(n4009), .ck(clk), .q(m2DataIn[9]) );
  dp_1 \ROUTEDATA/DataToM2_reg[10]  ( .ip(n4008), .ck(clk), .q(m2DataIn[10])
         );
  dp_1 \ROUTEDATA/DataToM2_reg[11]  ( .ip(n4007), .ck(clk), .q(m2DataIn[11])
         );
  dp_1 \ROUTEDATA/DataToM2_reg[12]  ( .ip(n4006), .ck(clk), .q(m2DataIn[12])
         );
  dp_1 \ROUTEDATA/DataToM2_reg[13]  ( .ip(n4005), .ck(clk), .q(m2DataIn[13])
         );
  dp_1 \ROUTEDATA/DataToM2_reg[14]  ( .ip(n4004), .ck(clk), .q(m2DataIn[14])
         );
  dp_1 \ROUTEDATA/DataToM2_reg[15]  ( .ip(n4003), .ck(clk), .q(m2DataIn[15])
         );
  dp_1 \WEIGHT_2/mem_w2_reg[0][0]  ( .ip(n4002), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][0] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][1]  ( .ip(n4001), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][1] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][2]  ( .ip(n4000), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][2] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][3]  ( .ip(n3999), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][3] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][4]  ( .ip(n3998), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][4] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][5]  ( .ip(n3997), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][5] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][6]  ( .ip(n3996), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][6] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][7]  ( .ip(n3995), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][7] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][8]  ( .ip(n3994), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][8] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][9]  ( .ip(n3993), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][9] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][10]  ( .ip(n3992), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][10] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][11]  ( .ip(n3991), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][11] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][12]  ( .ip(n3990), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][12] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][13]  ( .ip(n3989), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][13] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][14]  ( .ip(n3988), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][14] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][15]  ( .ip(n3987), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][15] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][0]  ( .ip(n3986), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][0] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][1]  ( .ip(n3985), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][1] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][2]  ( .ip(n3984), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][2] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][3]  ( .ip(n3983), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][3] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][4]  ( .ip(n3982), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][4] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][5]  ( .ip(n3981), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][5] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][6]  ( .ip(n3980), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][6] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][7]  ( .ip(n3979), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][7] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][8]  ( .ip(n3978), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][8] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][9]  ( .ip(n3977), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][9] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][10]  ( .ip(n3976), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][10] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][11]  ( .ip(n3975), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][11] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][12]  ( .ip(n3974), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][12] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][13]  ( .ip(n3973), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][13] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][14]  ( .ip(n3972), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][14] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][15]  ( .ip(n3971), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][15] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][0]  ( .ip(n3970), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][0] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][1]  ( .ip(n3969), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][1] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][2]  ( .ip(n3968), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][2] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][3]  ( .ip(n3967), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][3] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][4]  ( .ip(n3966), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][4] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][5]  ( .ip(n3965), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][5] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][6]  ( .ip(n3964), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][6] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][7]  ( .ip(n3963), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][7] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][8]  ( .ip(n3962), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][8] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][9]  ( .ip(n3961), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][9] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][10]  ( .ip(n3960), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][10] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][11]  ( .ip(n3959), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][11] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][12]  ( .ip(n3958), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][12] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][13]  ( .ip(n3957), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][13] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][14]  ( .ip(n3956), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][14] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][15]  ( .ip(n3955), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][15] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][0]  ( .ip(n3954), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][0] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][1]  ( .ip(n3953), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][1] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][2]  ( .ip(n3952), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][2] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][3]  ( .ip(n3951), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][3] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][4]  ( .ip(n3950), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][4] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][5]  ( .ip(n3949), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][5] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][6]  ( .ip(n3948), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][6] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][7]  ( .ip(n3947), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][7] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][8]  ( .ip(n3946), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][8] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][9]  ( .ip(n3945), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][9] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][10]  ( .ip(n3944), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][10] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][11]  ( .ip(n3943), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][11] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][12]  ( .ip(n3942), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][12] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][13]  ( .ip(n3941), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][13] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][14]  ( .ip(n3940), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][14] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][15]  ( .ip(n3939), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][15] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][0]  ( .ip(n3938), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][0] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][1]  ( .ip(n3937), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][1] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][2]  ( .ip(n3936), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][2] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][3]  ( .ip(n3935), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][3] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][4]  ( .ip(n3934), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][4] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][5]  ( .ip(n3933), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][5] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][6]  ( .ip(n3932), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][6] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][7]  ( .ip(n3931), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][7] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][8]  ( .ip(n3930), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][8] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][9]  ( .ip(n3929), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][9] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][10]  ( .ip(n3928), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][10] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][11]  ( .ip(n3927), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][11] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][12]  ( .ip(n3926), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][12] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][13]  ( .ip(n3925), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][13] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][14]  ( .ip(n3924), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][14] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][15]  ( .ip(n3923), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][15] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][0]  ( .ip(n3922), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][0] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][1]  ( .ip(n3921), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][1] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][2]  ( .ip(n3920), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][2] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][3]  ( .ip(n3919), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][3] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][4]  ( .ip(n3918), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][4] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][5]  ( .ip(n3917), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][5] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][6]  ( .ip(n3916), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][6] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][7]  ( .ip(n3915), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][7] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][8]  ( .ip(n3914), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][8] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][9]  ( .ip(n3913), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][9] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][10]  ( .ip(n3912), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][10] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][11]  ( .ip(n3911), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][11] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][12]  ( .ip(n3910), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][12] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][13]  ( .ip(n3909), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][13] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][14]  ( .ip(n3908), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][14] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][15]  ( .ip(n3907), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][15] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][0]  ( .ip(n3906), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][0] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][1]  ( .ip(n3905), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][1] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][2]  ( .ip(n3904), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][2] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][3]  ( .ip(n3903), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][3] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][4]  ( .ip(n3902), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][4] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][5]  ( .ip(n3901), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][5] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][6]  ( .ip(n3900), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][6] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][7]  ( .ip(n3899), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][7] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][8]  ( .ip(n3898), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][8] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][9]  ( .ip(n3897), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][9] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][10]  ( .ip(n3896), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][10] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][11]  ( .ip(n3895), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][11] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][12]  ( .ip(n3894), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][12] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][13]  ( .ip(n3893), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][13] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][14]  ( .ip(n3892), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][14] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][15]  ( .ip(n3891), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][15] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][0]  ( .ip(n3890), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][0] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][1]  ( .ip(n3889), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][1] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][2]  ( .ip(n3888), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][2] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][3]  ( .ip(n3887), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][3] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][4]  ( .ip(n3886), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][4] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][5]  ( .ip(n3885), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][5] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][6]  ( .ip(n3884), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][6] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][7]  ( .ip(n3883), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][7] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][8]  ( .ip(n3882), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][8] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][9]  ( .ip(n3881), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][9] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][10]  ( .ip(n3880), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][10] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][11]  ( .ip(n3879), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][11] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][12]  ( .ip(n3878), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][12] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][13]  ( .ip(n3877), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][13] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][14]  ( .ip(n3876), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][14] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][15]  ( .ip(n3875), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][15] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][0]  ( .ip(n3874), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][0] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][1]  ( .ip(n3873), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][1] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][2]  ( .ip(n3872), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][2] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][3]  ( .ip(n3871), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][3] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][4]  ( .ip(n3870), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][4] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][5]  ( .ip(n3869), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][5] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][6]  ( .ip(n3868), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][6] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][7]  ( .ip(n3867), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][7] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][8]  ( .ip(n3866), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][8] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][9]  ( .ip(n3865), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][9] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][10]  ( .ip(n3864), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][10] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][11]  ( .ip(n3863), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][11] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][12]  ( .ip(n3862), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][12] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][13]  ( .ip(n3861), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][13] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][14]  ( .ip(n3860), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][14] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][15]  ( .ip(n3859), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][15] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][0]  ( .ip(n3858), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][0] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][1]  ( .ip(n3857), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][1] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][2]  ( .ip(n3856), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][2] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][3]  ( .ip(n3855), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][3] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][4]  ( .ip(n3854), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][4] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][5]  ( .ip(n3853), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][5] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][6]  ( .ip(n3852), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][6] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][7]  ( .ip(n3851), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][7] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][8]  ( .ip(n3850), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][8] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][9]  ( .ip(n3849), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][9] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][10]  ( .ip(n3848), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][10] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][11]  ( .ip(n3847), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][11] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][12]  ( .ip(n3846), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][12] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][13]  ( .ip(n3845), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][13] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][14]  ( .ip(n3844), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][14] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][15]  ( .ip(n3843), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][15] ) );
  dp_1 \ANSWER/rdata_reg[0]  ( .ip(\ANSWER/N487 ), .ck(clk), .q(rdata[0]) );
  dp_1 \ANSWER/rdata_reg[1]  ( .ip(\ANSWER/N486 ), .ck(clk), .q(rdata[1]) );
  dp_1 \ANSWER/rdata_reg[2]  ( .ip(\ANSWER/N485 ), .ck(clk), .q(rdata[2]) );
  dp_1 \ANSWER/rdata_reg[3]  ( .ip(\ANSWER/N484 ), .ck(clk), .q(rdata[3]) );
  dp_1 \ANSWER/rdata_reg[4]  ( .ip(\ANSWER/N483 ), .ck(clk), .q(rdata[4]) );
  dp_1 \ANSWER/rdata_reg[5]  ( .ip(\ANSWER/N482 ), .ck(clk), .q(rdata[5]) );
  dp_1 \ANSWER/rdata_reg[6]  ( .ip(\ANSWER/N481 ), .ck(clk), .q(rdata[6]) );
  dp_1 \ANSWER/rdata_reg[7]  ( .ip(\ANSWER/N480 ), .ck(clk), .q(rdata[7]) );
  dp_1 \ANSWER/rdata_reg[8]  ( .ip(\ANSWER/N479 ), .ck(clk), .q(rdata[8]) );
  dp_1 \ANSWER/rdata_reg[9]  ( .ip(\ANSWER/N478 ), .ck(clk), .q(rdata[9]) );
  dp_1 \ANSWER/rdata_reg[10]  ( .ip(\ANSWER/N477 ), .ck(clk), .q(rdata[10]) );
  dp_1 \ANSWER/rdata_reg[11]  ( .ip(\ANSWER/N476 ), .ck(clk), .q(rdata[11]) );
  dp_1 \ANSWER/rdata_reg[12]  ( .ip(\ANSWER/N475 ), .ck(clk), .q(rdata[12]) );
  dp_1 \ANSWER/rdata_reg[13]  ( .ip(\ANSWER/N474 ), .ck(clk), .q(rdata[13]) );
  dp_1 \ANSWER/rdata_reg[14]  ( .ip(\ANSWER/N473 ), .ck(clk), .q(rdata[14]) );
  dp_1 \ANSWER/rdata_reg[15]  ( .ip(\ANSWER/N472 ), .ck(clk), .q(rdata[15]) );
  dp_1 \SIGMOID/sign_bit_reg  ( .ip(\sig_in[15] ), .ck(clk), .q(
        \SIGMOID/sign_bit ) );
  dp_1 \ANSWER/mem_reg[0][0][8]  ( .ip(n3034), .ck(clk), .q(
        \ANSWER/mem[0][0][8] ) );
  dp_1 \ANSWER/mem_reg[0][1][8]  ( .ip(n3033), .ck(clk), .q(
        \ANSWER/mem[0][1][8] ) );
  dp_1 \ANSWER/mem_reg[0][2][8]  ( .ip(n3032), .ck(clk), .q(
        \ANSWER/mem[0][2][8] ) );
  dp_1 \ANSWER/mem_reg[0][3][8]  ( .ip(n3031), .ck(clk), .q(
        \ANSWER/mem[0][3][8] ) );
  dp_1 \ANSWER/mem_reg[0][4][8]  ( .ip(n3030), .ck(clk), .q(
        \ANSWER/mem[0][4][8] ) );
  dp_1 \ANSWER/mem_reg[0][5][8]  ( .ip(n3029), .ck(clk), .q(
        \ANSWER/mem[0][5][8] ) );
  dp_1 \ANSWER/mem_reg[0][6][8]  ( .ip(n3028), .ck(clk), .q(
        \ANSWER/mem[0][6][8] ) );
  dp_1 \ANSWER/mem_reg[0][7][8]  ( .ip(n3027), .ck(clk), .q(
        \ANSWER/mem[0][7][8] ) );
  dp_1 \ANSWER/mem_reg[0][8][8]  ( .ip(n3026), .ck(clk), .q(
        \ANSWER/mem[0][8][8] ) );
  dp_1 \ANSWER/mem_reg[0][9][8]  ( .ip(n3025), .ck(clk), .q(
        \ANSWER/mem[0][9][8] ) );
  dp_1 \ANSWER/mem_reg[1][0][8]  ( .ip(n3024), .ck(clk), .q(
        \ANSWER/mem[1][0][8] ) );
  dp_1 \ANSWER/mem_reg[1][1][8]  ( .ip(n3023), .ck(clk), .q(
        \ANSWER/mem[1][1][8] ) );
  dp_1 \ANSWER/mem_reg[1][2][8]  ( .ip(n3022), .ck(clk), .q(
        \ANSWER/mem[1][2][8] ) );
  dp_1 \ANSWER/mem_reg[1][3][8]  ( .ip(n3021), .ck(clk), .q(
        \ANSWER/mem[1][3][8] ) );
  dp_1 \ANSWER/mem_reg[1][4][8]  ( .ip(n3020), .ck(clk), .q(
        \ANSWER/mem[1][4][8] ) );
  dp_1 \ANSWER/mem_reg[1][5][8]  ( .ip(n3019), .ck(clk), .q(
        \ANSWER/mem[1][5][8] ) );
  dp_1 \ANSWER/mem_reg[1][6][8]  ( .ip(n3018), .ck(clk), .q(
        \ANSWER/mem[1][6][8] ) );
  dp_1 \ANSWER/mem_reg[1][7][8]  ( .ip(n3017), .ck(clk), .q(
        \ANSWER/mem[1][7][8] ) );
  dp_1 \ANSWER/mem_reg[1][8][8]  ( .ip(n3016), .ck(clk), .q(
        \ANSWER/mem[1][8][8] ) );
  dp_1 \ANSWER/mem_reg[1][9][8]  ( .ip(n3015), .ck(clk), .q(
        \ANSWER/mem[1][9][8] ) );
  dp_1 \ANSWER/mem_reg[2][0][8]  ( .ip(n3014), .ck(clk), .q(
        \ANSWER/mem[2][0][8] ) );
  dp_1 \ANSWER/mem_reg[2][1][8]  ( .ip(n3013), .ck(clk), .q(
        \ANSWER/mem[2][1][8] ) );
  dp_1 \ANSWER/mem_reg[2][2][8]  ( .ip(n3012), .ck(clk), .q(
        \ANSWER/mem[2][2][8] ) );
  dp_1 \ANSWER/mem_reg[2][3][8]  ( .ip(n3011), .ck(clk), .q(
        \ANSWER/mem[2][3][8] ) );
  dp_1 \ANSWER/mem_reg[2][4][8]  ( .ip(n3010), .ck(clk), .q(
        \ANSWER/mem[2][4][8] ) );
  dp_1 \ANSWER/mem_reg[2][5][8]  ( .ip(n3009), .ck(clk), .q(
        \ANSWER/mem[2][5][8] ) );
  dp_1 \ANSWER/mem_reg[2][6][8]  ( .ip(n3008), .ck(clk), .q(
        \ANSWER/mem[2][6][8] ) );
  dp_1 \ANSWER/mem_reg[2][7][8]  ( .ip(n3007), .ck(clk), .q(
        \ANSWER/mem[2][7][8] ) );
  dp_1 \ANSWER/mem_reg[2][8][8]  ( .ip(n3006), .ck(clk), .q(
        \ANSWER/mem[2][8][8] ) );
  dp_1 \ANSWER/mem_reg[2][9][8]  ( .ip(n3005), .ck(clk), .q(
        \ANSWER/mem[2][9][8] ) );
  dp_1 \ANSWER/mem_reg[3][0][8]  ( .ip(n3004), .ck(clk), .q(
        \ANSWER/mem[3][0][8] ) );
  dp_1 \ANSWER/mem_reg[3][1][8]  ( .ip(n3003), .ck(clk), .q(
        \ANSWER/mem[3][1][8] ) );
  dp_1 \ANSWER/mem_reg[3][2][8]  ( .ip(n3002), .ck(clk), .q(
        \ANSWER/mem[3][2][8] ) );
  dp_1 \ANSWER/mem_reg[3][3][8]  ( .ip(n3001), .ck(clk), .q(
        \ANSWER/mem[3][3][8] ) );
  dp_1 \ANSWER/mem_reg[3][4][8]  ( .ip(n3000), .ck(clk), .q(
        \ANSWER/mem[3][4][8] ) );
  dp_1 \ANSWER/mem_reg[3][5][8]  ( .ip(n2999), .ck(clk), .q(
        \ANSWER/mem[3][5][8] ) );
  dp_1 \ANSWER/mem_reg[3][6][8]  ( .ip(n2998), .ck(clk), .q(
        \ANSWER/mem[3][6][8] ) );
  dp_1 \ANSWER/mem_reg[3][7][8]  ( .ip(n2997), .ck(clk), .q(
        \ANSWER/mem[3][7][8] ) );
  dp_1 \ANSWER/mem_reg[3][8][8]  ( .ip(n2996), .ck(clk), .q(
        \ANSWER/mem[3][8][8] ) );
  dp_1 \ANSWER/mem_reg[3][9][8]  ( .ip(n2995), .ck(clk), .q(
        \ANSWER/mem[3][9][8] ) );
  dp_1 \ANSWER/mem_reg[4][0][8]  ( .ip(n2994), .ck(clk), .q(
        \ANSWER/mem[4][0][8] ) );
  dp_1 \ANSWER/mem_reg[4][1][8]  ( .ip(n2993), .ck(clk), .q(
        \ANSWER/mem[4][1][8] ) );
  dp_1 \ANSWER/mem_reg[4][2][8]  ( .ip(n2992), .ck(clk), .q(
        \ANSWER/mem[4][2][8] ) );
  dp_1 \ANSWER/mem_reg[4][3][8]  ( .ip(n2991), .ck(clk), .q(
        \ANSWER/mem[4][3][8] ) );
  dp_1 \ANSWER/mem_reg[4][4][8]  ( .ip(n2990), .ck(clk), .q(
        \ANSWER/mem[4][4][8] ) );
  dp_1 \ANSWER/mem_reg[4][5][8]  ( .ip(n2989), .ck(clk), .q(
        \ANSWER/mem[4][5][8] ) );
  dp_1 \ANSWER/mem_reg[4][6][8]  ( .ip(n2988), .ck(clk), .q(
        \ANSWER/mem[4][6][8] ) );
  dp_1 \ANSWER/mem_reg[4][7][8]  ( .ip(n2987), .ck(clk), .q(
        \ANSWER/mem[4][7][8] ) );
  dp_1 \ANSWER/mem_reg[4][8][8]  ( .ip(n2986), .ck(clk), .q(
        \ANSWER/mem[4][8][8] ) );
  dp_1 \ANSWER/mem_reg[4][9][8]  ( .ip(n2985), .ck(clk), .q(
        \ANSWER/mem[4][9][8] ) );
  dp_1 \ANSWER/mem_reg[5][0][8]  ( .ip(n2984), .ck(clk), .q(
        \ANSWER/mem[5][0][8] ) );
  dp_1 \ANSWER/mem_reg[5][1][8]  ( .ip(n2983), .ck(clk), .q(
        \ANSWER/mem[5][1][8] ) );
  dp_1 \ANSWER/mem_reg[5][2][8]  ( .ip(n2982), .ck(clk), .q(
        \ANSWER/mem[5][2][8] ) );
  dp_1 \ANSWER/mem_reg[5][3][8]  ( .ip(n2981), .ck(clk), .q(
        \ANSWER/mem[5][3][8] ) );
  dp_1 \ANSWER/mem_reg[5][4][8]  ( .ip(n2980), .ck(clk), .q(
        \ANSWER/mem[5][4][8] ) );
  dp_1 \ANSWER/mem_reg[5][5][8]  ( .ip(n2979), .ck(clk), .q(
        \ANSWER/mem[5][5][8] ) );
  dp_1 \ANSWER/mem_reg[5][6][8]  ( .ip(n2978), .ck(clk), .q(
        \ANSWER/mem[5][6][8] ) );
  dp_1 \ANSWER/mem_reg[5][7][8]  ( .ip(n2977), .ck(clk), .q(
        \ANSWER/mem[5][7][8] ) );
  dp_1 \ANSWER/mem_reg[5][8][8]  ( .ip(n2976), .ck(clk), .q(
        \ANSWER/mem[5][8][8] ) );
  dp_1 \ANSWER/mem_reg[5][9][8]  ( .ip(n2975), .ck(clk), .q(
        \ANSWER/mem[5][9][8] ) );
  dp_1 \ANSWER/mem_reg[6][0][8]  ( .ip(n2974), .ck(clk), .q(
        \ANSWER/mem[6][0][8] ) );
  dp_1 \ANSWER/mem_reg[6][1][8]  ( .ip(n2973), .ck(clk), .q(
        \ANSWER/mem[6][1][8] ) );
  dp_1 \ANSWER/mem_reg[6][2][8]  ( .ip(n2972), .ck(clk), .q(
        \ANSWER/mem[6][2][8] ) );
  dp_1 \ANSWER/mem_reg[6][3][8]  ( .ip(n2971), .ck(clk), .q(
        \ANSWER/mem[6][3][8] ) );
  dp_1 \ANSWER/mem_reg[6][4][8]  ( .ip(n2970), .ck(clk), .q(
        \ANSWER/mem[6][4][8] ) );
  dp_1 \ANSWER/mem_reg[6][5][8]  ( .ip(n2969), .ck(clk), .q(
        \ANSWER/mem[6][5][8] ) );
  dp_1 \ANSWER/mem_reg[6][6][8]  ( .ip(n2968), .ck(clk), .q(
        \ANSWER/mem[6][6][8] ) );
  dp_1 \ANSWER/mem_reg[6][7][8]  ( .ip(n2967), .ck(clk), .q(
        \ANSWER/mem[6][7][8] ) );
  dp_1 \ANSWER/mem_reg[6][8][8]  ( .ip(n2966), .ck(clk), .q(
        \ANSWER/mem[6][8][8] ) );
  dp_1 \ANSWER/mem_reg[6][9][8]  ( .ip(n2965), .ck(clk), .q(
        \ANSWER/mem[6][9][8] ) );
  dp_1 \ANSWER/mem_reg[7][0][8]  ( .ip(n2964), .ck(clk), .q(
        \ANSWER/mem[7][0][8] ) );
  dp_1 \ANSWER/mem_reg[7][1][8]  ( .ip(n2963), .ck(clk), .q(
        \ANSWER/mem[7][1][8] ) );
  dp_1 \ANSWER/mem_reg[7][2][8]  ( .ip(n2962), .ck(clk), .q(
        \ANSWER/mem[7][2][8] ) );
  dp_1 \ANSWER/mem_reg[7][3][8]  ( .ip(n2961), .ck(clk), .q(
        \ANSWER/mem[7][3][8] ) );
  dp_1 \ANSWER/mem_reg[7][4][8]  ( .ip(n2960), .ck(clk), .q(
        \ANSWER/mem[7][4][8] ) );
  dp_1 \ANSWER/mem_reg[7][5][8]  ( .ip(n2959), .ck(clk), .q(
        \ANSWER/mem[7][5][8] ) );
  dp_1 \ANSWER/mem_reg[7][6][8]  ( .ip(n2958), .ck(clk), .q(
        \ANSWER/mem[7][6][8] ) );
  dp_1 \ANSWER/mem_reg[7][7][8]  ( .ip(n2957), .ck(clk), .q(
        \ANSWER/mem[7][7][8] ) );
  dp_1 \ANSWER/mem_reg[7][8][8]  ( .ip(n2956), .ck(clk), .q(
        \ANSWER/mem[7][8][8] ) );
  dp_1 \ANSWER/mem_reg[7][9][8]  ( .ip(n2955), .ck(clk), .q(
        \ANSWER/mem[7][9][8] ) );
  dp_1 \ANSWER/mem_reg[8][0][8]  ( .ip(n2954), .ck(clk), .q(
        \ANSWER/mem[8][0][8] ) );
  dp_1 \ANSWER/mem_reg[8][1][8]  ( .ip(n2953), .ck(clk), .q(
        \ANSWER/mem[8][1][8] ) );
  dp_1 \ANSWER/mem_reg[8][2][8]  ( .ip(n2952), .ck(clk), .q(
        \ANSWER/mem[8][2][8] ) );
  dp_1 \ANSWER/mem_reg[8][3][8]  ( .ip(n2951), .ck(clk), .q(
        \ANSWER/mem[8][3][8] ) );
  dp_1 \ANSWER/mem_reg[8][4][8]  ( .ip(n2950), .ck(clk), .q(
        \ANSWER/mem[8][4][8] ) );
  dp_1 \ANSWER/mem_reg[8][5][8]  ( .ip(n2949), .ck(clk), .q(
        \ANSWER/mem[8][5][8] ) );
  dp_1 \ANSWER/mem_reg[8][6][8]  ( .ip(n2948), .ck(clk), .q(
        \ANSWER/mem[8][6][8] ) );
  dp_1 \ANSWER/mem_reg[8][7][8]  ( .ip(n2947), .ck(clk), .q(
        \ANSWER/mem[8][7][8] ) );
  dp_1 \ANSWER/mem_reg[8][8][8]  ( .ip(n2946), .ck(clk), .q(
        \ANSWER/mem[8][8][8] ) );
  dp_1 \ANSWER/mem_reg[8][9][8]  ( .ip(n2945), .ck(clk), .q(
        \ANSWER/mem[8][9][8] ) );
  dp_1 \ANSWER/mem_reg[9][0][8]  ( .ip(n2944), .ck(clk), .q(
        \ANSWER/mem[9][0][8] ) );
  dp_1 \ANSWER/mem_reg[9][1][8]  ( .ip(n2943), .ck(clk), .q(
        \ANSWER/mem[9][1][8] ) );
  dp_1 \ANSWER/mem_reg[9][2][8]  ( .ip(n2942), .ck(clk), .q(
        \ANSWER/mem[9][2][8] ) );
  dp_1 \ANSWER/mem_reg[9][3][8]  ( .ip(n2941), .ck(clk), .q(
        \ANSWER/mem[9][3][8] ) );
  dp_1 \ANSWER/mem_reg[9][4][8]  ( .ip(n2940), .ck(clk), .q(
        \ANSWER/mem[9][4][8] ) );
  dp_1 \ANSWER/mem_reg[9][5][8]  ( .ip(n2939), .ck(clk), .q(
        \ANSWER/mem[9][5][8] ) );
  dp_1 \ANSWER/mem_reg[9][6][8]  ( .ip(n2938), .ck(clk), .q(
        \ANSWER/mem[9][6][8] ) );
  dp_1 \ANSWER/mem_reg[9][7][8]  ( .ip(n2937), .ck(clk), .q(
        \ANSWER/mem[9][7][8] ) );
  dp_1 \ANSWER/mem_reg[9][8][8]  ( .ip(n2936), .ck(clk), .q(
        \ANSWER/mem[9][8][8] ) );
  dp_1 \ANSWER/mem_reg[9][9][8]  ( .ip(n2935), .ck(clk), .q(
        \ANSWER/mem[9][9][8] ) );
  dp_1 \ANSWER/mem_reg[0][0][9]  ( .ip(n2934), .ck(clk), .q(
        \ANSWER/mem[0][0][9] ) );
  dp_1 \ANSWER/mem_reg[0][1][9]  ( .ip(n2933), .ck(clk), .q(
        \ANSWER/mem[0][1][9] ) );
  dp_1 \ANSWER/mem_reg[0][2][9]  ( .ip(n2932), .ck(clk), .q(
        \ANSWER/mem[0][2][9] ) );
  dp_1 \ANSWER/mem_reg[0][3][9]  ( .ip(n2931), .ck(clk), .q(
        \ANSWER/mem[0][3][9] ) );
  dp_1 \ANSWER/mem_reg[0][4][9]  ( .ip(n2930), .ck(clk), .q(
        \ANSWER/mem[0][4][9] ) );
  dp_1 \ANSWER/mem_reg[0][5][9]  ( .ip(n2929), .ck(clk), .q(
        \ANSWER/mem[0][5][9] ) );
  dp_1 \ANSWER/mem_reg[0][6][9]  ( .ip(n2928), .ck(clk), .q(
        \ANSWER/mem[0][6][9] ) );
  dp_1 \ANSWER/mem_reg[0][7][9]  ( .ip(n2927), .ck(clk), .q(
        \ANSWER/mem[0][7][9] ) );
  dp_1 \ANSWER/mem_reg[0][8][9]  ( .ip(n2926), .ck(clk), .q(
        \ANSWER/mem[0][8][9] ) );
  dp_1 \ANSWER/mem_reg[0][9][9]  ( .ip(n2925), .ck(clk), .q(
        \ANSWER/mem[0][9][9] ) );
  dp_1 \ANSWER/mem_reg[1][0][9]  ( .ip(n2924), .ck(clk), .q(
        \ANSWER/mem[1][0][9] ) );
  dp_1 \ANSWER/mem_reg[1][1][9]  ( .ip(n2923), .ck(clk), .q(
        \ANSWER/mem[1][1][9] ) );
  dp_1 \ANSWER/mem_reg[1][2][9]  ( .ip(n2922), .ck(clk), .q(
        \ANSWER/mem[1][2][9] ) );
  dp_1 \ANSWER/mem_reg[1][3][9]  ( .ip(n2921), .ck(clk), .q(
        \ANSWER/mem[1][3][9] ) );
  dp_1 \ANSWER/mem_reg[1][4][9]  ( .ip(n2920), .ck(clk), .q(
        \ANSWER/mem[1][4][9] ) );
  dp_1 \ANSWER/mem_reg[1][5][9]  ( .ip(n2919), .ck(clk), .q(
        \ANSWER/mem[1][5][9] ) );
  dp_1 \ANSWER/mem_reg[1][6][9]  ( .ip(n2918), .ck(clk), .q(
        \ANSWER/mem[1][6][9] ) );
  dp_1 \ANSWER/mem_reg[1][7][9]  ( .ip(n2917), .ck(clk), .q(
        \ANSWER/mem[1][7][9] ) );
  dp_1 \ANSWER/mem_reg[1][8][9]  ( .ip(n2916), .ck(clk), .q(
        \ANSWER/mem[1][8][9] ) );
  dp_1 \ANSWER/mem_reg[1][9][9]  ( .ip(n2915), .ck(clk), .q(
        \ANSWER/mem[1][9][9] ) );
  dp_1 \ANSWER/mem_reg[2][0][9]  ( .ip(n2914), .ck(clk), .q(
        \ANSWER/mem[2][0][9] ) );
  dp_1 \ANSWER/mem_reg[2][1][9]  ( .ip(n2913), .ck(clk), .q(
        \ANSWER/mem[2][1][9] ) );
  dp_1 \ANSWER/mem_reg[2][2][9]  ( .ip(n2912), .ck(clk), .q(
        \ANSWER/mem[2][2][9] ) );
  dp_1 \ANSWER/mem_reg[2][3][9]  ( .ip(n2911), .ck(clk), .q(
        \ANSWER/mem[2][3][9] ) );
  dp_1 \ANSWER/mem_reg[2][4][9]  ( .ip(n2910), .ck(clk), .q(
        \ANSWER/mem[2][4][9] ) );
  dp_1 \ANSWER/mem_reg[2][5][9]  ( .ip(n2909), .ck(clk), .q(
        \ANSWER/mem[2][5][9] ) );
  dp_1 \ANSWER/mem_reg[2][6][9]  ( .ip(n2908), .ck(clk), .q(
        \ANSWER/mem[2][6][9] ) );
  dp_1 \ANSWER/mem_reg[2][7][9]  ( .ip(n2907), .ck(clk), .q(
        \ANSWER/mem[2][7][9] ) );
  dp_1 \ANSWER/mem_reg[2][8][9]  ( .ip(n2906), .ck(clk), .q(
        \ANSWER/mem[2][8][9] ) );
  dp_1 \ANSWER/mem_reg[2][9][9]  ( .ip(n2905), .ck(clk), .q(
        \ANSWER/mem[2][9][9] ) );
  dp_1 \ANSWER/mem_reg[3][0][9]  ( .ip(n2904), .ck(clk), .q(
        \ANSWER/mem[3][0][9] ) );
  dp_1 \ANSWER/mem_reg[3][1][9]  ( .ip(n2903), .ck(clk), .q(
        \ANSWER/mem[3][1][9] ) );
  dp_1 \ANSWER/mem_reg[3][2][9]  ( .ip(n2902), .ck(clk), .q(
        \ANSWER/mem[3][2][9] ) );
  dp_1 \ANSWER/mem_reg[3][3][9]  ( .ip(n2901), .ck(clk), .q(
        \ANSWER/mem[3][3][9] ) );
  dp_1 \ANSWER/mem_reg[3][4][9]  ( .ip(n2900), .ck(clk), .q(
        \ANSWER/mem[3][4][9] ) );
  dp_1 \ANSWER/mem_reg[3][5][9]  ( .ip(n2899), .ck(clk), .q(
        \ANSWER/mem[3][5][9] ) );
  dp_1 \ANSWER/mem_reg[3][6][9]  ( .ip(n2898), .ck(clk), .q(
        \ANSWER/mem[3][6][9] ) );
  dp_1 \ANSWER/mem_reg[3][7][9]  ( .ip(n2897), .ck(clk), .q(
        \ANSWER/mem[3][7][9] ) );
  dp_1 \ANSWER/mem_reg[3][8][9]  ( .ip(n2896), .ck(clk), .q(
        \ANSWER/mem[3][8][9] ) );
  dp_1 \ANSWER/mem_reg[3][9][9]  ( .ip(n2895), .ck(clk), .q(
        \ANSWER/mem[3][9][9] ) );
  dp_1 \ANSWER/mem_reg[4][0][9]  ( .ip(n2894), .ck(clk), .q(
        \ANSWER/mem[4][0][9] ) );
  dp_1 \ANSWER/mem_reg[4][1][9]  ( .ip(n2893), .ck(clk), .q(
        \ANSWER/mem[4][1][9] ) );
  dp_1 \ANSWER/mem_reg[4][2][9]  ( .ip(n2892), .ck(clk), .q(
        \ANSWER/mem[4][2][9] ) );
  dp_1 \ANSWER/mem_reg[4][3][9]  ( .ip(n2891), .ck(clk), .q(
        \ANSWER/mem[4][3][9] ) );
  dp_1 \ANSWER/mem_reg[4][4][9]  ( .ip(n2890), .ck(clk), .q(
        \ANSWER/mem[4][4][9] ) );
  dp_1 \ANSWER/mem_reg[4][5][9]  ( .ip(n2889), .ck(clk), .q(
        \ANSWER/mem[4][5][9] ) );
  dp_1 \ANSWER/mem_reg[4][6][9]  ( .ip(n2888), .ck(clk), .q(
        \ANSWER/mem[4][6][9] ) );
  dp_1 \ANSWER/mem_reg[4][7][9]  ( .ip(n2887), .ck(clk), .q(
        \ANSWER/mem[4][7][9] ) );
  dp_1 \ANSWER/mem_reg[4][8][9]  ( .ip(n2886), .ck(clk), .q(
        \ANSWER/mem[4][8][9] ) );
  dp_1 \ANSWER/mem_reg[4][9][9]  ( .ip(n2885), .ck(clk), .q(
        \ANSWER/mem[4][9][9] ) );
  dp_1 \ANSWER/mem_reg[5][0][9]  ( .ip(n2884), .ck(clk), .q(
        \ANSWER/mem[5][0][9] ) );
  dp_1 \ANSWER/mem_reg[5][1][9]  ( .ip(n2883), .ck(clk), .q(
        \ANSWER/mem[5][1][9] ) );
  dp_1 \ANSWER/mem_reg[5][2][9]  ( .ip(n2882), .ck(clk), .q(
        \ANSWER/mem[5][2][9] ) );
  dp_1 \ANSWER/mem_reg[5][3][9]  ( .ip(n2881), .ck(clk), .q(
        \ANSWER/mem[5][3][9] ) );
  dp_1 \ANSWER/mem_reg[5][4][9]  ( .ip(n2880), .ck(clk), .q(
        \ANSWER/mem[5][4][9] ) );
  dp_1 \ANSWER/mem_reg[5][5][9]  ( .ip(n2879), .ck(clk), .q(
        \ANSWER/mem[5][5][9] ) );
  dp_1 \ANSWER/mem_reg[5][6][9]  ( .ip(n2878), .ck(clk), .q(
        \ANSWER/mem[5][6][9] ) );
  dp_1 \ANSWER/mem_reg[5][7][9]  ( .ip(n2877), .ck(clk), .q(
        \ANSWER/mem[5][7][9] ) );
  dp_1 \ANSWER/mem_reg[5][8][9]  ( .ip(n2876), .ck(clk), .q(
        \ANSWER/mem[5][8][9] ) );
  dp_1 \ANSWER/mem_reg[5][9][9]  ( .ip(n2875), .ck(clk), .q(
        \ANSWER/mem[5][9][9] ) );
  dp_1 \ANSWER/mem_reg[6][0][9]  ( .ip(n2874), .ck(clk), .q(
        \ANSWER/mem[6][0][9] ) );
  dp_1 \ANSWER/mem_reg[6][1][9]  ( .ip(n2873), .ck(clk), .q(
        \ANSWER/mem[6][1][9] ) );
  dp_1 \ANSWER/mem_reg[6][2][9]  ( .ip(n2872), .ck(clk), .q(
        \ANSWER/mem[6][2][9] ) );
  dp_1 \ANSWER/mem_reg[6][3][9]  ( .ip(n2871), .ck(clk), .q(
        \ANSWER/mem[6][3][9] ) );
  dp_1 \ANSWER/mem_reg[6][4][9]  ( .ip(n2870), .ck(clk), .q(
        \ANSWER/mem[6][4][9] ) );
  dp_1 \ANSWER/mem_reg[6][5][9]  ( .ip(n2869), .ck(clk), .q(
        \ANSWER/mem[6][5][9] ) );
  dp_1 \ANSWER/mem_reg[6][6][9]  ( .ip(n2868), .ck(clk), .q(
        \ANSWER/mem[6][6][9] ) );
  dp_1 \ANSWER/mem_reg[6][7][9]  ( .ip(n2867), .ck(clk), .q(
        \ANSWER/mem[6][7][9] ) );
  dp_1 \ANSWER/mem_reg[6][8][9]  ( .ip(n2866), .ck(clk), .q(
        \ANSWER/mem[6][8][9] ) );
  dp_1 \ANSWER/mem_reg[6][9][9]  ( .ip(n2865), .ck(clk), .q(
        \ANSWER/mem[6][9][9] ) );
  dp_1 \ANSWER/mem_reg[7][0][9]  ( .ip(n2864), .ck(clk), .q(
        \ANSWER/mem[7][0][9] ) );
  dp_1 \ANSWER/mem_reg[7][1][9]  ( .ip(n2863), .ck(clk), .q(
        \ANSWER/mem[7][1][9] ) );
  dp_1 \ANSWER/mem_reg[7][2][9]  ( .ip(n2862), .ck(clk), .q(
        \ANSWER/mem[7][2][9] ) );
  dp_1 \ANSWER/mem_reg[7][3][9]  ( .ip(n2861), .ck(clk), .q(
        \ANSWER/mem[7][3][9] ) );
  dp_1 \ANSWER/mem_reg[7][4][9]  ( .ip(n2860), .ck(clk), .q(
        \ANSWER/mem[7][4][9] ) );
  dp_1 \ANSWER/mem_reg[7][5][9]  ( .ip(n2859), .ck(clk), .q(
        \ANSWER/mem[7][5][9] ) );
  dp_1 \ANSWER/mem_reg[7][6][9]  ( .ip(n2858), .ck(clk), .q(
        \ANSWER/mem[7][6][9] ) );
  dp_1 \ANSWER/mem_reg[7][7][9]  ( .ip(n2857), .ck(clk), .q(
        \ANSWER/mem[7][7][9] ) );
  dp_1 \ANSWER/mem_reg[7][8][9]  ( .ip(n2856), .ck(clk), .q(
        \ANSWER/mem[7][8][9] ) );
  dp_1 \ANSWER/mem_reg[7][9][9]  ( .ip(n2855), .ck(clk), .q(
        \ANSWER/mem[7][9][9] ) );
  dp_1 \ANSWER/mem_reg[8][0][9]  ( .ip(n2854), .ck(clk), .q(
        \ANSWER/mem[8][0][9] ) );
  dp_1 \ANSWER/mem_reg[8][1][9]  ( .ip(n2853), .ck(clk), .q(
        \ANSWER/mem[8][1][9] ) );
  dp_1 \ANSWER/mem_reg[8][2][9]  ( .ip(n2852), .ck(clk), .q(
        \ANSWER/mem[8][2][9] ) );
  dp_1 \ANSWER/mem_reg[8][3][9]  ( .ip(n2851), .ck(clk), .q(
        \ANSWER/mem[8][3][9] ) );
  dp_1 \ANSWER/mem_reg[8][4][9]  ( .ip(n2850), .ck(clk), .q(
        \ANSWER/mem[8][4][9] ) );
  dp_1 \ANSWER/mem_reg[8][5][9]  ( .ip(n2849), .ck(clk), .q(
        \ANSWER/mem[8][5][9] ) );
  dp_1 \ANSWER/mem_reg[8][6][9]  ( .ip(n2848), .ck(clk), .q(
        \ANSWER/mem[8][6][9] ) );
  dp_1 \ANSWER/mem_reg[8][7][9]  ( .ip(n2847), .ck(clk), .q(
        \ANSWER/mem[8][7][9] ) );
  dp_1 \ANSWER/mem_reg[8][8][9]  ( .ip(n2846), .ck(clk), .q(
        \ANSWER/mem[8][8][9] ) );
  dp_1 \ANSWER/mem_reg[8][9][9]  ( .ip(n2845), .ck(clk), .q(
        \ANSWER/mem[8][9][9] ) );
  dp_1 \ANSWER/mem_reg[9][0][9]  ( .ip(n2844), .ck(clk), .q(
        \ANSWER/mem[9][0][9] ) );
  dp_1 \ANSWER/mem_reg[9][1][9]  ( .ip(n2843), .ck(clk), .q(
        \ANSWER/mem[9][1][9] ) );
  dp_1 \ANSWER/mem_reg[9][2][9]  ( .ip(n2842), .ck(clk), .q(
        \ANSWER/mem[9][2][9] ) );
  dp_1 \ANSWER/mem_reg[9][3][9]  ( .ip(n2841), .ck(clk), .q(
        \ANSWER/mem[9][3][9] ) );
  dp_1 \ANSWER/mem_reg[9][4][9]  ( .ip(n2840), .ck(clk), .q(
        \ANSWER/mem[9][4][9] ) );
  dp_1 \ANSWER/mem_reg[9][5][9]  ( .ip(n2839), .ck(clk), .q(
        \ANSWER/mem[9][5][9] ) );
  dp_1 \ANSWER/mem_reg[9][6][9]  ( .ip(n2838), .ck(clk), .q(
        \ANSWER/mem[9][6][9] ) );
  dp_1 \ANSWER/mem_reg[9][7][9]  ( .ip(n2837), .ck(clk), .q(
        \ANSWER/mem[9][7][9] ) );
  dp_1 \ANSWER/mem_reg[9][8][9]  ( .ip(n2836), .ck(clk), .q(
        \ANSWER/mem[9][8][9] ) );
  dp_1 \ANSWER/mem_reg[9][9][9]  ( .ip(n2835), .ck(clk), .q(
        \ANSWER/mem[9][9][9] ) );
  dp_1 \ANSWER/mem_reg[0][0][10]  ( .ip(n2834), .ck(clk), .q(
        \ANSWER/mem[0][0][10] ) );
  dp_1 \ANSWER/mem_reg[0][1][10]  ( .ip(n2833), .ck(clk), .q(
        \ANSWER/mem[0][1][10] ) );
  dp_1 \ANSWER/mem_reg[0][2][10]  ( .ip(n2832), .ck(clk), .q(
        \ANSWER/mem[0][2][10] ) );
  dp_1 \ANSWER/mem_reg[0][3][10]  ( .ip(n2831), .ck(clk), .q(
        \ANSWER/mem[0][3][10] ) );
  dp_1 \ANSWER/mem_reg[0][4][10]  ( .ip(n2830), .ck(clk), .q(
        \ANSWER/mem[0][4][10] ) );
  dp_1 \ANSWER/mem_reg[0][5][10]  ( .ip(n2829), .ck(clk), .q(
        \ANSWER/mem[0][5][10] ) );
  dp_1 \ANSWER/mem_reg[0][6][10]  ( .ip(n2828), .ck(clk), .q(
        \ANSWER/mem[0][6][10] ) );
  dp_1 \ANSWER/mem_reg[0][7][10]  ( .ip(n2827), .ck(clk), .q(
        \ANSWER/mem[0][7][10] ) );
  dp_1 \ANSWER/mem_reg[0][8][10]  ( .ip(n2826), .ck(clk), .q(
        \ANSWER/mem[0][8][10] ) );
  dp_1 \ANSWER/mem_reg[0][9][10]  ( .ip(n2825), .ck(clk), .q(
        \ANSWER/mem[0][9][10] ) );
  dp_1 \ANSWER/mem_reg[1][0][10]  ( .ip(n2824), .ck(clk), .q(
        \ANSWER/mem[1][0][10] ) );
  dp_1 \ANSWER/mem_reg[1][1][10]  ( .ip(n2823), .ck(clk), .q(
        \ANSWER/mem[1][1][10] ) );
  dp_1 \ANSWER/mem_reg[1][2][10]  ( .ip(n2822), .ck(clk), .q(
        \ANSWER/mem[1][2][10] ) );
  dp_1 \ANSWER/mem_reg[1][3][10]  ( .ip(n2821), .ck(clk), .q(
        \ANSWER/mem[1][3][10] ) );
  dp_1 \ANSWER/mem_reg[1][4][10]  ( .ip(n2820), .ck(clk), .q(
        \ANSWER/mem[1][4][10] ) );
  dp_1 \ANSWER/mem_reg[1][5][10]  ( .ip(n2819), .ck(clk), .q(
        \ANSWER/mem[1][5][10] ) );
  dp_1 \ANSWER/mem_reg[1][6][10]  ( .ip(n2818), .ck(clk), .q(
        \ANSWER/mem[1][6][10] ) );
  dp_1 \ANSWER/mem_reg[1][7][10]  ( .ip(n2817), .ck(clk), .q(
        \ANSWER/mem[1][7][10] ) );
  dp_1 \ANSWER/mem_reg[1][8][10]  ( .ip(n2816), .ck(clk), .q(
        \ANSWER/mem[1][8][10] ) );
  dp_1 \ANSWER/mem_reg[1][9][10]  ( .ip(n2815), .ck(clk), .q(
        \ANSWER/mem[1][9][10] ) );
  dp_1 \ANSWER/mem_reg[2][0][10]  ( .ip(n2814), .ck(clk), .q(
        \ANSWER/mem[2][0][10] ) );
  dp_1 \ANSWER/mem_reg[2][1][10]  ( .ip(n2813), .ck(clk), .q(
        \ANSWER/mem[2][1][10] ) );
  dp_1 \ANSWER/mem_reg[2][2][10]  ( .ip(n2812), .ck(clk), .q(
        \ANSWER/mem[2][2][10] ) );
  dp_1 \ANSWER/mem_reg[2][3][10]  ( .ip(n2811), .ck(clk), .q(
        \ANSWER/mem[2][3][10] ) );
  dp_1 \ANSWER/mem_reg[2][4][10]  ( .ip(n2810), .ck(clk), .q(
        \ANSWER/mem[2][4][10] ) );
  dp_1 \ANSWER/mem_reg[2][5][10]  ( .ip(n2809), .ck(clk), .q(
        \ANSWER/mem[2][5][10] ) );
  dp_1 \ANSWER/mem_reg[2][6][10]  ( .ip(n2808), .ck(clk), .q(
        \ANSWER/mem[2][6][10] ) );
  dp_1 \ANSWER/mem_reg[2][7][10]  ( .ip(n2807), .ck(clk), .q(
        \ANSWER/mem[2][7][10] ) );
  dp_1 \ANSWER/mem_reg[2][8][10]  ( .ip(n2806), .ck(clk), .q(
        \ANSWER/mem[2][8][10] ) );
  dp_1 \ANSWER/mem_reg[2][9][10]  ( .ip(n2805), .ck(clk), .q(
        \ANSWER/mem[2][9][10] ) );
  dp_1 \ANSWER/mem_reg[3][0][10]  ( .ip(n2804), .ck(clk), .q(
        \ANSWER/mem[3][0][10] ) );
  dp_1 \ANSWER/mem_reg[3][1][10]  ( .ip(n2803), .ck(clk), .q(
        \ANSWER/mem[3][1][10] ) );
  dp_1 \ANSWER/mem_reg[3][2][10]  ( .ip(n2802), .ck(clk), .q(
        \ANSWER/mem[3][2][10] ) );
  dp_1 \ANSWER/mem_reg[3][3][10]  ( .ip(n2801), .ck(clk), .q(
        \ANSWER/mem[3][3][10] ) );
  dp_1 \ANSWER/mem_reg[3][4][10]  ( .ip(n2800), .ck(clk), .q(
        \ANSWER/mem[3][4][10] ) );
  dp_1 \ANSWER/mem_reg[3][5][10]  ( .ip(n2799), .ck(clk), .q(
        \ANSWER/mem[3][5][10] ) );
  dp_1 \ANSWER/mem_reg[3][6][10]  ( .ip(n2798), .ck(clk), .q(
        \ANSWER/mem[3][6][10] ) );
  dp_1 \ANSWER/mem_reg[3][7][10]  ( .ip(n2797), .ck(clk), .q(
        \ANSWER/mem[3][7][10] ) );
  dp_1 \ANSWER/mem_reg[3][8][10]  ( .ip(n2796), .ck(clk), .q(
        \ANSWER/mem[3][8][10] ) );
  dp_1 \ANSWER/mem_reg[3][9][10]  ( .ip(n2795), .ck(clk), .q(
        \ANSWER/mem[3][9][10] ) );
  dp_1 \ANSWER/mem_reg[4][0][10]  ( .ip(n2794), .ck(clk), .q(
        \ANSWER/mem[4][0][10] ) );
  dp_1 \ANSWER/mem_reg[4][1][10]  ( .ip(n2793), .ck(clk), .q(
        \ANSWER/mem[4][1][10] ) );
  dp_1 \ANSWER/mem_reg[4][2][10]  ( .ip(n2792), .ck(clk), .q(
        \ANSWER/mem[4][2][10] ) );
  dp_1 \ANSWER/mem_reg[4][3][10]  ( .ip(n2791), .ck(clk), .q(
        \ANSWER/mem[4][3][10] ) );
  dp_1 \ANSWER/mem_reg[4][4][10]  ( .ip(n2790), .ck(clk), .q(
        \ANSWER/mem[4][4][10] ) );
  dp_1 \ANSWER/mem_reg[4][5][10]  ( .ip(n2789), .ck(clk), .q(
        \ANSWER/mem[4][5][10] ) );
  dp_1 \ANSWER/mem_reg[4][6][10]  ( .ip(n2788), .ck(clk), .q(
        \ANSWER/mem[4][6][10] ) );
  dp_1 \ANSWER/mem_reg[4][7][10]  ( .ip(n2787), .ck(clk), .q(
        \ANSWER/mem[4][7][10] ) );
  dp_1 \ANSWER/mem_reg[4][8][10]  ( .ip(n2786), .ck(clk), .q(
        \ANSWER/mem[4][8][10] ) );
  dp_1 \ANSWER/mem_reg[4][9][10]  ( .ip(n2785), .ck(clk), .q(
        \ANSWER/mem[4][9][10] ) );
  dp_1 \ANSWER/mem_reg[5][0][10]  ( .ip(n2784), .ck(clk), .q(
        \ANSWER/mem[5][0][10] ) );
  dp_1 \ANSWER/mem_reg[5][1][10]  ( .ip(n2783), .ck(clk), .q(
        \ANSWER/mem[5][1][10] ) );
  dp_1 \ANSWER/mem_reg[5][2][10]  ( .ip(n2782), .ck(clk), .q(
        \ANSWER/mem[5][2][10] ) );
  dp_1 \ANSWER/mem_reg[5][3][10]  ( .ip(n2781), .ck(clk), .q(
        \ANSWER/mem[5][3][10] ) );
  dp_1 \ANSWER/mem_reg[5][4][10]  ( .ip(n2780), .ck(clk), .q(
        \ANSWER/mem[5][4][10] ) );
  dp_1 \ANSWER/mem_reg[5][5][10]  ( .ip(n2779), .ck(clk), .q(
        \ANSWER/mem[5][5][10] ) );
  dp_1 \ANSWER/mem_reg[5][6][10]  ( .ip(n2778), .ck(clk), .q(
        \ANSWER/mem[5][6][10] ) );
  dp_1 \ANSWER/mem_reg[5][7][10]  ( .ip(n2777), .ck(clk), .q(
        \ANSWER/mem[5][7][10] ) );
  dp_1 \ANSWER/mem_reg[5][8][10]  ( .ip(n2776), .ck(clk), .q(
        \ANSWER/mem[5][8][10] ) );
  dp_1 \ANSWER/mem_reg[5][9][10]  ( .ip(n2775), .ck(clk), .q(
        \ANSWER/mem[5][9][10] ) );
  dp_1 \ANSWER/mem_reg[6][0][10]  ( .ip(n2774), .ck(clk), .q(
        \ANSWER/mem[6][0][10] ) );
  dp_1 \ANSWER/mem_reg[6][1][10]  ( .ip(n2773), .ck(clk), .q(
        \ANSWER/mem[6][1][10] ) );
  dp_1 \ANSWER/mem_reg[6][2][10]  ( .ip(n2772), .ck(clk), .q(
        \ANSWER/mem[6][2][10] ) );
  dp_1 \ANSWER/mem_reg[6][3][10]  ( .ip(n2771), .ck(clk), .q(
        \ANSWER/mem[6][3][10] ) );
  dp_1 \ANSWER/mem_reg[6][4][10]  ( .ip(n2770), .ck(clk), .q(
        \ANSWER/mem[6][4][10] ) );
  dp_1 \ANSWER/mem_reg[6][5][10]  ( .ip(n2769), .ck(clk), .q(
        \ANSWER/mem[6][5][10] ) );
  dp_1 \ANSWER/mem_reg[6][6][10]  ( .ip(n2768), .ck(clk), .q(
        \ANSWER/mem[6][6][10] ) );
  dp_1 \ANSWER/mem_reg[6][7][10]  ( .ip(n2767), .ck(clk), .q(
        \ANSWER/mem[6][7][10] ) );
  dp_1 \ANSWER/mem_reg[6][8][10]  ( .ip(n2766), .ck(clk), .q(
        \ANSWER/mem[6][8][10] ) );
  dp_1 \ANSWER/mem_reg[6][9][10]  ( .ip(n2765), .ck(clk), .q(
        \ANSWER/mem[6][9][10] ) );
  dp_1 \ANSWER/mem_reg[7][0][10]  ( .ip(n2764), .ck(clk), .q(
        \ANSWER/mem[7][0][10] ) );
  dp_1 \ANSWER/mem_reg[7][1][10]  ( .ip(n2763), .ck(clk), .q(
        \ANSWER/mem[7][1][10] ) );
  dp_1 \ANSWER/mem_reg[7][2][10]  ( .ip(n2762), .ck(clk), .q(
        \ANSWER/mem[7][2][10] ) );
  dp_1 \ANSWER/mem_reg[7][3][10]  ( .ip(n2761), .ck(clk), .q(
        \ANSWER/mem[7][3][10] ) );
  dp_1 \ANSWER/mem_reg[7][4][10]  ( .ip(n2760), .ck(clk), .q(
        \ANSWER/mem[7][4][10] ) );
  dp_1 \ANSWER/mem_reg[7][5][10]  ( .ip(n2759), .ck(clk), .q(
        \ANSWER/mem[7][5][10] ) );
  dp_1 \ANSWER/mem_reg[7][6][10]  ( .ip(n2758), .ck(clk), .q(
        \ANSWER/mem[7][6][10] ) );
  dp_1 \ANSWER/mem_reg[7][7][10]  ( .ip(n2757), .ck(clk), .q(
        \ANSWER/mem[7][7][10] ) );
  dp_1 \ANSWER/mem_reg[7][8][10]  ( .ip(n2756), .ck(clk), .q(
        \ANSWER/mem[7][8][10] ) );
  dp_1 \ANSWER/mem_reg[7][9][10]  ( .ip(n2755), .ck(clk), .q(
        \ANSWER/mem[7][9][10] ) );
  dp_1 \ANSWER/mem_reg[8][0][10]  ( .ip(n2754), .ck(clk), .q(
        \ANSWER/mem[8][0][10] ) );
  dp_1 \ANSWER/mem_reg[8][1][10]  ( .ip(n2753), .ck(clk), .q(
        \ANSWER/mem[8][1][10] ) );
  dp_1 \ANSWER/mem_reg[8][2][10]  ( .ip(n2752), .ck(clk), .q(
        \ANSWER/mem[8][2][10] ) );
  dp_1 \ANSWER/mem_reg[8][3][10]  ( .ip(n2751), .ck(clk), .q(
        \ANSWER/mem[8][3][10] ) );
  dp_1 \ANSWER/mem_reg[8][4][10]  ( .ip(n2750), .ck(clk), .q(
        \ANSWER/mem[8][4][10] ) );
  dp_1 \ANSWER/mem_reg[8][5][10]  ( .ip(n2749), .ck(clk), .q(
        \ANSWER/mem[8][5][10] ) );
  dp_1 \ANSWER/mem_reg[8][6][10]  ( .ip(n2748), .ck(clk), .q(
        \ANSWER/mem[8][6][10] ) );
  dp_1 \ANSWER/mem_reg[8][7][10]  ( .ip(n2747), .ck(clk), .q(
        \ANSWER/mem[8][7][10] ) );
  dp_1 \ANSWER/mem_reg[8][8][10]  ( .ip(n2746), .ck(clk), .q(
        \ANSWER/mem[8][8][10] ) );
  dp_1 \ANSWER/mem_reg[8][9][10]  ( .ip(n2745), .ck(clk), .q(
        \ANSWER/mem[8][9][10] ) );
  dp_1 \ANSWER/mem_reg[9][0][10]  ( .ip(n2744), .ck(clk), .q(
        \ANSWER/mem[9][0][10] ) );
  dp_1 \ANSWER/mem_reg[9][1][10]  ( .ip(n2743), .ck(clk), .q(
        \ANSWER/mem[9][1][10] ) );
  dp_1 \ANSWER/mem_reg[9][2][10]  ( .ip(n2742), .ck(clk), .q(
        \ANSWER/mem[9][2][10] ) );
  dp_1 \ANSWER/mem_reg[9][3][10]  ( .ip(n2741), .ck(clk), .q(
        \ANSWER/mem[9][3][10] ) );
  dp_1 \ANSWER/mem_reg[9][4][10]  ( .ip(n2740), .ck(clk), .q(
        \ANSWER/mem[9][4][10] ) );
  dp_1 \ANSWER/mem_reg[9][5][10]  ( .ip(n2739), .ck(clk), .q(
        \ANSWER/mem[9][5][10] ) );
  dp_1 \ANSWER/mem_reg[9][6][10]  ( .ip(n2738), .ck(clk), .q(
        \ANSWER/mem[9][6][10] ) );
  dp_1 \ANSWER/mem_reg[9][7][10]  ( .ip(n2737), .ck(clk), .q(
        \ANSWER/mem[9][7][10] ) );
  dp_1 \ANSWER/mem_reg[9][8][10]  ( .ip(n2736), .ck(clk), .q(
        \ANSWER/mem[9][8][10] ) );
  dp_1 \ANSWER/mem_reg[9][9][10]  ( .ip(n2735), .ck(clk), .q(
        \ANSWER/mem[9][9][10] ) );
  dp_1 \ANSWER/mem_reg[0][0][11]  ( .ip(n2734), .ck(clk), .q(
        \ANSWER/mem[0][0][11] ) );
  dp_1 \ANSWER/mem_reg[0][1][11]  ( .ip(n2733), .ck(clk), .q(
        \ANSWER/mem[0][1][11] ) );
  dp_1 \ANSWER/mem_reg[0][2][11]  ( .ip(n2732), .ck(clk), .q(
        \ANSWER/mem[0][2][11] ) );
  dp_1 \ANSWER/mem_reg[0][3][11]  ( .ip(n2731), .ck(clk), .q(
        \ANSWER/mem[0][3][11] ) );
  dp_1 \ANSWER/mem_reg[0][4][11]  ( .ip(n2730), .ck(clk), .q(
        \ANSWER/mem[0][4][11] ) );
  dp_1 \ANSWER/mem_reg[0][5][11]  ( .ip(n2729), .ck(clk), .q(
        \ANSWER/mem[0][5][11] ) );
  dp_1 \ANSWER/mem_reg[0][6][11]  ( .ip(n2728), .ck(clk), .q(
        \ANSWER/mem[0][6][11] ) );
  dp_1 \ANSWER/mem_reg[0][7][11]  ( .ip(n2727), .ck(clk), .q(
        \ANSWER/mem[0][7][11] ) );
  dp_1 \ANSWER/mem_reg[0][8][11]  ( .ip(n2726), .ck(clk), .q(
        \ANSWER/mem[0][8][11] ) );
  dp_1 \ANSWER/mem_reg[0][9][11]  ( .ip(n2725), .ck(clk), .q(
        \ANSWER/mem[0][9][11] ) );
  dp_1 \ANSWER/mem_reg[1][0][11]  ( .ip(n2724), .ck(clk), .q(
        \ANSWER/mem[1][0][11] ) );
  dp_1 \ANSWER/mem_reg[1][1][11]  ( .ip(n2723), .ck(clk), .q(
        \ANSWER/mem[1][1][11] ) );
  dp_1 \ANSWER/mem_reg[1][2][11]  ( .ip(n2722), .ck(clk), .q(
        \ANSWER/mem[1][2][11] ) );
  dp_1 \ANSWER/mem_reg[1][3][11]  ( .ip(n2721), .ck(clk), .q(
        \ANSWER/mem[1][3][11] ) );
  dp_1 \ANSWER/mem_reg[1][4][11]  ( .ip(n2720), .ck(clk), .q(
        \ANSWER/mem[1][4][11] ) );
  dp_1 \ANSWER/mem_reg[1][5][11]  ( .ip(n2719), .ck(clk), .q(
        \ANSWER/mem[1][5][11] ) );
  dp_1 \ANSWER/mem_reg[1][6][11]  ( .ip(n2718), .ck(clk), .q(
        \ANSWER/mem[1][6][11] ) );
  dp_1 \ANSWER/mem_reg[1][7][11]  ( .ip(n2717), .ck(clk), .q(
        \ANSWER/mem[1][7][11] ) );
  dp_1 \ANSWER/mem_reg[1][8][11]  ( .ip(n2716), .ck(clk), .q(
        \ANSWER/mem[1][8][11] ) );
  dp_1 \ANSWER/mem_reg[1][9][11]  ( .ip(n2715), .ck(clk), .q(
        \ANSWER/mem[1][9][11] ) );
  dp_1 \ANSWER/mem_reg[2][0][11]  ( .ip(n2714), .ck(clk), .q(
        \ANSWER/mem[2][0][11] ) );
  dp_1 \ANSWER/mem_reg[2][1][11]  ( .ip(n2713), .ck(clk), .q(
        \ANSWER/mem[2][1][11] ) );
  dp_1 \ANSWER/mem_reg[2][2][11]  ( .ip(n2712), .ck(clk), .q(
        \ANSWER/mem[2][2][11] ) );
  dp_1 \ANSWER/mem_reg[2][3][11]  ( .ip(n2711), .ck(clk), .q(
        \ANSWER/mem[2][3][11] ) );
  dp_1 \ANSWER/mem_reg[2][4][11]  ( .ip(n2710), .ck(clk), .q(
        \ANSWER/mem[2][4][11] ) );
  dp_1 \ANSWER/mem_reg[2][5][11]  ( .ip(n2709), .ck(clk), .q(
        \ANSWER/mem[2][5][11] ) );
  dp_1 \ANSWER/mem_reg[2][6][11]  ( .ip(n2708), .ck(clk), .q(
        \ANSWER/mem[2][6][11] ) );
  dp_1 \ANSWER/mem_reg[2][7][11]  ( .ip(n2707), .ck(clk), .q(
        \ANSWER/mem[2][7][11] ) );
  dp_1 \ANSWER/mem_reg[2][8][11]  ( .ip(n2706), .ck(clk), .q(
        \ANSWER/mem[2][8][11] ) );
  dp_1 \ANSWER/mem_reg[2][9][11]  ( .ip(n2705), .ck(clk), .q(
        \ANSWER/mem[2][9][11] ) );
  dp_1 \ANSWER/mem_reg[3][0][11]  ( .ip(n2704), .ck(clk), .q(
        \ANSWER/mem[3][0][11] ) );
  dp_1 \ANSWER/mem_reg[3][1][11]  ( .ip(n2703), .ck(clk), .q(
        \ANSWER/mem[3][1][11] ) );
  dp_1 \ANSWER/mem_reg[3][2][11]  ( .ip(n2702), .ck(clk), .q(
        \ANSWER/mem[3][2][11] ) );
  dp_1 \ANSWER/mem_reg[3][3][11]  ( .ip(n2701), .ck(clk), .q(
        \ANSWER/mem[3][3][11] ) );
  dp_1 \ANSWER/mem_reg[3][4][11]  ( .ip(n2700), .ck(clk), .q(
        \ANSWER/mem[3][4][11] ) );
  dp_1 \ANSWER/mem_reg[3][5][11]  ( .ip(n2699), .ck(clk), .q(
        \ANSWER/mem[3][5][11] ) );
  dp_1 \ANSWER/mem_reg[3][6][11]  ( .ip(n2698), .ck(clk), .q(
        \ANSWER/mem[3][6][11] ) );
  dp_1 \ANSWER/mem_reg[3][7][11]  ( .ip(n2697), .ck(clk), .q(
        \ANSWER/mem[3][7][11] ) );
  dp_1 \ANSWER/mem_reg[3][8][11]  ( .ip(n2696), .ck(clk), .q(
        \ANSWER/mem[3][8][11] ) );
  dp_1 \ANSWER/mem_reg[3][9][11]  ( .ip(n2695), .ck(clk), .q(
        \ANSWER/mem[3][9][11] ) );
  dp_1 \ANSWER/mem_reg[4][0][11]  ( .ip(n2694), .ck(clk), .q(
        \ANSWER/mem[4][0][11] ) );
  dp_1 \ANSWER/mem_reg[4][1][11]  ( .ip(n2693), .ck(clk), .q(
        \ANSWER/mem[4][1][11] ) );
  dp_1 \ANSWER/mem_reg[4][2][11]  ( .ip(n2692), .ck(clk), .q(
        \ANSWER/mem[4][2][11] ) );
  dp_1 \ANSWER/mem_reg[4][3][11]  ( .ip(n2691), .ck(clk), .q(
        \ANSWER/mem[4][3][11] ) );
  dp_1 \ANSWER/mem_reg[4][4][11]  ( .ip(n2690), .ck(clk), .q(
        \ANSWER/mem[4][4][11] ) );
  dp_1 \ANSWER/mem_reg[4][5][11]  ( .ip(n2689), .ck(clk), .q(
        \ANSWER/mem[4][5][11] ) );
  dp_1 \ANSWER/mem_reg[4][6][11]  ( .ip(n2688), .ck(clk), .q(
        \ANSWER/mem[4][6][11] ) );
  dp_1 \ANSWER/mem_reg[4][7][11]  ( .ip(n2687), .ck(clk), .q(
        \ANSWER/mem[4][7][11] ) );
  dp_1 \ANSWER/mem_reg[4][8][11]  ( .ip(n2686), .ck(clk), .q(
        \ANSWER/mem[4][8][11] ) );
  dp_1 \ANSWER/mem_reg[4][9][11]  ( .ip(n2685), .ck(clk), .q(
        \ANSWER/mem[4][9][11] ) );
  dp_1 \ANSWER/mem_reg[5][0][11]  ( .ip(n2684), .ck(clk), .q(
        \ANSWER/mem[5][0][11] ) );
  dp_1 \ANSWER/mem_reg[5][1][11]  ( .ip(n2683), .ck(clk), .q(
        \ANSWER/mem[5][1][11] ) );
  dp_1 \ANSWER/mem_reg[5][2][11]  ( .ip(n2682), .ck(clk), .q(
        \ANSWER/mem[5][2][11] ) );
  dp_1 \ANSWER/mem_reg[5][3][11]  ( .ip(n2681), .ck(clk), .q(
        \ANSWER/mem[5][3][11] ) );
  dp_1 \ANSWER/mem_reg[5][4][11]  ( .ip(n2680), .ck(clk), .q(
        \ANSWER/mem[5][4][11] ) );
  dp_1 \ANSWER/mem_reg[5][5][11]  ( .ip(n2679), .ck(clk), .q(
        \ANSWER/mem[5][5][11] ) );
  dp_1 \ANSWER/mem_reg[5][6][11]  ( .ip(n2678), .ck(clk), .q(
        \ANSWER/mem[5][6][11] ) );
  dp_1 \ANSWER/mem_reg[5][7][11]  ( .ip(n2677), .ck(clk), .q(
        \ANSWER/mem[5][7][11] ) );
  dp_1 \ANSWER/mem_reg[5][8][11]  ( .ip(n2676), .ck(clk), .q(
        \ANSWER/mem[5][8][11] ) );
  dp_1 \ANSWER/mem_reg[5][9][11]  ( .ip(n2675), .ck(clk), .q(
        \ANSWER/mem[5][9][11] ) );
  dp_1 \ANSWER/mem_reg[6][0][11]  ( .ip(n2674), .ck(clk), .q(
        \ANSWER/mem[6][0][11] ) );
  dp_1 \ANSWER/mem_reg[6][1][11]  ( .ip(n2673), .ck(clk), .q(
        \ANSWER/mem[6][1][11] ) );
  dp_1 \ANSWER/mem_reg[6][2][11]  ( .ip(n2672), .ck(clk), .q(
        \ANSWER/mem[6][2][11] ) );
  dp_1 \ANSWER/mem_reg[6][3][11]  ( .ip(n2671), .ck(clk), .q(
        \ANSWER/mem[6][3][11] ) );
  dp_1 \ANSWER/mem_reg[6][4][11]  ( .ip(n2670), .ck(clk), .q(
        \ANSWER/mem[6][4][11] ) );
  dp_1 \ANSWER/mem_reg[6][5][11]  ( .ip(n2669), .ck(clk), .q(
        \ANSWER/mem[6][5][11] ) );
  dp_1 \ANSWER/mem_reg[6][6][11]  ( .ip(n2668), .ck(clk), .q(
        \ANSWER/mem[6][6][11] ) );
  dp_1 \ANSWER/mem_reg[6][7][11]  ( .ip(n2667), .ck(clk), .q(
        \ANSWER/mem[6][7][11] ) );
  dp_1 \ANSWER/mem_reg[6][8][11]  ( .ip(n2666), .ck(clk), .q(
        \ANSWER/mem[6][8][11] ) );
  dp_1 \ANSWER/mem_reg[6][9][11]  ( .ip(n2665), .ck(clk), .q(
        \ANSWER/mem[6][9][11] ) );
  dp_1 \ANSWER/mem_reg[7][0][11]  ( .ip(n2664), .ck(clk), .q(
        \ANSWER/mem[7][0][11] ) );
  dp_1 \ANSWER/mem_reg[7][1][11]  ( .ip(n2663), .ck(clk), .q(
        \ANSWER/mem[7][1][11] ) );
  dp_1 \ANSWER/mem_reg[7][2][11]  ( .ip(n2662), .ck(clk), .q(
        \ANSWER/mem[7][2][11] ) );
  dp_1 \ANSWER/mem_reg[7][3][11]  ( .ip(n2661), .ck(clk), .q(
        \ANSWER/mem[7][3][11] ) );
  dp_1 \ANSWER/mem_reg[7][4][11]  ( .ip(n2660), .ck(clk), .q(
        \ANSWER/mem[7][4][11] ) );
  dp_1 \ANSWER/mem_reg[7][5][11]  ( .ip(n2659), .ck(clk), .q(
        \ANSWER/mem[7][5][11] ) );
  dp_1 \ANSWER/mem_reg[7][6][11]  ( .ip(n2658), .ck(clk), .q(
        \ANSWER/mem[7][6][11] ) );
  dp_1 \ANSWER/mem_reg[7][7][11]  ( .ip(n2657), .ck(clk), .q(
        \ANSWER/mem[7][7][11] ) );
  dp_1 \ANSWER/mem_reg[7][8][11]  ( .ip(n2656), .ck(clk), .q(
        \ANSWER/mem[7][8][11] ) );
  dp_1 \ANSWER/mem_reg[7][9][11]  ( .ip(n2655), .ck(clk), .q(
        \ANSWER/mem[7][9][11] ) );
  dp_1 \ANSWER/mem_reg[8][0][11]  ( .ip(n2654), .ck(clk), .q(
        \ANSWER/mem[8][0][11] ) );
  dp_1 \ANSWER/mem_reg[8][1][11]  ( .ip(n2653), .ck(clk), .q(
        \ANSWER/mem[8][1][11] ) );
  dp_1 \ANSWER/mem_reg[8][2][11]  ( .ip(n2652), .ck(clk), .q(
        \ANSWER/mem[8][2][11] ) );
  dp_1 \ANSWER/mem_reg[8][3][11]  ( .ip(n2651), .ck(clk), .q(
        \ANSWER/mem[8][3][11] ) );
  dp_1 \ANSWER/mem_reg[8][4][11]  ( .ip(n2650), .ck(clk), .q(
        \ANSWER/mem[8][4][11] ) );
  dp_1 \ANSWER/mem_reg[8][5][11]  ( .ip(n2649), .ck(clk), .q(
        \ANSWER/mem[8][5][11] ) );
  dp_1 \ANSWER/mem_reg[8][6][11]  ( .ip(n2648), .ck(clk), .q(
        \ANSWER/mem[8][6][11] ) );
  dp_1 \ANSWER/mem_reg[8][7][11]  ( .ip(n2647), .ck(clk), .q(
        \ANSWER/mem[8][7][11] ) );
  dp_1 \ANSWER/mem_reg[8][8][11]  ( .ip(n2646), .ck(clk), .q(
        \ANSWER/mem[8][8][11] ) );
  dp_1 \ANSWER/mem_reg[8][9][11]  ( .ip(n2645), .ck(clk), .q(
        \ANSWER/mem[8][9][11] ) );
  dp_1 \ANSWER/mem_reg[9][0][11]  ( .ip(n2644), .ck(clk), .q(
        \ANSWER/mem[9][0][11] ) );
  dp_1 \ANSWER/mem_reg[9][1][11]  ( .ip(n2643), .ck(clk), .q(
        \ANSWER/mem[9][1][11] ) );
  dp_1 \ANSWER/mem_reg[9][2][11]  ( .ip(n2642), .ck(clk), .q(
        \ANSWER/mem[9][2][11] ) );
  dp_1 \ANSWER/mem_reg[9][3][11]  ( .ip(n2641), .ck(clk), .q(
        \ANSWER/mem[9][3][11] ) );
  dp_1 \ANSWER/mem_reg[9][4][11]  ( .ip(n2640), .ck(clk), .q(
        \ANSWER/mem[9][4][11] ) );
  dp_1 \ANSWER/mem_reg[9][5][11]  ( .ip(n2639), .ck(clk), .q(
        \ANSWER/mem[9][5][11] ) );
  dp_1 \ANSWER/mem_reg[9][6][11]  ( .ip(n2638), .ck(clk), .q(
        \ANSWER/mem[9][6][11] ) );
  dp_1 \ANSWER/mem_reg[9][7][11]  ( .ip(n2637), .ck(clk), .q(
        \ANSWER/mem[9][7][11] ) );
  dp_1 \ANSWER/mem_reg[9][8][11]  ( .ip(n2636), .ck(clk), .q(
        \ANSWER/mem[9][8][11] ) );
  dp_1 \ANSWER/mem_reg[9][9][11]  ( .ip(n2635), .ck(clk), .q(
        \ANSWER/mem[9][9][11] ) );
  dp_1 \ANSWER/mem_reg[0][0][12]  ( .ip(n2634), .ck(clk), .q(
        \ANSWER/mem[0][0][12] ) );
  dp_1 \ANSWER/mem_reg[0][1][12]  ( .ip(n2633), .ck(clk), .q(
        \ANSWER/mem[0][1][12] ) );
  dp_1 \ANSWER/mem_reg[0][2][12]  ( .ip(n2632), .ck(clk), .q(
        \ANSWER/mem[0][2][12] ) );
  dp_1 \ANSWER/mem_reg[0][3][12]  ( .ip(n2631), .ck(clk), .q(
        \ANSWER/mem[0][3][12] ) );
  dp_1 \ANSWER/mem_reg[0][4][12]  ( .ip(n2630), .ck(clk), .q(
        \ANSWER/mem[0][4][12] ) );
  dp_1 \ANSWER/mem_reg[0][5][12]  ( .ip(n2629), .ck(clk), .q(
        \ANSWER/mem[0][5][12] ) );
  dp_1 \ANSWER/mem_reg[0][6][12]  ( .ip(n2628), .ck(clk), .q(
        \ANSWER/mem[0][6][12] ) );
  dp_1 \ANSWER/mem_reg[0][7][12]  ( .ip(n2627), .ck(clk), .q(
        \ANSWER/mem[0][7][12] ) );
  dp_1 \ANSWER/mem_reg[0][8][12]  ( .ip(n2626), .ck(clk), .q(
        \ANSWER/mem[0][8][12] ) );
  dp_1 \ANSWER/mem_reg[0][9][12]  ( .ip(n2625), .ck(clk), .q(
        \ANSWER/mem[0][9][12] ) );
  dp_1 \ANSWER/mem_reg[1][0][12]  ( .ip(n2624), .ck(clk), .q(
        \ANSWER/mem[1][0][12] ) );
  dp_1 \ANSWER/mem_reg[1][1][12]  ( .ip(n2623), .ck(clk), .q(
        \ANSWER/mem[1][1][12] ) );
  dp_1 \ANSWER/mem_reg[1][2][12]  ( .ip(n2622), .ck(clk), .q(
        \ANSWER/mem[1][2][12] ) );
  dp_1 \ANSWER/mem_reg[1][3][12]  ( .ip(n2621), .ck(clk), .q(
        \ANSWER/mem[1][3][12] ) );
  dp_1 \ANSWER/mem_reg[1][4][12]  ( .ip(n2620), .ck(clk), .q(
        \ANSWER/mem[1][4][12] ) );
  dp_1 \ANSWER/mem_reg[1][5][12]  ( .ip(n2619), .ck(clk), .q(
        \ANSWER/mem[1][5][12] ) );
  dp_1 \ANSWER/mem_reg[1][6][12]  ( .ip(n2618), .ck(clk), .q(
        \ANSWER/mem[1][6][12] ) );
  dp_1 \ANSWER/mem_reg[1][7][12]  ( .ip(n2617), .ck(clk), .q(
        \ANSWER/mem[1][7][12] ) );
  dp_1 \ANSWER/mem_reg[1][8][12]  ( .ip(n2616), .ck(clk), .q(
        \ANSWER/mem[1][8][12] ) );
  dp_1 \ANSWER/mem_reg[1][9][12]  ( .ip(n2615), .ck(clk), .q(
        \ANSWER/mem[1][9][12] ) );
  dp_1 \ANSWER/mem_reg[2][0][12]  ( .ip(n2614), .ck(clk), .q(
        \ANSWER/mem[2][0][12] ) );
  dp_1 \ANSWER/mem_reg[2][1][12]  ( .ip(n2613), .ck(clk), .q(
        \ANSWER/mem[2][1][12] ) );
  dp_1 \ANSWER/mem_reg[2][2][12]  ( .ip(n2612), .ck(clk), .q(
        \ANSWER/mem[2][2][12] ) );
  dp_1 \ANSWER/mem_reg[2][3][12]  ( .ip(n2611), .ck(clk), .q(
        \ANSWER/mem[2][3][12] ) );
  dp_1 \ANSWER/mem_reg[2][4][12]  ( .ip(n2610), .ck(clk), .q(
        \ANSWER/mem[2][4][12] ) );
  dp_1 \ANSWER/mem_reg[2][5][12]  ( .ip(n2609), .ck(clk), .q(
        \ANSWER/mem[2][5][12] ) );
  dp_1 \ANSWER/mem_reg[2][6][12]  ( .ip(n2608), .ck(clk), .q(
        \ANSWER/mem[2][6][12] ) );
  dp_1 \ANSWER/mem_reg[2][7][12]  ( .ip(n2607), .ck(clk), .q(
        \ANSWER/mem[2][7][12] ) );
  dp_1 \ANSWER/mem_reg[2][8][12]  ( .ip(n2606), .ck(clk), .q(
        \ANSWER/mem[2][8][12] ) );
  dp_1 \ANSWER/mem_reg[2][9][12]  ( .ip(n2605), .ck(clk), .q(
        \ANSWER/mem[2][9][12] ) );
  dp_1 \ANSWER/mem_reg[3][0][12]  ( .ip(n2604), .ck(clk), .q(
        \ANSWER/mem[3][0][12] ) );
  dp_1 \ANSWER/mem_reg[3][1][12]  ( .ip(n2603), .ck(clk), .q(
        \ANSWER/mem[3][1][12] ) );
  dp_1 \ANSWER/mem_reg[3][2][12]  ( .ip(n2602), .ck(clk), .q(
        \ANSWER/mem[3][2][12] ) );
  dp_1 \ANSWER/mem_reg[3][3][12]  ( .ip(n2601), .ck(clk), .q(
        \ANSWER/mem[3][3][12] ) );
  dp_1 \ANSWER/mem_reg[3][4][12]  ( .ip(n2600), .ck(clk), .q(
        \ANSWER/mem[3][4][12] ) );
  dp_1 \ANSWER/mem_reg[3][5][12]  ( .ip(n2599), .ck(clk), .q(
        \ANSWER/mem[3][5][12] ) );
  dp_1 \ANSWER/mem_reg[3][6][12]  ( .ip(n2598), .ck(clk), .q(
        \ANSWER/mem[3][6][12] ) );
  dp_1 \ANSWER/mem_reg[3][7][12]  ( .ip(n2597), .ck(clk), .q(
        \ANSWER/mem[3][7][12] ) );
  dp_1 \ANSWER/mem_reg[3][8][12]  ( .ip(n2596), .ck(clk), .q(
        \ANSWER/mem[3][8][12] ) );
  dp_1 \ANSWER/mem_reg[3][9][12]  ( .ip(n2595), .ck(clk), .q(
        \ANSWER/mem[3][9][12] ) );
  dp_1 \ANSWER/mem_reg[4][0][12]  ( .ip(n2594), .ck(clk), .q(
        \ANSWER/mem[4][0][12] ) );
  dp_1 \ANSWER/mem_reg[4][1][12]  ( .ip(n2593), .ck(clk), .q(
        \ANSWER/mem[4][1][12] ) );
  dp_1 \ANSWER/mem_reg[4][2][12]  ( .ip(n2592), .ck(clk), .q(
        \ANSWER/mem[4][2][12] ) );
  dp_1 \ANSWER/mem_reg[4][3][12]  ( .ip(n2591), .ck(clk), .q(
        \ANSWER/mem[4][3][12] ) );
  dp_1 \ANSWER/mem_reg[4][4][12]  ( .ip(n2590), .ck(clk), .q(
        \ANSWER/mem[4][4][12] ) );
  dp_1 \ANSWER/mem_reg[4][5][12]  ( .ip(n2589), .ck(clk), .q(
        \ANSWER/mem[4][5][12] ) );
  dp_1 \ANSWER/mem_reg[4][6][12]  ( .ip(n2588), .ck(clk), .q(
        \ANSWER/mem[4][6][12] ) );
  dp_1 \ANSWER/mem_reg[4][7][12]  ( .ip(n2587), .ck(clk), .q(
        \ANSWER/mem[4][7][12] ) );
  dp_1 \ANSWER/mem_reg[4][8][12]  ( .ip(n2586), .ck(clk), .q(
        \ANSWER/mem[4][8][12] ) );
  dp_1 \ANSWER/mem_reg[4][9][12]  ( .ip(n2585), .ck(clk), .q(
        \ANSWER/mem[4][9][12] ) );
  dp_1 \ANSWER/mem_reg[5][0][12]  ( .ip(n2584), .ck(clk), .q(
        \ANSWER/mem[5][0][12] ) );
  dp_1 \ANSWER/mem_reg[5][1][12]  ( .ip(n2583), .ck(clk), .q(
        \ANSWER/mem[5][1][12] ) );
  dp_1 \ANSWER/mem_reg[5][2][12]  ( .ip(n2582), .ck(clk), .q(
        \ANSWER/mem[5][2][12] ) );
  dp_1 \ANSWER/mem_reg[5][3][12]  ( .ip(n2581), .ck(clk), .q(
        \ANSWER/mem[5][3][12] ) );
  dp_1 \ANSWER/mem_reg[5][4][12]  ( .ip(n2580), .ck(clk), .q(
        \ANSWER/mem[5][4][12] ) );
  dp_1 \ANSWER/mem_reg[5][5][12]  ( .ip(n2579), .ck(clk), .q(
        \ANSWER/mem[5][5][12] ) );
  dp_1 \ANSWER/mem_reg[5][6][12]  ( .ip(n2578), .ck(clk), .q(
        \ANSWER/mem[5][6][12] ) );
  dp_1 \ANSWER/mem_reg[5][7][12]  ( .ip(n2577), .ck(clk), .q(
        \ANSWER/mem[5][7][12] ) );
  dp_1 \ANSWER/mem_reg[5][8][12]  ( .ip(n2576), .ck(clk), .q(
        \ANSWER/mem[5][8][12] ) );
  dp_1 \ANSWER/mem_reg[5][9][12]  ( .ip(n2575), .ck(clk), .q(
        \ANSWER/mem[5][9][12] ) );
  dp_1 \ANSWER/mem_reg[6][0][12]  ( .ip(n2574), .ck(clk), .q(
        \ANSWER/mem[6][0][12] ) );
  dp_1 \ANSWER/mem_reg[6][1][12]  ( .ip(n2573), .ck(clk), .q(
        \ANSWER/mem[6][1][12] ) );
  dp_1 \ANSWER/mem_reg[6][2][12]  ( .ip(n2572), .ck(clk), .q(
        \ANSWER/mem[6][2][12] ) );
  dp_1 \ANSWER/mem_reg[6][3][12]  ( .ip(n2571), .ck(clk), .q(
        \ANSWER/mem[6][3][12] ) );
  dp_1 \ANSWER/mem_reg[6][4][12]  ( .ip(n2570), .ck(clk), .q(
        \ANSWER/mem[6][4][12] ) );
  dp_1 \ANSWER/mem_reg[6][5][12]  ( .ip(n2569), .ck(clk), .q(
        \ANSWER/mem[6][5][12] ) );
  dp_1 \ANSWER/mem_reg[6][6][12]  ( .ip(n2568), .ck(clk), .q(
        \ANSWER/mem[6][6][12] ) );
  dp_1 \ANSWER/mem_reg[6][7][12]  ( .ip(n2567), .ck(clk), .q(
        \ANSWER/mem[6][7][12] ) );
  dp_1 \ANSWER/mem_reg[6][8][12]  ( .ip(n2566), .ck(clk), .q(
        \ANSWER/mem[6][8][12] ) );
  dp_1 \ANSWER/mem_reg[6][9][12]  ( .ip(n2565), .ck(clk), .q(
        \ANSWER/mem[6][9][12] ) );
  dp_1 \ANSWER/mem_reg[7][0][12]  ( .ip(n2564), .ck(clk), .q(
        \ANSWER/mem[7][0][12] ) );
  dp_1 \ANSWER/mem_reg[7][1][12]  ( .ip(n2563), .ck(clk), .q(
        \ANSWER/mem[7][1][12] ) );
  dp_1 \ANSWER/mem_reg[7][2][12]  ( .ip(n2562), .ck(clk), .q(
        \ANSWER/mem[7][2][12] ) );
  dp_1 \ANSWER/mem_reg[7][3][12]  ( .ip(n2561), .ck(clk), .q(
        \ANSWER/mem[7][3][12] ) );
  dp_1 \ANSWER/mem_reg[7][4][12]  ( .ip(n2560), .ck(clk), .q(
        \ANSWER/mem[7][4][12] ) );
  dp_1 \ANSWER/mem_reg[7][5][12]  ( .ip(n2559), .ck(clk), .q(
        \ANSWER/mem[7][5][12] ) );
  dp_1 \ANSWER/mem_reg[7][6][12]  ( .ip(n2558), .ck(clk), .q(
        \ANSWER/mem[7][6][12] ) );
  dp_1 \ANSWER/mem_reg[7][7][12]  ( .ip(n2557), .ck(clk), .q(
        \ANSWER/mem[7][7][12] ) );
  dp_1 \ANSWER/mem_reg[7][8][12]  ( .ip(n2556), .ck(clk), .q(
        \ANSWER/mem[7][8][12] ) );
  dp_1 \ANSWER/mem_reg[7][9][12]  ( .ip(n2555), .ck(clk), .q(
        \ANSWER/mem[7][9][12] ) );
  dp_1 \ANSWER/mem_reg[8][0][12]  ( .ip(n2554), .ck(clk), .q(
        \ANSWER/mem[8][0][12] ) );
  dp_1 \ANSWER/mem_reg[8][1][12]  ( .ip(n2553), .ck(clk), .q(
        \ANSWER/mem[8][1][12] ) );
  dp_1 \ANSWER/mem_reg[8][2][12]  ( .ip(n2552), .ck(clk), .q(
        \ANSWER/mem[8][2][12] ) );
  dp_1 \ANSWER/mem_reg[8][3][12]  ( .ip(n2551), .ck(clk), .q(
        \ANSWER/mem[8][3][12] ) );
  dp_1 \ANSWER/mem_reg[8][4][12]  ( .ip(n2550), .ck(clk), .q(
        \ANSWER/mem[8][4][12] ) );
  dp_1 \ANSWER/mem_reg[8][5][12]  ( .ip(n2549), .ck(clk), .q(
        \ANSWER/mem[8][5][12] ) );
  dp_1 \ANSWER/mem_reg[8][6][12]  ( .ip(n2548), .ck(clk), .q(
        \ANSWER/mem[8][6][12] ) );
  dp_1 \ANSWER/mem_reg[8][7][12]  ( .ip(n2547), .ck(clk), .q(
        \ANSWER/mem[8][7][12] ) );
  dp_1 \ANSWER/mem_reg[8][8][12]  ( .ip(n2546), .ck(clk), .q(
        \ANSWER/mem[8][8][12] ) );
  dp_1 \ANSWER/mem_reg[8][9][12]  ( .ip(n2545), .ck(clk), .q(
        \ANSWER/mem[8][9][12] ) );
  dp_1 \ANSWER/mem_reg[9][0][12]  ( .ip(n2544), .ck(clk), .q(
        \ANSWER/mem[9][0][12] ) );
  dp_1 \ANSWER/mem_reg[9][1][12]  ( .ip(n2543), .ck(clk), .q(
        \ANSWER/mem[9][1][12] ) );
  dp_1 \ANSWER/mem_reg[9][2][12]  ( .ip(n2542), .ck(clk), .q(
        \ANSWER/mem[9][2][12] ) );
  dp_1 \ANSWER/mem_reg[9][3][12]  ( .ip(n2541), .ck(clk), .q(
        \ANSWER/mem[9][3][12] ) );
  dp_1 \ANSWER/mem_reg[9][4][12]  ( .ip(n2540), .ck(clk), .q(
        \ANSWER/mem[9][4][12] ) );
  dp_1 \ANSWER/mem_reg[9][5][12]  ( .ip(n2539), .ck(clk), .q(
        \ANSWER/mem[9][5][12] ) );
  dp_1 \ANSWER/mem_reg[9][6][12]  ( .ip(n2538), .ck(clk), .q(
        \ANSWER/mem[9][6][12] ) );
  dp_1 \ANSWER/mem_reg[9][7][12]  ( .ip(n2537), .ck(clk), .q(
        \ANSWER/mem[9][7][12] ) );
  dp_1 \ANSWER/mem_reg[9][8][12]  ( .ip(n2536), .ck(clk), .q(
        \ANSWER/mem[9][8][12] ) );
  dp_1 \ANSWER/mem_reg[9][9][12]  ( .ip(n2535), .ck(clk), .q(
        \ANSWER/mem[9][9][12] ) );
  dp_1 \ANSWER/mem_reg[0][0][13]  ( .ip(n2534), .ck(clk), .q(
        \ANSWER/mem[0][0][13] ) );
  dp_1 \ANSWER/mem_reg[0][1][13]  ( .ip(n2533), .ck(clk), .q(
        \ANSWER/mem[0][1][13] ) );
  dp_1 \ANSWER/mem_reg[0][2][13]  ( .ip(n2532), .ck(clk), .q(
        \ANSWER/mem[0][2][13] ) );
  dp_1 \ANSWER/mem_reg[0][3][13]  ( .ip(n2531), .ck(clk), .q(
        \ANSWER/mem[0][3][13] ) );
  dp_1 \ANSWER/mem_reg[0][4][13]  ( .ip(n2530), .ck(clk), .q(
        \ANSWER/mem[0][4][13] ) );
  dp_1 \ANSWER/mem_reg[0][5][13]  ( .ip(n2529), .ck(clk), .q(
        \ANSWER/mem[0][5][13] ) );
  dp_1 \ANSWER/mem_reg[0][6][13]  ( .ip(n2528), .ck(clk), .q(
        \ANSWER/mem[0][6][13] ) );
  dp_1 \ANSWER/mem_reg[0][7][13]  ( .ip(n2527), .ck(clk), .q(
        \ANSWER/mem[0][7][13] ) );
  dp_1 \ANSWER/mem_reg[0][8][13]  ( .ip(n2526), .ck(clk), .q(
        \ANSWER/mem[0][8][13] ) );
  dp_1 \ANSWER/mem_reg[0][9][13]  ( .ip(n2525), .ck(clk), .q(
        \ANSWER/mem[0][9][13] ) );
  dp_1 \ANSWER/mem_reg[1][0][13]  ( .ip(n2524), .ck(clk), .q(
        \ANSWER/mem[1][0][13] ) );
  dp_1 \ANSWER/mem_reg[1][1][13]  ( .ip(n2523), .ck(clk), .q(
        \ANSWER/mem[1][1][13] ) );
  dp_1 \ANSWER/mem_reg[1][2][13]  ( .ip(n2522), .ck(clk), .q(
        \ANSWER/mem[1][2][13] ) );
  dp_1 \ANSWER/mem_reg[1][3][13]  ( .ip(n2521), .ck(clk), .q(
        \ANSWER/mem[1][3][13] ) );
  dp_1 \ANSWER/mem_reg[1][4][13]  ( .ip(n2520), .ck(clk), .q(
        \ANSWER/mem[1][4][13] ) );
  dp_1 \ANSWER/mem_reg[1][5][13]  ( .ip(n2519), .ck(clk), .q(
        \ANSWER/mem[1][5][13] ) );
  dp_1 \ANSWER/mem_reg[1][6][13]  ( .ip(n2518), .ck(clk), .q(
        \ANSWER/mem[1][6][13] ) );
  dp_1 \ANSWER/mem_reg[1][7][13]  ( .ip(n2517), .ck(clk), .q(
        \ANSWER/mem[1][7][13] ) );
  dp_1 \ANSWER/mem_reg[1][8][13]  ( .ip(n2516), .ck(clk), .q(
        \ANSWER/mem[1][8][13] ) );
  dp_1 \ANSWER/mem_reg[1][9][13]  ( .ip(n2515), .ck(clk), .q(
        \ANSWER/mem[1][9][13] ) );
  dp_1 \ANSWER/mem_reg[2][0][13]  ( .ip(n2514), .ck(clk), .q(
        \ANSWER/mem[2][0][13] ) );
  dp_1 \ANSWER/mem_reg[2][1][13]  ( .ip(n2513), .ck(clk), .q(
        \ANSWER/mem[2][1][13] ) );
  dp_1 \ANSWER/mem_reg[2][2][13]  ( .ip(n2512), .ck(clk), .q(
        \ANSWER/mem[2][2][13] ) );
  dp_1 \ANSWER/mem_reg[2][3][13]  ( .ip(n2511), .ck(clk), .q(
        \ANSWER/mem[2][3][13] ) );
  dp_1 \ANSWER/mem_reg[2][4][13]  ( .ip(n2510), .ck(clk), .q(
        \ANSWER/mem[2][4][13] ) );
  dp_1 \ANSWER/mem_reg[2][5][13]  ( .ip(n2509), .ck(clk), .q(
        \ANSWER/mem[2][5][13] ) );
  dp_1 \ANSWER/mem_reg[2][6][13]  ( .ip(n2508), .ck(clk), .q(
        \ANSWER/mem[2][6][13] ) );
  dp_1 \ANSWER/mem_reg[2][7][13]  ( .ip(n2507), .ck(clk), .q(
        \ANSWER/mem[2][7][13] ) );
  dp_1 \ANSWER/mem_reg[2][8][13]  ( .ip(n2506), .ck(clk), .q(
        \ANSWER/mem[2][8][13] ) );
  dp_1 \ANSWER/mem_reg[2][9][13]  ( .ip(n2505), .ck(clk), .q(
        \ANSWER/mem[2][9][13] ) );
  dp_1 \ANSWER/mem_reg[3][0][13]  ( .ip(n2504), .ck(clk), .q(
        \ANSWER/mem[3][0][13] ) );
  dp_1 \ANSWER/mem_reg[3][1][13]  ( .ip(n2503), .ck(clk), .q(
        \ANSWER/mem[3][1][13] ) );
  dp_1 \ANSWER/mem_reg[3][2][13]  ( .ip(n2502), .ck(clk), .q(
        \ANSWER/mem[3][2][13] ) );
  dp_1 \ANSWER/mem_reg[3][3][13]  ( .ip(n2501), .ck(clk), .q(
        \ANSWER/mem[3][3][13] ) );
  dp_1 \ANSWER/mem_reg[3][4][13]  ( .ip(n2500), .ck(clk), .q(
        \ANSWER/mem[3][4][13] ) );
  dp_1 \ANSWER/mem_reg[3][5][13]  ( .ip(n2499), .ck(clk), .q(
        \ANSWER/mem[3][5][13] ) );
  dp_1 \ANSWER/mem_reg[3][6][13]  ( .ip(n2498), .ck(clk), .q(
        \ANSWER/mem[3][6][13] ) );
  dp_1 \ANSWER/mem_reg[3][7][13]  ( .ip(n2497), .ck(clk), .q(
        \ANSWER/mem[3][7][13] ) );
  dp_1 \ANSWER/mem_reg[3][8][13]  ( .ip(n2496), .ck(clk), .q(
        \ANSWER/mem[3][8][13] ) );
  dp_1 \ANSWER/mem_reg[3][9][13]  ( .ip(n2495), .ck(clk), .q(
        \ANSWER/mem[3][9][13] ) );
  dp_1 \ANSWER/mem_reg[4][0][13]  ( .ip(n2494), .ck(clk), .q(
        \ANSWER/mem[4][0][13] ) );
  dp_1 \ANSWER/mem_reg[4][1][13]  ( .ip(n2493), .ck(clk), .q(
        \ANSWER/mem[4][1][13] ) );
  dp_1 \ANSWER/mem_reg[4][2][13]  ( .ip(n2492), .ck(clk), .q(
        \ANSWER/mem[4][2][13] ) );
  dp_1 \ANSWER/mem_reg[4][3][13]  ( .ip(n2491), .ck(clk), .q(
        \ANSWER/mem[4][3][13] ) );
  dp_1 \ANSWER/mem_reg[4][4][13]  ( .ip(n2490), .ck(clk), .q(
        \ANSWER/mem[4][4][13] ) );
  dp_1 \ANSWER/mem_reg[4][5][13]  ( .ip(n2489), .ck(clk), .q(
        \ANSWER/mem[4][5][13] ) );
  dp_1 \ANSWER/mem_reg[4][6][13]  ( .ip(n2488), .ck(clk), .q(
        \ANSWER/mem[4][6][13] ) );
  dp_1 \ANSWER/mem_reg[4][7][13]  ( .ip(n2487), .ck(clk), .q(
        \ANSWER/mem[4][7][13] ) );
  dp_1 \ANSWER/mem_reg[4][8][13]  ( .ip(n2486), .ck(clk), .q(
        \ANSWER/mem[4][8][13] ) );
  dp_1 \ANSWER/mem_reg[4][9][13]  ( .ip(n2485), .ck(clk), .q(
        \ANSWER/mem[4][9][13] ) );
  dp_1 \ANSWER/mem_reg[5][0][13]  ( .ip(n2484), .ck(clk), .q(
        \ANSWER/mem[5][0][13] ) );
  dp_1 \ANSWER/mem_reg[5][1][13]  ( .ip(n2483), .ck(clk), .q(
        \ANSWER/mem[5][1][13] ) );
  dp_1 \ANSWER/mem_reg[5][2][13]  ( .ip(n2482), .ck(clk), .q(
        \ANSWER/mem[5][2][13] ) );
  dp_1 \ANSWER/mem_reg[5][3][13]  ( .ip(n2481), .ck(clk), .q(
        \ANSWER/mem[5][3][13] ) );
  dp_1 \ANSWER/mem_reg[5][4][13]  ( .ip(n2480), .ck(clk), .q(
        \ANSWER/mem[5][4][13] ) );
  dp_1 \ANSWER/mem_reg[5][5][13]  ( .ip(n2479), .ck(clk), .q(
        \ANSWER/mem[5][5][13] ) );
  dp_1 \ANSWER/mem_reg[5][6][13]  ( .ip(n2478), .ck(clk), .q(
        \ANSWER/mem[5][6][13] ) );
  dp_1 \ANSWER/mem_reg[5][7][13]  ( .ip(n2477), .ck(clk), .q(
        \ANSWER/mem[5][7][13] ) );
  dp_1 \ANSWER/mem_reg[5][8][13]  ( .ip(n2476), .ck(clk), .q(
        \ANSWER/mem[5][8][13] ) );
  dp_1 \ANSWER/mem_reg[5][9][13]  ( .ip(n2475), .ck(clk), .q(
        \ANSWER/mem[5][9][13] ) );
  dp_1 \ANSWER/mem_reg[6][0][13]  ( .ip(n2474), .ck(clk), .q(
        \ANSWER/mem[6][0][13] ) );
  dp_1 \ANSWER/mem_reg[6][1][13]  ( .ip(n2473), .ck(clk), .q(
        \ANSWER/mem[6][1][13] ) );
  dp_1 \ANSWER/mem_reg[6][2][13]  ( .ip(n2472), .ck(clk), .q(
        \ANSWER/mem[6][2][13] ) );
  dp_1 \ANSWER/mem_reg[6][3][13]  ( .ip(n2471), .ck(clk), .q(
        \ANSWER/mem[6][3][13] ) );
  dp_1 \ANSWER/mem_reg[6][4][13]  ( .ip(n2470), .ck(clk), .q(
        \ANSWER/mem[6][4][13] ) );
  dp_1 \ANSWER/mem_reg[6][5][13]  ( .ip(n2469), .ck(clk), .q(
        \ANSWER/mem[6][5][13] ) );
  dp_1 \ANSWER/mem_reg[6][6][13]  ( .ip(n2468), .ck(clk), .q(
        \ANSWER/mem[6][6][13] ) );
  dp_1 \ANSWER/mem_reg[6][7][13]  ( .ip(n2467), .ck(clk), .q(
        \ANSWER/mem[6][7][13] ) );
  dp_1 \ANSWER/mem_reg[6][8][13]  ( .ip(n2466), .ck(clk), .q(
        \ANSWER/mem[6][8][13] ) );
  dp_1 \ANSWER/mem_reg[6][9][13]  ( .ip(n2465), .ck(clk), .q(
        \ANSWER/mem[6][9][13] ) );
  dp_1 \ANSWER/mem_reg[7][0][13]  ( .ip(n2464), .ck(clk), .q(
        \ANSWER/mem[7][0][13] ) );
  dp_1 \ANSWER/mem_reg[7][1][13]  ( .ip(n2463), .ck(clk), .q(
        \ANSWER/mem[7][1][13] ) );
  dp_1 \ANSWER/mem_reg[7][2][13]  ( .ip(n2462), .ck(clk), .q(
        \ANSWER/mem[7][2][13] ) );
  dp_1 \ANSWER/mem_reg[7][3][13]  ( .ip(n2461), .ck(clk), .q(
        \ANSWER/mem[7][3][13] ) );
  dp_1 \ANSWER/mem_reg[7][4][13]  ( .ip(n2460), .ck(clk), .q(
        \ANSWER/mem[7][4][13] ) );
  dp_1 \ANSWER/mem_reg[7][5][13]  ( .ip(n2459), .ck(clk), .q(
        \ANSWER/mem[7][5][13] ) );
  dp_1 \ANSWER/mem_reg[7][6][13]  ( .ip(n2458), .ck(clk), .q(
        \ANSWER/mem[7][6][13] ) );
  dp_1 \ANSWER/mem_reg[7][7][13]  ( .ip(n2457), .ck(clk), .q(
        \ANSWER/mem[7][7][13] ) );
  dp_1 \ANSWER/mem_reg[7][8][13]  ( .ip(n2456), .ck(clk), .q(
        \ANSWER/mem[7][8][13] ) );
  dp_1 \ANSWER/mem_reg[7][9][13]  ( .ip(n2455), .ck(clk), .q(
        \ANSWER/mem[7][9][13] ) );
  dp_1 \ANSWER/mem_reg[8][0][13]  ( .ip(n2454), .ck(clk), .q(
        \ANSWER/mem[8][0][13] ) );
  dp_1 \ANSWER/mem_reg[8][1][13]  ( .ip(n2453), .ck(clk), .q(
        \ANSWER/mem[8][1][13] ) );
  dp_1 \ANSWER/mem_reg[8][2][13]  ( .ip(n2452), .ck(clk), .q(
        \ANSWER/mem[8][2][13] ) );
  dp_1 \ANSWER/mem_reg[8][3][13]  ( .ip(n2451), .ck(clk), .q(
        \ANSWER/mem[8][3][13] ) );
  dp_1 \ANSWER/mem_reg[8][4][13]  ( .ip(n2450), .ck(clk), .q(
        \ANSWER/mem[8][4][13] ) );
  dp_1 \ANSWER/mem_reg[8][5][13]  ( .ip(n2449), .ck(clk), .q(
        \ANSWER/mem[8][5][13] ) );
  dp_1 \ANSWER/mem_reg[8][6][13]  ( .ip(n2448), .ck(clk), .q(
        \ANSWER/mem[8][6][13] ) );
  dp_1 \ANSWER/mem_reg[8][7][13]  ( .ip(n2447), .ck(clk), .q(
        \ANSWER/mem[8][7][13] ) );
  dp_1 \ANSWER/mem_reg[8][8][13]  ( .ip(n2446), .ck(clk), .q(
        \ANSWER/mem[8][8][13] ) );
  dp_1 \ANSWER/mem_reg[8][9][13]  ( .ip(n2445), .ck(clk), .q(
        \ANSWER/mem[8][9][13] ) );
  dp_1 \ANSWER/mem_reg[9][0][13]  ( .ip(n2444), .ck(clk), .q(
        \ANSWER/mem[9][0][13] ) );
  dp_1 \ANSWER/mem_reg[9][1][13]  ( .ip(n2443), .ck(clk), .q(
        \ANSWER/mem[9][1][13] ) );
  dp_1 \ANSWER/mem_reg[9][2][13]  ( .ip(n2442), .ck(clk), .q(
        \ANSWER/mem[9][2][13] ) );
  dp_1 \ANSWER/mem_reg[9][3][13]  ( .ip(n2441), .ck(clk), .q(
        \ANSWER/mem[9][3][13] ) );
  dp_1 \ANSWER/mem_reg[9][4][13]  ( .ip(n2440), .ck(clk), .q(
        \ANSWER/mem[9][4][13] ) );
  dp_1 \ANSWER/mem_reg[9][5][13]  ( .ip(n2439), .ck(clk), .q(
        \ANSWER/mem[9][5][13] ) );
  dp_1 \ANSWER/mem_reg[9][6][13]  ( .ip(n2438), .ck(clk), .q(
        \ANSWER/mem[9][6][13] ) );
  dp_1 \ANSWER/mem_reg[9][7][13]  ( .ip(n2437), .ck(clk), .q(
        \ANSWER/mem[9][7][13] ) );
  dp_1 \ANSWER/mem_reg[9][8][13]  ( .ip(n2436), .ck(clk), .q(
        \ANSWER/mem[9][8][13] ) );
  dp_1 \ANSWER/mem_reg[9][9][13]  ( .ip(n2435), .ck(clk), .q(
        \ANSWER/mem[9][9][13] ) );
  dp_1 \ANSWER/mem_reg[0][0][14]  ( .ip(n2434), .ck(clk), .q(
        \ANSWER/mem[0][0][14] ) );
  dp_1 \ANSWER/mem_reg[0][1][14]  ( .ip(n2433), .ck(clk), .q(
        \ANSWER/mem[0][1][14] ) );
  dp_1 \ANSWER/mem_reg[0][2][14]  ( .ip(n2432), .ck(clk), .q(
        \ANSWER/mem[0][2][14] ) );
  dp_1 \ANSWER/mem_reg[0][3][14]  ( .ip(n2431), .ck(clk), .q(
        \ANSWER/mem[0][3][14] ) );
  dp_1 \ANSWER/mem_reg[0][4][14]  ( .ip(n2430), .ck(clk), .q(
        \ANSWER/mem[0][4][14] ) );
  dp_1 \ANSWER/mem_reg[0][5][14]  ( .ip(n2429), .ck(clk), .q(
        \ANSWER/mem[0][5][14] ) );
  dp_1 \ANSWER/mem_reg[0][6][14]  ( .ip(n2428), .ck(clk), .q(
        \ANSWER/mem[0][6][14] ) );
  dp_1 \ANSWER/mem_reg[0][7][14]  ( .ip(n2427), .ck(clk), .q(
        \ANSWER/mem[0][7][14] ) );
  dp_1 \ANSWER/mem_reg[0][8][14]  ( .ip(n2426), .ck(clk), .q(
        \ANSWER/mem[0][8][14] ) );
  dp_1 \ANSWER/mem_reg[0][9][14]  ( .ip(n2425), .ck(clk), .q(
        \ANSWER/mem[0][9][14] ) );
  dp_1 \ANSWER/mem_reg[1][0][14]  ( .ip(n2424), .ck(clk), .q(
        \ANSWER/mem[1][0][14] ) );
  dp_1 \ANSWER/mem_reg[1][1][14]  ( .ip(n2423), .ck(clk), .q(
        \ANSWER/mem[1][1][14] ) );
  dp_1 \ANSWER/mem_reg[1][2][14]  ( .ip(n2422), .ck(clk), .q(
        \ANSWER/mem[1][2][14] ) );
  dp_1 \ANSWER/mem_reg[1][3][14]  ( .ip(n2421), .ck(clk), .q(
        \ANSWER/mem[1][3][14] ) );
  dp_1 \ANSWER/mem_reg[1][4][14]  ( .ip(n2420), .ck(clk), .q(
        \ANSWER/mem[1][4][14] ) );
  dp_1 \ANSWER/mem_reg[1][5][14]  ( .ip(n2419), .ck(clk), .q(
        \ANSWER/mem[1][5][14] ) );
  dp_1 \ANSWER/mem_reg[1][6][14]  ( .ip(n2418), .ck(clk), .q(
        \ANSWER/mem[1][6][14] ) );
  dp_1 \ANSWER/mem_reg[1][7][14]  ( .ip(n2417), .ck(clk), .q(
        \ANSWER/mem[1][7][14] ) );
  dp_1 \ANSWER/mem_reg[1][8][14]  ( .ip(n2416), .ck(clk), .q(
        \ANSWER/mem[1][8][14] ) );
  dp_1 \ANSWER/mem_reg[1][9][14]  ( .ip(n2415), .ck(clk), .q(
        \ANSWER/mem[1][9][14] ) );
  dp_1 \ANSWER/mem_reg[2][0][14]  ( .ip(n2414), .ck(clk), .q(
        \ANSWER/mem[2][0][14] ) );
  dp_1 \ANSWER/mem_reg[2][1][14]  ( .ip(n2413), .ck(clk), .q(
        \ANSWER/mem[2][1][14] ) );
  dp_1 \ANSWER/mem_reg[2][2][14]  ( .ip(n2412), .ck(clk), .q(
        \ANSWER/mem[2][2][14] ) );
  dp_1 \ANSWER/mem_reg[2][3][14]  ( .ip(n2411), .ck(clk), .q(
        \ANSWER/mem[2][3][14] ) );
  dp_1 \ANSWER/mem_reg[2][4][14]  ( .ip(n2410), .ck(clk), .q(
        \ANSWER/mem[2][4][14] ) );
  dp_1 \ANSWER/mem_reg[2][5][14]  ( .ip(n2409), .ck(clk), .q(
        \ANSWER/mem[2][5][14] ) );
  dp_1 \ANSWER/mem_reg[2][6][14]  ( .ip(n2408), .ck(clk), .q(
        \ANSWER/mem[2][6][14] ) );
  dp_1 \ANSWER/mem_reg[2][7][14]  ( .ip(n2407), .ck(clk), .q(
        \ANSWER/mem[2][7][14] ) );
  dp_1 \ANSWER/mem_reg[2][8][14]  ( .ip(n2406), .ck(clk), .q(
        \ANSWER/mem[2][8][14] ) );
  dp_1 \ANSWER/mem_reg[2][9][14]  ( .ip(n2405), .ck(clk), .q(
        \ANSWER/mem[2][9][14] ) );
  dp_1 \ANSWER/mem_reg[3][0][14]  ( .ip(n2404), .ck(clk), .q(
        \ANSWER/mem[3][0][14] ) );
  dp_1 \ANSWER/mem_reg[3][1][14]  ( .ip(n2403), .ck(clk), .q(
        \ANSWER/mem[3][1][14] ) );
  dp_1 \ANSWER/mem_reg[3][2][14]  ( .ip(n2402), .ck(clk), .q(
        \ANSWER/mem[3][2][14] ) );
  dp_1 \ANSWER/mem_reg[3][3][14]  ( .ip(n2401), .ck(clk), .q(
        \ANSWER/mem[3][3][14] ) );
  dp_1 \ANSWER/mem_reg[3][4][14]  ( .ip(n2400), .ck(clk), .q(
        \ANSWER/mem[3][4][14] ) );
  dp_1 \ANSWER/mem_reg[3][5][14]  ( .ip(n2399), .ck(clk), .q(
        \ANSWER/mem[3][5][14] ) );
  dp_1 \ANSWER/mem_reg[3][6][14]  ( .ip(n2398), .ck(clk), .q(
        \ANSWER/mem[3][6][14] ) );
  dp_1 \ANSWER/mem_reg[3][7][14]  ( .ip(n2397), .ck(clk), .q(
        \ANSWER/mem[3][7][14] ) );
  dp_1 \ANSWER/mem_reg[3][8][14]  ( .ip(n2396), .ck(clk), .q(
        \ANSWER/mem[3][8][14] ) );
  dp_1 \ANSWER/mem_reg[3][9][14]  ( .ip(n2395), .ck(clk), .q(
        \ANSWER/mem[3][9][14] ) );
  dp_1 \ANSWER/mem_reg[4][0][14]  ( .ip(n2394), .ck(clk), .q(
        \ANSWER/mem[4][0][14] ) );
  dp_1 \ANSWER/mem_reg[4][1][14]  ( .ip(n2393), .ck(clk), .q(
        \ANSWER/mem[4][1][14] ) );
  dp_1 \ANSWER/mem_reg[4][2][14]  ( .ip(n2392), .ck(clk), .q(
        \ANSWER/mem[4][2][14] ) );
  dp_1 \ANSWER/mem_reg[4][3][14]  ( .ip(n2391), .ck(clk), .q(
        \ANSWER/mem[4][3][14] ) );
  dp_1 \ANSWER/mem_reg[4][4][14]  ( .ip(n2390), .ck(clk), .q(
        \ANSWER/mem[4][4][14] ) );
  dp_1 \ANSWER/mem_reg[4][5][14]  ( .ip(n2389), .ck(clk), .q(
        \ANSWER/mem[4][5][14] ) );
  dp_1 \ANSWER/mem_reg[4][6][14]  ( .ip(n2388), .ck(clk), .q(
        \ANSWER/mem[4][6][14] ) );
  dp_1 \ANSWER/mem_reg[4][7][14]  ( .ip(n2387), .ck(clk), .q(
        \ANSWER/mem[4][7][14] ) );
  dp_1 \ANSWER/mem_reg[4][8][14]  ( .ip(n2386), .ck(clk), .q(
        \ANSWER/mem[4][8][14] ) );
  dp_1 \ANSWER/mem_reg[4][9][14]  ( .ip(n2385), .ck(clk), .q(
        \ANSWER/mem[4][9][14] ) );
  dp_1 \ANSWER/mem_reg[5][0][14]  ( .ip(n2384), .ck(clk), .q(
        \ANSWER/mem[5][0][14] ) );
  dp_1 \ANSWER/mem_reg[5][1][14]  ( .ip(n2383), .ck(clk), .q(
        \ANSWER/mem[5][1][14] ) );
  dp_1 \ANSWER/mem_reg[5][2][14]  ( .ip(n2382), .ck(clk), .q(
        \ANSWER/mem[5][2][14] ) );
  dp_1 \ANSWER/mem_reg[5][3][14]  ( .ip(n2381), .ck(clk), .q(
        \ANSWER/mem[5][3][14] ) );
  dp_1 \ANSWER/mem_reg[5][4][14]  ( .ip(n2380), .ck(clk), .q(
        \ANSWER/mem[5][4][14] ) );
  dp_1 \ANSWER/mem_reg[5][5][14]  ( .ip(n2379), .ck(clk), .q(
        \ANSWER/mem[5][5][14] ) );
  dp_1 \ANSWER/mem_reg[5][6][14]  ( .ip(n2378), .ck(clk), .q(
        \ANSWER/mem[5][6][14] ) );
  dp_1 \ANSWER/mem_reg[5][7][14]  ( .ip(n2377), .ck(clk), .q(
        \ANSWER/mem[5][7][14] ) );
  dp_1 \ANSWER/mem_reg[5][8][14]  ( .ip(n2376), .ck(clk), .q(
        \ANSWER/mem[5][8][14] ) );
  dp_1 \ANSWER/mem_reg[5][9][14]  ( .ip(n2375), .ck(clk), .q(
        \ANSWER/mem[5][9][14] ) );
  dp_1 \ANSWER/mem_reg[6][0][14]  ( .ip(n2374), .ck(clk), .q(
        \ANSWER/mem[6][0][14] ) );
  dp_1 \ANSWER/mem_reg[6][1][14]  ( .ip(n2373), .ck(clk), .q(
        \ANSWER/mem[6][1][14] ) );
  dp_1 \ANSWER/mem_reg[6][2][14]  ( .ip(n2372), .ck(clk), .q(
        \ANSWER/mem[6][2][14] ) );
  dp_1 \ANSWER/mem_reg[6][3][14]  ( .ip(n2371), .ck(clk), .q(
        \ANSWER/mem[6][3][14] ) );
  dp_1 \ANSWER/mem_reg[6][4][14]  ( .ip(n2370), .ck(clk), .q(
        \ANSWER/mem[6][4][14] ) );
  dp_1 \ANSWER/mem_reg[6][5][14]  ( .ip(n2369), .ck(clk), .q(
        \ANSWER/mem[6][5][14] ) );
  dp_1 \ANSWER/mem_reg[6][6][14]  ( .ip(n2368), .ck(clk), .q(
        \ANSWER/mem[6][6][14] ) );
  dp_1 \ANSWER/mem_reg[6][7][14]  ( .ip(n2367), .ck(clk), .q(
        \ANSWER/mem[6][7][14] ) );
  dp_1 \ANSWER/mem_reg[6][8][14]  ( .ip(n2366), .ck(clk), .q(
        \ANSWER/mem[6][8][14] ) );
  dp_1 \ANSWER/mem_reg[6][9][14]  ( .ip(n2365), .ck(clk), .q(
        \ANSWER/mem[6][9][14] ) );
  dp_1 \ANSWER/mem_reg[7][0][14]  ( .ip(n2364), .ck(clk), .q(
        \ANSWER/mem[7][0][14] ) );
  dp_1 \ANSWER/mem_reg[7][1][14]  ( .ip(n2363), .ck(clk), .q(
        \ANSWER/mem[7][1][14] ) );
  dp_1 \ANSWER/mem_reg[7][2][14]  ( .ip(n2362), .ck(clk), .q(
        \ANSWER/mem[7][2][14] ) );
  dp_1 \ANSWER/mem_reg[7][3][14]  ( .ip(n2361), .ck(clk), .q(
        \ANSWER/mem[7][3][14] ) );
  dp_1 \ANSWER/mem_reg[7][4][14]  ( .ip(n2360), .ck(clk), .q(
        \ANSWER/mem[7][4][14] ) );
  dp_1 \ANSWER/mem_reg[7][5][14]  ( .ip(n2359), .ck(clk), .q(
        \ANSWER/mem[7][5][14] ) );
  dp_1 \ANSWER/mem_reg[7][6][14]  ( .ip(n2358), .ck(clk), .q(
        \ANSWER/mem[7][6][14] ) );
  dp_1 \ANSWER/mem_reg[7][7][14]  ( .ip(n2357), .ck(clk), .q(
        \ANSWER/mem[7][7][14] ) );
  dp_1 \ANSWER/mem_reg[7][8][14]  ( .ip(n2356), .ck(clk), .q(
        \ANSWER/mem[7][8][14] ) );
  dp_1 \ANSWER/mem_reg[7][9][14]  ( .ip(n2355), .ck(clk), .q(
        \ANSWER/mem[7][9][14] ) );
  dp_1 \ANSWER/mem_reg[8][0][14]  ( .ip(n2354), .ck(clk), .q(
        \ANSWER/mem[8][0][14] ) );
  dp_1 \ANSWER/mem_reg[8][1][14]  ( .ip(n2353), .ck(clk), .q(
        \ANSWER/mem[8][1][14] ) );
  dp_1 \ANSWER/mem_reg[8][2][14]  ( .ip(n2352), .ck(clk), .q(
        \ANSWER/mem[8][2][14] ) );
  dp_1 \ANSWER/mem_reg[8][3][14]  ( .ip(n2351), .ck(clk), .q(
        \ANSWER/mem[8][3][14] ) );
  dp_1 \ANSWER/mem_reg[8][4][14]  ( .ip(n2350), .ck(clk), .q(
        \ANSWER/mem[8][4][14] ) );
  dp_1 \ANSWER/mem_reg[8][5][14]  ( .ip(n2349), .ck(clk), .q(
        \ANSWER/mem[8][5][14] ) );
  dp_1 \ANSWER/mem_reg[8][6][14]  ( .ip(n2348), .ck(clk), .q(
        \ANSWER/mem[8][6][14] ) );
  dp_1 \ANSWER/mem_reg[8][7][14]  ( .ip(n2347), .ck(clk), .q(
        \ANSWER/mem[8][7][14] ) );
  dp_1 \ANSWER/mem_reg[8][8][14]  ( .ip(n2346), .ck(clk), .q(
        \ANSWER/mem[8][8][14] ) );
  dp_1 \ANSWER/mem_reg[8][9][14]  ( .ip(n2345), .ck(clk), .q(
        \ANSWER/mem[8][9][14] ) );
  dp_1 \ANSWER/mem_reg[9][0][14]  ( .ip(n2344), .ck(clk), .q(
        \ANSWER/mem[9][0][14] ) );
  dp_1 \ANSWER/mem_reg[9][1][14]  ( .ip(n2343), .ck(clk), .q(
        \ANSWER/mem[9][1][14] ) );
  dp_1 \ANSWER/mem_reg[9][2][14]  ( .ip(n2342), .ck(clk), .q(
        \ANSWER/mem[9][2][14] ) );
  dp_1 \ANSWER/mem_reg[9][3][14]  ( .ip(n2341), .ck(clk), .q(
        \ANSWER/mem[9][3][14] ) );
  dp_1 \ANSWER/mem_reg[9][4][14]  ( .ip(n2340), .ck(clk), .q(
        \ANSWER/mem[9][4][14] ) );
  dp_1 \ANSWER/mem_reg[9][5][14]  ( .ip(n2339), .ck(clk), .q(
        \ANSWER/mem[9][5][14] ) );
  dp_1 \ANSWER/mem_reg[9][6][14]  ( .ip(n2338), .ck(clk), .q(
        \ANSWER/mem[9][6][14] ) );
  dp_1 \ANSWER/mem_reg[9][7][14]  ( .ip(n2337), .ck(clk), .q(
        \ANSWER/mem[9][7][14] ) );
  dp_1 \ANSWER/mem_reg[9][8][14]  ( .ip(n2336), .ck(clk), .q(
        \ANSWER/mem[9][8][14] ) );
  dp_1 \ANSWER/mem_reg[9][9][14]  ( .ip(n2335), .ck(clk), .q(
        \ANSWER/mem[9][9][14] ) );
  dp_1 \ANSWER/mem_reg[0][0][15]  ( .ip(n2334), .ck(clk), .q(
        \ANSWER/mem[0][0][15] ) );
  dp_1 \ANSWER/mem_reg[0][1][15]  ( .ip(n2333), .ck(clk), .q(
        \ANSWER/mem[0][1][15] ) );
  dp_1 \ANSWER/mem_reg[0][2][15]  ( .ip(n2332), .ck(clk), .q(
        \ANSWER/mem[0][2][15] ) );
  dp_1 \ANSWER/mem_reg[0][3][15]  ( .ip(n2331), .ck(clk), .q(
        \ANSWER/mem[0][3][15] ) );
  dp_1 \ANSWER/mem_reg[0][4][15]  ( .ip(n2330), .ck(clk), .q(
        \ANSWER/mem[0][4][15] ) );
  dp_1 \ANSWER/mem_reg[0][5][15]  ( .ip(n2329), .ck(clk), .q(
        \ANSWER/mem[0][5][15] ) );
  dp_1 \ANSWER/mem_reg[0][6][15]  ( .ip(n2328), .ck(clk), .q(
        \ANSWER/mem[0][6][15] ) );
  dp_1 \ANSWER/mem_reg[0][7][15]  ( .ip(n2327), .ck(clk), .q(
        \ANSWER/mem[0][7][15] ) );
  dp_1 \ANSWER/mem_reg[0][8][15]  ( .ip(n2326), .ck(clk), .q(
        \ANSWER/mem[0][8][15] ) );
  dp_1 \ANSWER/mem_reg[0][9][15]  ( .ip(n2325), .ck(clk), .q(
        \ANSWER/mem[0][9][15] ) );
  dp_1 \ANSWER/mem_reg[1][0][15]  ( .ip(n2324), .ck(clk), .q(
        \ANSWER/mem[1][0][15] ) );
  dp_1 \ANSWER/mem_reg[1][1][15]  ( .ip(n2323), .ck(clk), .q(
        \ANSWER/mem[1][1][15] ) );
  dp_1 \ANSWER/mem_reg[1][2][15]  ( .ip(n2322), .ck(clk), .q(
        \ANSWER/mem[1][2][15] ) );
  dp_1 \ANSWER/mem_reg[1][3][15]  ( .ip(n2321), .ck(clk), .q(
        \ANSWER/mem[1][3][15] ) );
  dp_1 \ANSWER/mem_reg[1][4][15]  ( .ip(n2320), .ck(clk), .q(
        \ANSWER/mem[1][4][15] ) );
  dp_1 \ANSWER/mem_reg[1][5][15]  ( .ip(n2319), .ck(clk), .q(
        \ANSWER/mem[1][5][15] ) );
  dp_1 \ANSWER/mem_reg[1][6][15]  ( .ip(n2318), .ck(clk), .q(
        \ANSWER/mem[1][6][15] ) );
  dp_1 \ANSWER/mem_reg[1][7][15]  ( .ip(n2317), .ck(clk), .q(
        \ANSWER/mem[1][7][15] ) );
  dp_1 \ANSWER/mem_reg[1][8][15]  ( .ip(n2316), .ck(clk), .q(
        \ANSWER/mem[1][8][15] ) );
  dp_1 \ANSWER/mem_reg[1][9][15]  ( .ip(n2315), .ck(clk), .q(
        \ANSWER/mem[1][9][15] ) );
  dp_1 \ANSWER/mem_reg[2][0][15]  ( .ip(n2314), .ck(clk), .q(
        \ANSWER/mem[2][0][15] ) );
  dp_1 \ANSWER/mem_reg[2][1][15]  ( .ip(n2313), .ck(clk), .q(
        \ANSWER/mem[2][1][15] ) );
  dp_1 \ANSWER/mem_reg[2][2][15]  ( .ip(n2312), .ck(clk), .q(
        \ANSWER/mem[2][2][15] ) );
  dp_1 \ANSWER/mem_reg[2][3][15]  ( .ip(n2311), .ck(clk), .q(
        \ANSWER/mem[2][3][15] ) );
  dp_1 \ANSWER/mem_reg[2][4][15]  ( .ip(n2310), .ck(clk), .q(
        \ANSWER/mem[2][4][15] ) );
  dp_1 \ANSWER/mem_reg[2][5][15]  ( .ip(n2309), .ck(clk), .q(
        \ANSWER/mem[2][5][15] ) );
  dp_1 \ANSWER/mem_reg[2][6][15]  ( .ip(n2308), .ck(clk), .q(
        \ANSWER/mem[2][6][15] ) );
  dp_1 \ANSWER/mem_reg[2][7][15]  ( .ip(n2307), .ck(clk), .q(
        \ANSWER/mem[2][7][15] ) );
  dp_1 \ANSWER/mem_reg[2][8][15]  ( .ip(n2306), .ck(clk), .q(
        \ANSWER/mem[2][8][15] ) );
  dp_1 \ANSWER/mem_reg[2][9][15]  ( .ip(n2305), .ck(clk), .q(
        \ANSWER/mem[2][9][15] ) );
  dp_1 \ANSWER/mem_reg[3][0][15]  ( .ip(n2304), .ck(clk), .q(
        \ANSWER/mem[3][0][15] ) );
  dp_1 \ANSWER/mem_reg[3][1][15]  ( .ip(n2303), .ck(clk), .q(
        \ANSWER/mem[3][1][15] ) );
  dp_1 \ANSWER/mem_reg[3][2][15]  ( .ip(n2302), .ck(clk), .q(
        \ANSWER/mem[3][2][15] ) );
  dp_1 \ANSWER/mem_reg[3][3][15]  ( .ip(n2301), .ck(clk), .q(
        \ANSWER/mem[3][3][15] ) );
  dp_1 \ANSWER/mem_reg[3][4][15]  ( .ip(n2300), .ck(clk), .q(
        \ANSWER/mem[3][4][15] ) );
  dp_1 \ANSWER/mem_reg[3][5][15]  ( .ip(n2299), .ck(clk), .q(
        \ANSWER/mem[3][5][15] ) );
  dp_1 \ANSWER/mem_reg[3][6][15]  ( .ip(n2298), .ck(clk), .q(
        \ANSWER/mem[3][6][15] ) );
  dp_1 \ANSWER/mem_reg[3][7][15]  ( .ip(n2297), .ck(clk), .q(
        \ANSWER/mem[3][7][15] ) );
  dp_1 \ANSWER/mem_reg[3][8][15]  ( .ip(n2296), .ck(clk), .q(
        \ANSWER/mem[3][8][15] ) );
  dp_1 \ANSWER/mem_reg[3][9][15]  ( .ip(n2295), .ck(clk), .q(
        \ANSWER/mem[3][9][15] ) );
  dp_1 \ANSWER/mem_reg[4][0][15]  ( .ip(n2294), .ck(clk), .q(
        \ANSWER/mem[4][0][15] ) );
  dp_1 \ANSWER/mem_reg[4][1][15]  ( .ip(n2293), .ck(clk), .q(
        \ANSWER/mem[4][1][15] ) );
  dp_1 \ANSWER/mem_reg[4][2][15]  ( .ip(n2292), .ck(clk), .q(
        \ANSWER/mem[4][2][15] ) );
  dp_1 \ANSWER/mem_reg[4][3][15]  ( .ip(n2291), .ck(clk), .q(
        \ANSWER/mem[4][3][15] ) );
  dp_1 \ANSWER/mem_reg[4][4][15]  ( .ip(n2290), .ck(clk), .q(
        \ANSWER/mem[4][4][15] ) );
  dp_1 \ANSWER/mem_reg[4][5][15]  ( .ip(n2289), .ck(clk), .q(
        \ANSWER/mem[4][5][15] ) );
  dp_1 \ANSWER/mem_reg[4][6][15]  ( .ip(n2288), .ck(clk), .q(
        \ANSWER/mem[4][6][15] ) );
  dp_1 \ANSWER/mem_reg[4][7][15]  ( .ip(n2287), .ck(clk), .q(
        \ANSWER/mem[4][7][15] ) );
  dp_1 \ANSWER/mem_reg[4][8][15]  ( .ip(n2286), .ck(clk), .q(
        \ANSWER/mem[4][8][15] ) );
  dp_1 \ANSWER/mem_reg[4][9][15]  ( .ip(n2285), .ck(clk), .q(
        \ANSWER/mem[4][9][15] ) );
  dp_1 \ANSWER/mem_reg[5][0][15]  ( .ip(n2284), .ck(clk), .q(
        \ANSWER/mem[5][0][15] ) );
  dp_1 \ANSWER/mem_reg[5][1][15]  ( .ip(n2283), .ck(clk), .q(
        \ANSWER/mem[5][1][15] ) );
  dp_1 \ANSWER/mem_reg[5][2][15]  ( .ip(n2282), .ck(clk), .q(
        \ANSWER/mem[5][2][15] ) );
  dp_1 \ANSWER/mem_reg[5][3][15]  ( .ip(n2281), .ck(clk), .q(
        \ANSWER/mem[5][3][15] ) );
  dp_1 \ANSWER/mem_reg[5][4][15]  ( .ip(n2280), .ck(clk), .q(
        \ANSWER/mem[5][4][15] ) );
  dp_1 \ANSWER/mem_reg[5][5][15]  ( .ip(n2279), .ck(clk), .q(
        \ANSWER/mem[5][5][15] ) );
  dp_1 \ANSWER/mem_reg[5][6][15]  ( .ip(n2278), .ck(clk), .q(
        \ANSWER/mem[5][6][15] ) );
  dp_1 \ANSWER/mem_reg[5][7][15]  ( .ip(n2277), .ck(clk), .q(
        \ANSWER/mem[5][7][15] ) );
  dp_1 \ANSWER/mem_reg[5][8][15]  ( .ip(n2276), .ck(clk), .q(
        \ANSWER/mem[5][8][15] ) );
  dp_1 \ANSWER/mem_reg[5][9][15]  ( .ip(n2275), .ck(clk), .q(
        \ANSWER/mem[5][9][15] ) );
  dp_1 \ANSWER/mem_reg[6][0][15]  ( .ip(n2274), .ck(clk), .q(
        \ANSWER/mem[6][0][15] ) );
  dp_1 \ANSWER/mem_reg[6][1][15]  ( .ip(n2273), .ck(clk), .q(
        \ANSWER/mem[6][1][15] ) );
  dp_1 \ANSWER/mem_reg[6][2][15]  ( .ip(n2272), .ck(clk), .q(
        \ANSWER/mem[6][2][15] ) );
  dp_1 \ANSWER/mem_reg[6][3][15]  ( .ip(n2271), .ck(clk), .q(
        \ANSWER/mem[6][3][15] ) );
  dp_1 \ANSWER/mem_reg[6][4][15]  ( .ip(n2270), .ck(clk), .q(
        \ANSWER/mem[6][4][15] ) );
  dp_1 \ANSWER/mem_reg[6][5][15]  ( .ip(n2269), .ck(clk), .q(
        \ANSWER/mem[6][5][15] ) );
  dp_1 \ANSWER/mem_reg[6][6][15]  ( .ip(n2268), .ck(clk), .q(
        \ANSWER/mem[6][6][15] ) );
  dp_1 \ANSWER/mem_reg[6][7][15]  ( .ip(n2267), .ck(clk), .q(
        \ANSWER/mem[6][7][15] ) );
  dp_1 \ANSWER/mem_reg[6][8][15]  ( .ip(n2266), .ck(clk), .q(
        \ANSWER/mem[6][8][15] ) );
  dp_1 \ANSWER/mem_reg[6][9][15]  ( .ip(n2265), .ck(clk), .q(
        \ANSWER/mem[6][9][15] ) );
  dp_1 \ANSWER/mem_reg[7][0][15]  ( .ip(n2264), .ck(clk), .q(
        \ANSWER/mem[7][0][15] ) );
  dp_1 \ANSWER/mem_reg[7][1][15]  ( .ip(n2263), .ck(clk), .q(
        \ANSWER/mem[7][1][15] ) );
  dp_1 \ANSWER/mem_reg[7][2][15]  ( .ip(n2262), .ck(clk), .q(
        \ANSWER/mem[7][2][15] ) );
  dp_1 \ANSWER/mem_reg[7][3][15]  ( .ip(n2261), .ck(clk), .q(
        \ANSWER/mem[7][3][15] ) );
  dp_1 \ANSWER/mem_reg[7][4][15]  ( .ip(n2260), .ck(clk), .q(
        \ANSWER/mem[7][4][15] ) );
  dp_1 \ANSWER/mem_reg[7][5][15]  ( .ip(n2259), .ck(clk), .q(
        \ANSWER/mem[7][5][15] ) );
  dp_1 \ANSWER/mem_reg[7][6][15]  ( .ip(n2258), .ck(clk), .q(
        \ANSWER/mem[7][6][15] ) );
  dp_1 \ANSWER/mem_reg[7][7][15]  ( .ip(n2257), .ck(clk), .q(
        \ANSWER/mem[7][7][15] ) );
  dp_1 \ANSWER/mem_reg[7][8][15]  ( .ip(n2256), .ck(clk), .q(
        \ANSWER/mem[7][8][15] ) );
  dp_1 \ANSWER/mem_reg[7][9][15]  ( .ip(n2255), .ck(clk), .q(
        \ANSWER/mem[7][9][15] ) );
  dp_1 \ANSWER/mem_reg[8][0][15]  ( .ip(n2254), .ck(clk), .q(
        \ANSWER/mem[8][0][15] ) );
  dp_1 \ANSWER/mem_reg[8][1][15]  ( .ip(n2253), .ck(clk), .q(
        \ANSWER/mem[8][1][15] ) );
  dp_1 \ANSWER/mem_reg[8][2][15]  ( .ip(n2252), .ck(clk), .q(
        \ANSWER/mem[8][2][15] ) );
  dp_1 \ANSWER/mem_reg[8][3][15]  ( .ip(n2251), .ck(clk), .q(
        \ANSWER/mem[8][3][15] ) );
  dp_1 \ANSWER/mem_reg[8][4][15]  ( .ip(n2250), .ck(clk), .q(
        \ANSWER/mem[8][4][15] ) );
  dp_1 \ANSWER/mem_reg[8][5][15]  ( .ip(n2249), .ck(clk), .q(
        \ANSWER/mem[8][5][15] ) );
  dp_1 \ANSWER/mem_reg[8][6][15]  ( .ip(n2248), .ck(clk), .q(
        \ANSWER/mem[8][6][15] ) );
  dp_1 \ANSWER/mem_reg[8][7][15]  ( .ip(n2247), .ck(clk), .q(
        \ANSWER/mem[8][7][15] ) );
  dp_1 \ANSWER/mem_reg[8][8][15]  ( .ip(n2246), .ck(clk), .q(
        \ANSWER/mem[8][8][15] ) );
  dp_1 \ANSWER/mem_reg[8][9][15]  ( .ip(n2245), .ck(clk), .q(
        \ANSWER/mem[8][9][15] ) );
  dp_1 \ANSWER/mem_reg[9][0][15]  ( .ip(n2244), .ck(clk), .q(
        \ANSWER/mem[9][0][15] ) );
  dp_1 \ANSWER/mem_reg[9][1][15]  ( .ip(n2243), .ck(clk), .q(
        \ANSWER/mem[9][1][15] ) );
  dp_1 \ANSWER/mem_reg[9][2][15]  ( .ip(n2242), .ck(clk), .q(
        \ANSWER/mem[9][2][15] ) );
  dp_1 \ANSWER/mem_reg[9][3][15]  ( .ip(n2241), .ck(clk), .q(
        \ANSWER/mem[9][3][15] ) );
  dp_1 \ANSWER/mem_reg[9][4][15]  ( .ip(n2240), .ck(clk), .q(
        \ANSWER/mem[9][4][15] ) );
  dp_1 \ANSWER/mem_reg[9][5][15]  ( .ip(n2239), .ck(clk), .q(
        \ANSWER/mem[9][5][15] ) );
  dp_1 \ANSWER/mem_reg[9][6][15]  ( .ip(n2238), .ck(clk), .q(
        \ANSWER/mem[9][6][15] ) );
  dp_1 \ANSWER/mem_reg[9][7][15]  ( .ip(n2237), .ck(clk), .q(
        \ANSWER/mem[9][7][15] ) );
  dp_1 \ANSWER/mem_reg[9][8][15]  ( .ip(n2236), .ck(clk), .q(
        \ANSWER/mem[9][8][15] ) );
  dp_1 \ANSWER/mem_reg[9][9][15]  ( .ip(n2235), .ck(clk), .q(
        \ANSWER/mem[9][9][15] ) );
  dp_1 \SIGMOID/lut_out_reg[0]  ( .ip(n3842), .ck(clk), .q(\SIGMOID/N64 ) );
  dp_1 \ANSWER/mem_reg[0][0][0]  ( .ip(n3834), .ck(clk), .q(
        \ANSWER/mem[0][0][0] ) );
  dp_1 \ANSWER/mem_reg[0][1][0]  ( .ip(n3833), .ck(clk), .q(
        \ANSWER/mem[0][1][0] ) );
  dp_1 \ANSWER/mem_reg[0][2][0]  ( .ip(n3832), .ck(clk), .q(
        \ANSWER/mem[0][2][0] ) );
  dp_1 \ANSWER/mem_reg[0][3][0]  ( .ip(n3831), .ck(clk), .q(
        \ANSWER/mem[0][3][0] ) );
  dp_1 \ANSWER/mem_reg[0][4][0]  ( .ip(n3830), .ck(clk), .q(
        \ANSWER/mem[0][4][0] ) );
  dp_1 \ANSWER/mem_reg[0][5][0]  ( .ip(n3829), .ck(clk), .q(
        \ANSWER/mem[0][5][0] ) );
  dp_1 \ANSWER/mem_reg[0][6][0]  ( .ip(n3828), .ck(clk), .q(
        \ANSWER/mem[0][6][0] ) );
  dp_1 \ANSWER/mem_reg[0][7][0]  ( .ip(n3827), .ck(clk), .q(
        \ANSWER/mem[0][7][0] ) );
  dp_1 \ANSWER/mem_reg[0][8][0]  ( .ip(n3826), .ck(clk), .q(
        \ANSWER/mem[0][8][0] ) );
  dp_1 \ANSWER/mem_reg[0][9][0]  ( .ip(n3825), .ck(clk), .q(
        \ANSWER/mem[0][9][0] ) );
  dp_1 \ANSWER/mem_reg[1][0][0]  ( .ip(n3824), .ck(clk), .q(
        \ANSWER/mem[1][0][0] ) );
  dp_1 \ANSWER/mem_reg[1][1][0]  ( .ip(n3823), .ck(clk), .q(
        \ANSWER/mem[1][1][0] ) );
  dp_1 \ANSWER/mem_reg[1][2][0]  ( .ip(n3822), .ck(clk), .q(
        \ANSWER/mem[1][2][0] ) );
  dp_1 \ANSWER/mem_reg[1][3][0]  ( .ip(n3821), .ck(clk), .q(
        \ANSWER/mem[1][3][0] ) );
  dp_1 \ANSWER/mem_reg[1][4][0]  ( .ip(n3820), .ck(clk), .q(
        \ANSWER/mem[1][4][0] ) );
  dp_1 \ANSWER/mem_reg[1][5][0]  ( .ip(n3819), .ck(clk), .q(
        \ANSWER/mem[1][5][0] ) );
  dp_1 \ANSWER/mem_reg[1][6][0]  ( .ip(n3818), .ck(clk), .q(
        \ANSWER/mem[1][6][0] ) );
  dp_1 \ANSWER/mem_reg[1][7][0]  ( .ip(n3817), .ck(clk), .q(
        \ANSWER/mem[1][7][0] ) );
  dp_1 \ANSWER/mem_reg[1][8][0]  ( .ip(n3816), .ck(clk), .q(
        \ANSWER/mem[1][8][0] ) );
  dp_1 \ANSWER/mem_reg[1][9][0]  ( .ip(n3815), .ck(clk), .q(
        \ANSWER/mem[1][9][0] ) );
  dp_1 \ANSWER/mem_reg[2][0][0]  ( .ip(n3814), .ck(clk), .q(
        \ANSWER/mem[2][0][0] ) );
  dp_1 \ANSWER/mem_reg[2][1][0]  ( .ip(n3813), .ck(clk), .q(
        \ANSWER/mem[2][1][0] ) );
  dp_1 \ANSWER/mem_reg[2][2][0]  ( .ip(n3812), .ck(clk), .q(
        \ANSWER/mem[2][2][0] ) );
  dp_1 \ANSWER/mem_reg[2][3][0]  ( .ip(n3811), .ck(clk), .q(
        \ANSWER/mem[2][3][0] ) );
  dp_1 \ANSWER/mem_reg[2][4][0]  ( .ip(n3810), .ck(clk), .q(
        \ANSWER/mem[2][4][0] ) );
  dp_1 \ANSWER/mem_reg[2][5][0]  ( .ip(n3809), .ck(clk), .q(
        \ANSWER/mem[2][5][0] ) );
  dp_1 \ANSWER/mem_reg[2][6][0]  ( .ip(n3808), .ck(clk), .q(
        \ANSWER/mem[2][6][0] ) );
  dp_1 \ANSWER/mem_reg[2][7][0]  ( .ip(n3807), .ck(clk), .q(
        \ANSWER/mem[2][7][0] ) );
  dp_1 \ANSWER/mem_reg[2][8][0]  ( .ip(n3806), .ck(clk), .q(
        \ANSWER/mem[2][8][0] ) );
  dp_1 \ANSWER/mem_reg[2][9][0]  ( .ip(n3805), .ck(clk), .q(
        \ANSWER/mem[2][9][0] ) );
  dp_1 \ANSWER/mem_reg[3][0][0]  ( .ip(n3804), .ck(clk), .q(
        \ANSWER/mem[3][0][0] ) );
  dp_1 \ANSWER/mem_reg[3][1][0]  ( .ip(n3803), .ck(clk), .q(
        \ANSWER/mem[3][1][0] ) );
  dp_1 \ANSWER/mem_reg[3][2][0]  ( .ip(n3802), .ck(clk), .q(
        \ANSWER/mem[3][2][0] ) );
  dp_1 \ANSWER/mem_reg[3][3][0]  ( .ip(n3801), .ck(clk), .q(
        \ANSWER/mem[3][3][0] ) );
  dp_1 \ANSWER/mem_reg[3][4][0]  ( .ip(n3800), .ck(clk), .q(
        \ANSWER/mem[3][4][0] ) );
  dp_1 \ANSWER/mem_reg[3][5][0]  ( .ip(n3799), .ck(clk), .q(
        \ANSWER/mem[3][5][0] ) );
  dp_1 \ANSWER/mem_reg[3][6][0]  ( .ip(n3798), .ck(clk), .q(
        \ANSWER/mem[3][6][0] ) );
  dp_1 \ANSWER/mem_reg[3][7][0]  ( .ip(n3797), .ck(clk), .q(
        \ANSWER/mem[3][7][0] ) );
  dp_1 \ANSWER/mem_reg[3][8][0]  ( .ip(n3796), .ck(clk), .q(
        \ANSWER/mem[3][8][0] ) );
  dp_1 \ANSWER/mem_reg[3][9][0]  ( .ip(n3795), .ck(clk), .q(
        \ANSWER/mem[3][9][0] ) );
  dp_1 \ANSWER/mem_reg[4][0][0]  ( .ip(n3794), .ck(clk), .q(
        \ANSWER/mem[4][0][0] ) );
  dp_1 \ANSWER/mem_reg[4][1][0]  ( .ip(n3793), .ck(clk), .q(
        \ANSWER/mem[4][1][0] ) );
  dp_1 \ANSWER/mem_reg[4][2][0]  ( .ip(n3792), .ck(clk), .q(
        \ANSWER/mem[4][2][0] ) );
  dp_1 \ANSWER/mem_reg[4][3][0]  ( .ip(n3791), .ck(clk), .q(
        \ANSWER/mem[4][3][0] ) );
  dp_1 \ANSWER/mem_reg[4][4][0]  ( .ip(n3790), .ck(clk), .q(
        \ANSWER/mem[4][4][0] ) );
  dp_1 \ANSWER/mem_reg[4][5][0]  ( .ip(n3789), .ck(clk), .q(
        \ANSWER/mem[4][5][0] ) );
  dp_1 \ANSWER/mem_reg[4][6][0]  ( .ip(n3788), .ck(clk), .q(
        \ANSWER/mem[4][6][0] ) );
  dp_1 \ANSWER/mem_reg[4][7][0]  ( .ip(n3787), .ck(clk), .q(
        \ANSWER/mem[4][7][0] ) );
  dp_1 \ANSWER/mem_reg[4][8][0]  ( .ip(n3786), .ck(clk), .q(
        \ANSWER/mem[4][8][0] ) );
  dp_1 \ANSWER/mem_reg[4][9][0]  ( .ip(n3785), .ck(clk), .q(
        \ANSWER/mem[4][9][0] ) );
  dp_1 \ANSWER/mem_reg[5][0][0]  ( .ip(n3784), .ck(clk), .q(
        \ANSWER/mem[5][0][0] ) );
  dp_1 \ANSWER/mem_reg[5][1][0]  ( .ip(n3783), .ck(clk), .q(
        \ANSWER/mem[5][1][0] ) );
  dp_1 \ANSWER/mem_reg[5][2][0]  ( .ip(n3782), .ck(clk), .q(
        \ANSWER/mem[5][2][0] ) );
  dp_1 \ANSWER/mem_reg[5][3][0]  ( .ip(n3781), .ck(clk), .q(
        \ANSWER/mem[5][3][0] ) );
  dp_1 \ANSWER/mem_reg[5][4][0]  ( .ip(n3780), .ck(clk), .q(
        \ANSWER/mem[5][4][0] ) );
  dp_1 \ANSWER/mem_reg[5][5][0]  ( .ip(n3779), .ck(clk), .q(
        \ANSWER/mem[5][5][0] ) );
  dp_1 \ANSWER/mem_reg[5][6][0]  ( .ip(n3778), .ck(clk), .q(
        \ANSWER/mem[5][6][0] ) );
  dp_1 \ANSWER/mem_reg[5][7][0]  ( .ip(n3777), .ck(clk), .q(
        \ANSWER/mem[5][7][0] ) );
  dp_1 \ANSWER/mem_reg[5][8][0]  ( .ip(n3776), .ck(clk), .q(
        \ANSWER/mem[5][8][0] ) );
  dp_1 \ANSWER/mem_reg[5][9][0]  ( .ip(n3775), .ck(clk), .q(
        \ANSWER/mem[5][9][0] ) );
  dp_1 \ANSWER/mem_reg[6][0][0]  ( .ip(n3774), .ck(clk), .q(
        \ANSWER/mem[6][0][0] ) );
  dp_1 \ANSWER/mem_reg[6][1][0]  ( .ip(n3773), .ck(clk), .q(
        \ANSWER/mem[6][1][0] ) );
  dp_1 \ANSWER/mem_reg[6][2][0]  ( .ip(n3772), .ck(clk), .q(
        \ANSWER/mem[6][2][0] ) );
  dp_1 \ANSWER/mem_reg[6][3][0]  ( .ip(n3771), .ck(clk), .q(
        \ANSWER/mem[6][3][0] ) );
  dp_1 \ANSWER/mem_reg[6][4][0]  ( .ip(n3770), .ck(clk), .q(
        \ANSWER/mem[6][4][0] ) );
  dp_1 \ANSWER/mem_reg[6][5][0]  ( .ip(n3769), .ck(clk), .q(
        \ANSWER/mem[6][5][0] ) );
  dp_1 \ANSWER/mem_reg[6][6][0]  ( .ip(n3768), .ck(clk), .q(
        \ANSWER/mem[6][6][0] ) );
  dp_1 \ANSWER/mem_reg[6][7][0]  ( .ip(n3767), .ck(clk), .q(
        \ANSWER/mem[6][7][0] ) );
  dp_1 \ANSWER/mem_reg[6][8][0]  ( .ip(n3766), .ck(clk), .q(
        \ANSWER/mem[6][8][0] ) );
  dp_1 \ANSWER/mem_reg[6][9][0]  ( .ip(n3765), .ck(clk), .q(
        \ANSWER/mem[6][9][0] ) );
  dp_1 \ANSWER/mem_reg[7][0][0]  ( .ip(n3764), .ck(clk), .q(
        \ANSWER/mem[7][0][0] ) );
  dp_1 \ANSWER/mem_reg[7][1][0]  ( .ip(n3763), .ck(clk), .q(
        \ANSWER/mem[7][1][0] ) );
  dp_1 \ANSWER/mem_reg[7][2][0]  ( .ip(n3762), .ck(clk), .q(
        \ANSWER/mem[7][2][0] ) );
  dp_1 \ANSWER/mem_reg[7][3][0]  ( .ip(n3761), .ck(clk), .q(
        \ANSWER/mem[7][3][0] ) );
  dp_1 \ANSWER/mem_reg[7][4][0]  ( .ip(n3760), .ck(clk), .q(
        \ANSWER/mem[7][4][0] ) );
  dp_1 \ANSWER/mem_reg[7][5][0]  ( .ip(n3759), .ck(clk), .q(
        \ANSWER/mem[7][5][0] ) );
  dp_1 \ANSWER/mem_reg[7][6][0]  ( .ip(n3758), .ck(clk), .q(
        \ANSWER/mem[7][6][0] ) );
  dp_1 \ANSWER/mem_reg[7][7][0]  ( .ip(n3757), .ck(clk), .q(
        \ANSWER/mem[7][7][0] ) );
  dp_1 \ANSWER/mem_reg[7][8][0]  ( .ip(n3756), .ck(clk), .q(
        \ANSWER/mem[7][8][0] ) );
  dp_1 \ANSWER/mem_reg[7][9][0]  ( .ip(n3755), .ck(clk), .q(
        \ANSWER/mem[7][9][0] ) );
  dp_1 \ANSWER/mem_reg[8][0][0]  ( .ip(n3754), .ck(clk), .q(
        \ANSWER/mem[8][0][0] ) );
  dp_1 \ANSWER/mem_reg[8][1][0]  ( .ip(n3753), .ck(clk), .q(
        \ANSWER/mem[8][1][0] ) );
  dp_1 \ANSWER/mem_reg[8][2][0]  ( .ip(n3752), .ck(clk), .q(
        \ANSWER/mem[8][2][0] ) );
  dp_1 \ANSWER/mem_reg[8][3][0]  ( .ip(n3751), .ck(clk), .q(
        \ANSWER/mem[8][3][0] ) );
  dp_1 \ANSWER/mem_reg[8][4][0]  ( .ip(n3750), .ck(clk), .q(
        \ANSWER/mem[8][4][0] ) );
  dp_1 \ANSWER/mem_reg[8][5][0]  ( .ip(n3749), .ck(clk), .q(
        \ANSWER/mem[8][5][0] ) );
  dp_1 \ANSWER/mem_reg[8][6][0]  ( .ip(n3748), .ck(clk), .q(
        \ANSWER/mem[8][6][0] ) );
  dp_1 \ANSWER/mem_reg[8][7][0]  ( .ip(n3747), .ck(clk), .q(
        \ANSWER/mem[8][7][0] ) );
  dp_1 \ANSWER/mem_reg[8][8][0]  ( .ip(n3746), .ck(clk), .q(
        \ANSWER/mem[8][8][0] ) );
  dp_1 \ANSWER/mem_reg[8][9][0]  ( .ip(n3745), .ck(clk), .q(
        \ANSWER/mem[8][9][0] ) );
  dp_1 \ANSWER/mem_reg[9][0][0]  ( .ip(n3744), .ck(clk), .q(
        \ANSWER/mem[9][0][0] ) );
  dp_1 \ANSWER/mem_reg[9][1][0]  ( .ip(n3743), .ck(clk), .q(
        \ANSWER/mem[9][1][0] ) );
  dp_1 \ANSWER/mem_reg[9][2][0]  ( .ip(n3742), .ck(clk), .q(
        \ANSWER/mem[9][2][0] ) );
  dp_1 \ANSWER/mem_reg[9][3][0]  ( .ip(n3741), .ck(clk), .q(
        \ANSWER/mem[9][3][0] ) );
  dp_1 \ANSWER/mem_reg[9][4][0]  ( .ip(n3740), .ck(clk), .q(
        \ANSWER/mem[9][4][0] ) );
  dp_1 \ANSWER/mem_reg[9][5][0]  ( .ip(n3739), .ck(clk), .q(
        \ANSWER/mem[9][5][0] ) );
  dp_1 \ANSWER/mem_reg[9][6][0]  ( .ip(n3738), .ck(clk), .q(
        \ANSWER/mem[9][6][0] ) );
  dp_1 \ANSWER/mem_reg[9][7][0]  ( .ip(n3737), .ck(clk), .q(
        \ANSWER/mem[9][7][0] ) );
  dp_1 \ANSWER/mem_reg[9][8][0]  ( .ip(n3736), .ck(clk), .q(
        \ANSWER/mem[9][8][0] ) );
  dp_1 \ANSWER/mem_reg[9][9][0]  ( .ip(n3735), .ck(clk), .q(
        \ANSWER/mem[9][9][0] ) );
  dp_1 \SIGMOID/lut_out_reg[1]  ( .ip(n3841), .ck(clk), .q(
        \SIGMOID/lut_out [1]) );
  dp_1 \ANSWER/mem_reg[0][0][1]  ( .ip(n3734), .ck(clk), .q(
        \ANSWER/mem[0][0][1] ) );
  dp_1 \ANSWER/mem_reg[0][1][1]  ( .ip(n3733), .ck(clk), .q(
        \ANSWER/mem[0][1][1] ) );
  dp_1 \ANSWER/mem_reg[0][2][1]  ( .ip(n3732), .ck(clk), .q(
        \ANSWER/mem[0][2][1] ) );
  dp_1 \ANSWER/mem_reg[0][3][1]  ( .ip(n3731), .ck(clk), .q(
        \ANSWER/mem[0][3][1] ) );
  dp_1 \ANSWER/mem_reg[0][4][1]  ( .ip(n3730), .ck(clk), .q(
        \ANSWER/mem[0][4][1] ) );
  dp_1 \ANSWER/mem_reg[0][5][1]  ( .ip(n3729), .ck(clk), .q(
        \ANSWER/mem[0][5][1] ) );
  dp_1 \ANSWER/mem_reg[0][6][1]  ( .ip(n3728), .ck(clk), .q(
        \ANSWER/mem[0][6][1] ) );
  dp_1 \ANSWER/mem_reg[0][7][1]  ( .ip(n3727), .ck(clk), .q(
        \ANSWER/mem[0][7][1] ) );
  dp_1 \ANSWER/mem_reg[0][8][1]  ( .ip(n3726), .ck(clk), .q(
        \ANSWER/mem[0][8][1] ) );
  dp_1 \ANSWER/mem_reg[0][9][1]  ( .ip(n3725), .ck(clk), .q(
        \ANSWER/mem[0][9][1] ) );
  dp_1 \ANSWER/mem_reg[1][0][1]  ( .ip(n3724), .ck(clk), .q(
        \ANSWER/mem[1][0][1] ) );
  dp_1 \ANSWER/mem_reg[1][1][1]  ( .ip(n3723), .ck(clk), .q(
        \ANSWER/mem[1][1][1] ) );
  dp_1 \ANSWER/mem_reg[1][2][1]  ( .ip(n3722), .ck(clk), .q(
        \ANSWER/mem[1][2][1] ) );
  dp_1 \ANSWER/mem_reg[1][3][1]  ( .ip(n3721), .ck(clk), .q(
        \ANSWER/mem[1][3][1] ) );
  dp_1 \ANSWER/mem_reg[1][4][1]  ( .ip(n3720), .ck(clk), .q(
        \ANSWER/mem[1][4][1] ) );
  dp_1 \ANSWER/mem_reg[1][5][1]  ( .ip(n3719), .ck(clk), .q(
        \ANSWER/mem[1][5][1] ) );
  dp_1 \ANSWER/mem_reg[1][6][1]  ( .ip(n3718), .ck(clk), .q(
        \ANSWER/mem[1][6][1] ) );
  dp_1 \ANSWER/mem_reg[1][7][1]  ( .ip(n3717), .ck(clk), .q(
        \ANSWER/mem[1][7][1] ) );
  dp_1 \ANSWER/mem_reg[1][8][1]  ( .ip(n3716), .ck(clk), .q(
        \ANSWER/mem[1][8][1] ) );
  dp_1 \ANSWER/mem_reg[1][9][1]  ( .ip(n3715), .ck(clk), .q(
        \ANSWER/mem[1][9][1] ) );
  dp_1 \ANSWER/mem_reg[2][0][1]  ( .ip(n3714), .ck(clk), .q(
        \ANSWER/mem[2][0][1] ) );
  dp_1 \ANSWER/mem_reg[2][1][1]  ( .ip(n3713), .ck(clk), .q(
        \ANSWER/mem[2][1][1] ) );
  dp_1 \ANSWER/mem_reg[2][2][1]  ( .ip(n3712), .ck(clk), .q(
        \ANSWER/mem[2][2][1] ) );
  dp_1 \ANSWER/mem_reg[2][3][1]  ( .ip(n3711), .ck(clk), .q(
        \ANSWER/mem[2][3][1] ) );
  dp_1 \ANSWER/mem_reg[2][4][1]  ( .ip(n3710), .ck(clk), .q(
        \ANSWER/mem[2][4][1] ) );
  dp_1 \ANSWER/mem_reg[2][5][1]  ( .ip(n3709), .ck(clk), .q(
        \ANSWER/mem[2][5][1] ) );
  dp_1 \ANSWER/mem_reg[2][6][1]  ( .ip(n3708), .ck(clk), .q(
        \ANSWER/mem[2][6][1] ) );
  dp_1 \ANSWER/mem_reg[2][7][1]  ( .ip(n3707), .ck(clk), .q(
        \ANSWER/mem[2][7][1] ) );
  dp_1 \ANSWER/mem_reg[2][8][1]  ( .ip(n3706), .ck(clk), .q(
        \ANSWER/mem[2][8][1] ) );
  dp_1 \ANSWER/mem_reg[2][9][1]  ( .ip(n3705), .ck(clk), .q(
        \ANSWER/mem[2][9][1] ) );
  dp_1 \ANSWER/mem_reg[3][0][1]  ( .ip(n3704), .ck(clk), .q(
        \ANSWER/mem[3][0][1] ) );
  dp_1 \ANSWER/mem_reg[3][1][1]  ( .ip(n3703), .ck(clk), .q(
        \ANSWER/mem[3][1][1] ) );
  dp_1 \ANSWER/mem_reg[3][2][1]  ( .ip(n3702), .ck(clk), .q(
        \ANSWER/mem[3][2][1] ) );
  dp_1 \ANSWER/mem_reg[3][3][1]  ( .ip(n3701), .ck(clk), .q(
        \ANSWER/mem[3][3][1] ) );
  dp_1 \ANSWER/mem_reg[3][4][1]  ( .ip(n3700), .ck(clk), .q(
        \ANSWER/mem[3][4][1] ) );
  dp_1 \ANSWER/mem_reg[3][5][1]  ( .ip(n3699), .ck(clk), .q(
        \ANSWER/mem[3][5][1] ) );
  dp_1 \ANSWER/mem_reg[3][6][1]  ( .ip(n3698), .ck(clk), .q(
        \ANSWER/mem[3][6][1] ) );
  dp_1 \ANSWER/mem_reg[3][7][1]  ( .ip(n3697), .ck(clk), .q(
        \ANSWER/mem[3][7][1] ) );
  dp_1 \ANSWER/mem_reg[3][8][1]  ( .ip(n3696), .ck(clk), .q(
        \ANSWER/mem[3][8][1] ) );
  dp_1 \ANSWER/mem_reg[3][9][1]  ( .ip(n3695), .ck(clk), .q(
        \ANSWER/mem[3][9][1] ) );
  dp_1 \ANSWER/mem_reg[4][0][1]  ( .ip(n3694), .ck(clk), .q(
        \ANSWER/mem[4][0][1] ) );
  dp_1 \ANSWER/mem_reg[4][1][1]  ( .ip(n3693), .ck(clk), .q(
        \ANSWER/mem[4][1][1] ) );
  dp_1 \ANSWER/mem_reg[4][2][1]  ( .ip(n3692), .ck(clk), .q(
        \ANSWER/mem[4][2][1] ) );
  dp_1 \ANSWER/mem_reg[4][3][1]  ( .ip(n3691), .ck(clk), .q(
        \ANSWER/mem[4][3][1] ) );
  dp_1 \ANSWER/mem_reg[4][4][1]  ( .ip(n3690), .ck(clk), .q(
        \ANSWER/mem[4][4][1] ) );
  dp_1 \ANSWER/mem_reg[4][5][1]  ( .ip(n3689), .ck(clk), .q(
        \ANSWER/mem[4][5][1] ) );
  dp_1 \ANSWER/mem_reg[4][6][1]  ( .ip(n3688), .ck(clk), .q(
        \ANSWER/mem[4][6][1] ) );
  dp_1 \ANSWER/mem_reg[4][7][1]  ( .ip(n3687), .ck(clk), .q(
        \ANSWER/mem[4][7][1] ) );
  dp_1 \ANSWER/mem_reg[4][8][1]  ( .ip(n3686), .ck(clk), .q(
        \ANSWER/mem[4][8][1] ) );
  dp_1 \ANSWER/mem_reg[4][9][1]  ( .ip(n3685), .ck(clk), .q(
        \ANSWER/mem[4][9][1] ) );
  dp_1 \ANSWER/mem_reg[5][0][1]  ( .ip(n3684), .ck(clk), .q(
        \ANSWER/mem[5][0][1] ) );
  dp_1 \ANSWER/mem_reg[5][1][1]  ( .ip(n3683), .ck(clk), .q(
        \ANSWER/mem[5][1][1] ) );
  dp_1 \ANSWER/mem_reg[5][2][1]  ( .ip(n3682), .ck(clk), .q(
        \ANSWER/mem[5][2][1] ) );
  dp_1 \ANSWER/mem_reg[5][3][1]  ( .ip(n3681), .ck(clk), .q(
        \ANSWER/mem[5][3][1] ) );
  dp_1 \ANSWER/mem_reg[5][4][1]  ( .ip(n3680), .ck(clk), .q(
        \ANSWER/mem[5][4][1] ) );
  dp_1 \ANSWER/mem_reg[5][5][1]  ( .ip(n3679), .ck(clk), .q(
        \ANSWER/mem[5][5][1] ) );
  dp_1 \ANSWER/mem_reg[5][6][1]  ( .ip(n3678), .ck(clk), .q(
        \ANSWER/mem[5][6][1] ) );
  dp_1 \ANSWER/mem_reg[5][7][1]  ( .ip(n3677), .ck(clk), .q(
        \ANSWER/mem[5][7][1] ) );
  dp_1 \ANSWER/mem_reg[5][8][1]  ( .ip(n3676), .ck(clk), .q(
        \ANSWER/mem[5][8][1] ) );
  dp_1 \ANSWER/mem_reg[5][9][1]  ( .ip(n3675), .ck(clk), .q(
        \ANSWER/mem[5][9][1] ) );
  dp_1 \ANSWER/mem_reg[6][0][1]  ( .ip(n3674), .ck(clk), .q(
        \ANSWER/mem[6][0][1] ) );
  dp_1 \ANSWER/mem_reg[6][1][1]  ( .ip(n3673), .ck(clk), .q(
        \ANSWER/mem[6][1][1] ) );
  dp_1 \ANSWER/mem_reg[6][2][1]  ( .ip(n3672), .ck(clk), .q(
        \ANSWER/mem[6][2][1] ) );
  dp_1 \ANSWER/mem_reg[6][3][1]  ( .ip(n3671), .ck(clk), .q(
        \ANSWER/mem[6][3][1] ) );
  dp_1 \ANSWER/mem_reg[6][4][1]  ( .ip(n3670), .ck(clk), .q(
        \ANSWER/mem[6][4][1] ) );
  dp_1 \ANSWER/mem_reg[6][5][1]  ( .ip(n3669), .ck(clk), .q(
        \ANSWER/mem[6][5][1] ) );
  dp_1 \ANSWER/mem_reg[6][6][1]  ( .ip(n3668), .ck(clk), .q(
        \ANSWER/mem[6][6][1] ) );
  dp_1 \ANSWER/mem_reg[6][7][1]  ( .ip(n3667), .ck(clk), .q(
        \ANSWER/mem[6][7][1] ) );
  dp_1 \ANSWER/mem_reg[6][8][1]  ( .ip(n3666), .ck(clk), .q(
        \ANSWER/mem[6][8][1] ) );
  dp_1 \ANSWER/mem_reg[6][9][1]  ( .ip(n3665), .ck(clk), .q(
        \ANSWER/mem[6][9][1] ) );
  dp_1 \ANSWER/mem_reg[7][0][1]  ( .ip(n3664), .ck(clk), .q(
        \ANSWER/mem[7][0][1] ) );
  dp_1 \ANSWER/mem_reg[7][1][1]  ( .ip(n3663), .ck(clk), .q(
        \ANSWER/mem[7][1][1] ) );
  dp_1 \ANSWER/mem_reg[7][2][1]  ( .ip(n3662), .ck(clk), .q(
        \ANSWER/mem[7][2][1] ) );
  dp_1 \ANSWER/mem_reg[7][3][1]  ( .ip(n3661), .ck(clk), .q(
        \ANSWER/mem[7][3][1] ) );
  dp_1 \ANSWER/mem_reg[7][4][1]  ( .ip(n3660), .ck(clk), .q(
        \ANSWER/mem[7][4][1] ) );
  dp_1 \ANSWER/mem_reg[7][5][1]  ( .ip(n3659), .ck(clk), .q(
        \ANSWER/mem[7][5][1] ) );
  dp_1 \ANSWER/mem_reg[7][6][1]  ( .ip(n3658), .ck(clk), .q(
        \ANSWER/mem[7][6][1] ) );
  dp_1 \ANSWER/mem_reg[7][7][1]  ( .ip(n3657), .ck(clk), .q(
        \ANSWER/mem[7][7][1] ) );
  dp_1 \ANSWER/mem_reg[7][8][1]  ( .ip(n3656), .ck(clk), .q(
        \ANSWER/mem[7][8][1] ) );
  dp_1 \ANSWER/mem_reg[7][9][1]  ( .ip(n3655), .ck(clk), .q(
        \ANSWER/mem[7][9][1] ) );
  dp_1 \ANSWER/mem_reg[8][0][1]  ( .ip(n3654), .ck(clk), .q(
        \ANSWER/mem[8][0][1] ) );
  dp_1 \ANSWER/mem_reg[8][1][1]  ( .ip(n3653), .ck(clk), .q(
        \ANSWER/mem[8][1][1] ) );
  dp_1 \ANSWER/mem_reg[8][2][1]  ( .ip(n3652), .ck(clk), .q(
        \ANSWER/mem[8][2][1] ) );
  dp_1 \ANSWER/mem_reg[8][3][1]  ( .ip(n3651), .ck(clk), .q(
        \ANSWER/mem[8][3][1] ) );
  dp_1 \ANSWER/mem_reg[8][4][1]  ( .ip(n3650), .ck(clk), .q(
        \ANSWER/mem[8][4][1] ) );
  dp_1 \ANSWER/mem_reg[8][5][1]  ( .ip(n3649), .ck(clk), .q(
        \ANSWER/mem[8][5][1] ) );
  dp_1 \ANSWER/mem_reg[8][6][1]  ( .ip(n3648), .ck(clk), .q(
        \ANSWER/mem[8][6][1] ) );
  dp_1 \ANSWER/mem_reg[8][7][1]  ( .ip(n3647), .ck(clk), .q(
        \ANSWER/mem[8][7][1] ) );
  dp_1 \ANSWER/mem_reg[8][8][1]  ( .ip(n3646), .ck(clk), .q(
        \ANSWER/mem[8][8][1] ) );
  dp_1 \ANSWER/mem_reg[8][9][1]  ( .ip(n3645), .ck(clk), .q(
        \ANSWER/mem[8][9][1] ) );
  dp_1 \ANSWER/mem_reg[9][0][1]  ( .ip(n3644), .ck(clk), .q(
        \ANSWER/mem[9][0][1] ) );
  dp_1 \ANSWER/mem_reg[9][1][1]  ( .ip(n3643), .ck(clk), .q(
        \ANSWER/mem[9][1][1] ) );
  dp_1 \ANSWER/mem_reg[9][2][1]  ( .ip(n3642), .ck(clk), .q(
        \ANSWER/mem[9][2][1] ) );
  dp_1 \ANSWER/mem_reg[9][3][1]  ( .ip(n3641), .ck(clk), .q(
        \ANSWER/mem[9][3][1] ) );
  dp_1 \ANSWER/mem_reg[9][4][1]  ( .ip(n3640), .ck(clk), .q(
        \ANSWER/mem[9][4][1] ) );
  dp_1 \ANSWER/mem_reg[9][5][1]  ( .ip(n3639), .ck(clk), .q(
        \ANSWER/mem[9][5][1] ) );
  dp_1 \ANSWER/mem_reg[9][6][1]  ( .ip(n3638), .ck(clk), .q(
        \ANSWER/mem[9][6][1] ) );
  dp_1 \ANSWER/mem_reg[9][7][1]  ( .ip(n3637), .ck(clk), .q(
        \ANSWER/mem[9][7][1] ) );
  dp_1 \ANSWER/mem_reg[9][8][1]  ( .ip(n3636), .ck(clk), .q(
        \ANSWER/mem[9][8][1] ) );
  dp_1 \ANSWER/mem_reg[9][9][1]  ( .ip(n3635), .ck(clk), .q(
        \ANSWER/mem[9][9][1] ) );
  dp_1 \SIGMOID/lut_out_reg[2]  ( .ip(n3840), .ck(clk), .q(
        \SIGMOID/lut_out [2]) );
  dp_1 \ANSWER/mem_reg[0][0][2]  ( .ip(n3634), .ck(clk), .q(
        \ANSWER/mem[0][0][2] ) );
  dp_1 \ANSWER/mem_reg[0][1][2]  ( .ip(n3633), .ck(clk), .q(
        \ANSWER/mem[0][1][2] ) );
  dp_1 \ANSWER/mem_reg[0][2][2]  ( .ip(n3632), .ck(clk), .q(
        \ANSWER/mem[0][2][2] ) );
  dp_1 \ANSWER/mem_reg[0][3][2]  ( .ip(n3631), .ck(clk), .q(
        \ANSWER/mem[0][3][2] ) );
  dp_1 \ANSWER/mem_reg[0][4][2]  ( .ip(n3630), .ck(clk), .q(
        \ANSWER/mem[0][4][2] ) );
  dp_1 \ANSWER/mem_reg[0][5][2]  ( .ip(n3629), .ck(clk), .q(
        \ANSWER/mem[0][5][2] ) );
  dp_1 \ANSWER/mem_reg[0][6][2]  ( .ip(n3628), .ck(clk), .q(
        \ANSWER/mem[0][6][2] ) );
  dp_1 \ANSWER/mem_reg[0][7][2]  ( .ip(n3627), .ck(clk), .q(
        \ANSWER/mem[0][7][2] ) );
  dp_1 \ANSWER/mem_reg[0][8][2]  ( .ip(n3626), .ck(clk), .q(
        \ANSWER/mem[0][8][2] ) );
  dp_1 \ANSWER/mem_reg[0][9][2]  ( .ip(n3625), .ck(clk), .q(
        \ANSWER/mem[0][9][2] ) );
  dp_1 \ANSWER/mem_reg[1][0][2]  ( .ip(n3624), .ck(clk), .q(
        \ANSWER/mem[1][0][2] ) );
  dp_1 \ANSWER/mem_reg[1][1][2]  ( .ip(n3623), .ck(clk), .q(
        \ANSWER/mem[1][1][2] ) );
  dp_1 \ANSWER/mem_reg[1][2][2]  ( .ip(n3622), .ck(clk), .q(
        \ANSWER/mem[1][2][2] ) );
  dp_1 \ANSWER/mem_reg[1][3][2]  ( .ip(n3621), .ck(clk), .q(
        \ANSWER/mem[1][3][2] ) );
  dp_1 \ANSWER/mem_reg[1][4][2]  ( .ip(n3620), .ck(clk), .q(
        \ANSWER/mem[1][4][2] ) );
  dp_1 \ANSWER/mem_reg[1][5][2]  ( .ip(n3619), .ck(clk), .q(
        \ANSWER/mem[1][5][2] ) );
  dp_1 \ANSWER/mem_reg[1][6][2]  ( .ip(n3618), .ck(clk), .q(
        \ANSWER/mem[1][6][2] ) );
  dp_1 \ANSWER/mem_reg[1][7][2]  ( .ip(n3617), .ck(clk), .q(
        \ANSWER/mem[1][7][2] ) );
  dp_1 \ANSWER/mem_reg[1][8][2]  ( .ip(n3616), .ck(clk), .q(
        \ANSWER/mem[1][8][2] ) );
  dp_1 \ANSWER/mem_reg[1][9][2]  ( .ip(n3615), .ck(clk), .q(
        \ANSWER/mem[1][9][2] ) );
  dp_1 \ANSWER/mem_reg[2][0][2]  ( .ip(n3614), .ck(clk), .q(
        \ANSWER/mem[2][0][2] ) );
  dp_1 \ANSWER/mem_reg[2][1][2]  ( .ip(n3613), .ck(clk), .q(
        \ANSWER/mem[2][1][2] ) );
  dp_1 \ANSWER/mem_reg[2][2][2]  ( .ip(n3612), .ck(clk), .q(
        \ANSWER/mem[2][2][2] ) );
  dp_1 \ANSWER/mem_reg[2][3][2]  ( .ip(n3611), .ck(clk), .q(
        \ANSWER/mem[2][3][2] ) );
  dp_1 \ANSWER/mem_reg[2][4][2]  ( .ip(n3610), .ck(clk), .q(
        \ANSWER/mem[2][4][2] ) );
  dp_1 \ANSWER/mem_reg[2][5][2]  ( .ip(n3609), .ck(clk), .q(
        \ANSWER/mem[2][5][2] ) );
  dp_1 \ANSWER/mem_reg[2][6][2]  ( .ip(n3608), .ck(clk), .q(
        \ANSWER/mem[2][6][2] ) );
  dp_1 \ANSWER/mem_reg[2][7][2]  ( .ip(n3607), .ck(clk), .q(
        \ANSWER/mem[2][7][2] ) );
  dp_1 \ANSWER/mem_reg[2][8][2]  ( .ip(n3606), .ck(clk), .q(
        \ANSWER/mem[2][8][2] ) );
  dp_1 \ANSWER/mem_reg[2][9][2]  ( .ip(n3605), .ck(clk), .q(
        \ANSWER/mem[2][9][2] ) );
  dp_1 \ANSWER/mem_reg[3][0][2]  ( .ip(n3604), .ck(clk), .q(
        \ANSWER/mem[3][0][2] ) );
  dp_1 \ANSWER/mem_reg[3][1][2]  ( .ip(n3603), .ck(clk), .q(
        \ANSWER/mem[3][1][2] ) );
  dp_1 \ANSWER/mem_reg[3][2][2]  ( .ip(n3602), .ck(clk), .q(
        \ANSWER/mem[3][2][2] ) );
  dp_1 \ANSWER/mem_reg[3][3][2]  ( .ip(n3601), .ck(clk), .q(
        \ANSWER/mem[3][3][2] ) );
  dp_1 \ANSWER/mem_reg[3][4][2]  ( .ip(n3600), .ck(clk), .q(
        \ANSWER/mem[3][4][2] ) );
  dp_1 \ANSWER/mem_reg[3][5][2]  ( .ip(n3599), .ck(clk), .q(
        \ANSWER/mem[3][5][2] ) );
  dp_1 \ANSWER/mem_reg[3][6][2]  ( .ip(n3598), .ck(clk), .q(
        \ANSWER/mem[3][6][2] ) );
  dp_1 \ANSWER/mem_reg[3][7][2]  ( .ip(n3597), .ck(clk), .q(
        \ANSWER/mem[3][7][2] ) );
  dp_1 \ANSWER/mem_reg[3][8][2]  ( .ip(n3596), .ck(clk), .q(
        \ANSWER/mem[3][8][2] ) );
  dp_1 \ANSWER/mem_reg[3][9][2]  ( .ip(n3595), .ck(clk), .q(
        \ANSWER/mem[3][9][2] ) );
  dp_1 \ANSWER/mem_reg[4][0][2]  ( .ip(n3594), .ck(clk), .q(
        \ANSWER/mem[4][0][2] ) );
  dp_1 \ANSWER/mem_reg[4][1][2]  ( .ip(n3593), .ck(clk), .q(
        \ANSWER/mem[4][1][2] ) );
  dp_1 \ANSWER/mem_reg[4][2][2]  ( .ip(n3592), .ck(clk), .q(
        \ANSWER/mem[4][2][2] ) );
  dp_1 \ANSWER/mem_reg[4][3][2]  ( .ip(n3591), .ck(clk), .q(
        \ANSWER/mem[4][3][2] ) );
  dp_1 \ANSWER/mem_reg[4][4][2]  ( .ip(n3590), .ck(clk), .q(
        \ANSWER/mem[4][4][2] ) );
  dp_1 \ANSWER/mem_reg[4][5][2]  ( .ip(n3589), .ck(clk), .q(
        \ANSWER/mem[4][5][2] ) );
  dp_1 \ANSWER/mem_reg[4][6][2]  ( .ip(n3588), .ck(clk), .q(
        \ANSWER/mem[4][6][2] ) );
  dp_1 \ANSWER/mem_reg[4][7][2]  ( .ip(n3587), .ck(clk), .q(
        \ANSWER/mem[4][7][2] ) );
  dp_1 \ANSWER/mem_reg[4][8][2]  ( .ip(n3586), .ck(clk), .q(
        \ANSWER/mem[4][8][2] ) );
  dp_1 \ANSWER/mem_reg[4][9][2]  ( .ip(n3585), .ck(clk), .q(
        \ANSWER/mem[4][9][2] ) );
  dp_1 \ANSWER/mem_reg[5][0][2]  ( .ip(n3584), .ck(clk), .q(
        \ANSWER/mem[5][0][2] ) );
  dp_1 \ANSWER/mem_reg[5][1][2]  ( .ip(n3583), .ck(clk), .q(
        \ANSWER/mem[5][1][2] ) );
  dp_1 \ANSWER/mem_reg[5][2][2]  ( .ip(n3582), .ck(clk), .q(
        \ANSWER/mem[5][2][2] ) );
  dp_1 \ANSWER/mem_reg[5][3][2]  ( .ip(n3581), .ck(clk), .q(
        \ANSWER/mem[5][3][2] ) );
  dp_1 \ANSWER/mem_reg[5][4][2]  ( .ip(n3580), .ck(clk), .q(
        \ANSWER/mem[5][4][2] ) );
  dp_1 \ANSWER/mem_reg[5][5][2]  ( .ip(n3579), .ck(clk), .q(
        \ANSWER/mem[5][5][2] ) );
  dp_1 \ANSWER/mem_reg[5][6][2]  ( .ip(n3578), .ck(clk), .q(
        \ANSWER/mem[5][6][2] ) );
  dp_1 \ANSWER/mem_reg[5][7][2]  ( .ip(n3577), .ck(clk), .q(
        \ANSWER/mem[5][7][2] ) );
  dp_1 \ANSWER/mem_reg[5][8][2]  ( .ip(n3576), .ck(clk), .q(
        \ANSWER/mem[5][8][2] ) );
  dp_1 \ANSWER/mem_reg[5][9][2]  ( .ip(n3575), .ck(clk), .q(
        \ANSWER/mem[5][9][2] ) );
  dp_1 \ANSWER/mem_reg[6][0][2]  ( .ip(n3574), .ck(clk), .q(
        \ANSWER/mem[6][0][2] ) );
  dp_1 \ANSWER/mem_reg[6][1][2]  ( .ip(n3573), .ck(clk), .q(
        \ANSWER/mem[6][1][2] ) );
  dp_1 \ANSWER/mem_reg[6][2][2]  ( .ip(n3572), .ck(clk), .q(
        \ANSWER/mem[6][2][2] ) );
  dp_1 \ANSWER/mem_reg[6][3][2]  ( .ip(n3571), .ck(clk), .q(
        \ANSWER/mem[6][3][2] ) );
  dp_1 \ANSWER/mem_reg[6][4][2]  ( .ip(n3570), .ck(clk), .q(
        \ANSWER/mem[6][4][2] ) );
  dp_1 \ANSWER/mem_reg[6][5][2]  ( .ip(n3569), .ck(clk), .q(
        \ANSWER/mem[6][5][2] ) );
  dp_1 \ANSWER/mem_reg[6][6][2]  ( .ip(n3568), .ck(clk), .q(
        \ANSWER/mem[6][6][2] ) );
  dp_1 \ANSWER/mem_reg[6][7][2]  ( .ip(n3567), .ck(clk), .q(
        \ANSWER/mem[6][7][2] ) );
  dp_1 \ANSWER/mem_reg[6][8][2]  ( .ip(n3566), .ck(clk), .q(
        \ANSWER/mem[6][8][2] ) );
  dp_1 \ANSWER/mem_reg[6][9][2]  ( .ip(n3565), .ck(clk), .q(
        \ANSWER/mem[6][9][2] ) );
  dp_1 \ANSWER/mem_reg[7][0][2]  ( .ip(n3564), .ck(clk), .q(
        \ANSWER/mem[7][0][2] ) );
  dp_1 \ANSWER/mem_reg[7][1][2]  ( .ip(n3563), .ck(clk), .q(
        \ANSWER/mem[7][1][2] ) );
  dp_1 \ANSWER/mem_reg[7][2][2]  ( .ip(n3562), .ck(clk), .q(
        \ANSWER/mem[7][2][2] ) );
  dp_1 \ANSWER/mem_reg[7][3][2]  ( .ip(n3561), .ck(clk), .q(
        \ANSWER/mem[7][3][2] ) );
  dp_1 \ANSWER/mem_reg[7][4][2]  ( .ip(n3560), .ck(clk), .q(
        \ANSWER/mem[7][4][2] ) );
  dp_1 \ANSWER/mem_reg[7][5][2]  ( .ip(n3559), .ck(clk), .q(
        \ANSWER/mem[7][5][2] ) );
  dp_1 \ANSWER/mem_reg[7][6][2]  ( .ip(n3558), .ck(clk), .q(
        \ANSWER/mem[7][6][2] ) );
  dp_1 \ANSWER/mem_reg[7][7][2]  ( .ip(n3557), .ck(clk), .q(
        \ANSWER/mem[7][7][2] ) );
  dp_1 \ANSWER/mem_reg[7][8][2]  ( .ip(n3556), .ck(clk), .q(
        \ANSWER/mem[7][8][2] ) );
  dp_1 \ANSWER/mem_reg[7][9][2]  ( .ip(n3555), .ck(clk), .q(
        \ANSWER/mem[7][9][2] ) );
  dp_1 \ANSWER/mem_reg[8][0][2]  ( .ip(n3554), .ck(clk), .q(
        \ANSWER/mem[8][0][2] ) );
  dp_1 \ANSWER/mem_reg[8][1][2]  ( .ip(n3553), .ck(clk), .q(
        \ANSWER/mem[8][1][2] ) );
  dp_1 \ANSWER/mem_reg[8][2][2]  ( .ip(n3552), .ck(clk), .q(
        \ANSWER/mem[8][2][2] ) );
  dp_1 \ANSWER/mem_reg[8][3][2]  ( .ip(n3551), .ck(clk), .q(
        \ANSWER/mem[8][3][2] ) );
  dp_1 \ANSWER/mem_reg[8][4][2]  ( .ip(n3550), .ck(clk), .q(
        \ANSWER/mem[8][4][2] ) );
  dp_1 \ANSWER/mem_reg[8][5][2]  ( .ip(n3549), .ck(clk), .q(
        \ANSWER/mem[8][5][2] ) );
  dp_1 \ANSWER/mem_reg[8][6][2]  ( .ip(n3548), .ck(clk), .q(
        \ANSWER/mem[8][6][2] ) );
  dp_1 \ANSWER/mem_reg[8][7][2]  ( .ip(n3547), .ck(clk), .q(
        \ANSWER/mem[8][7][2] ) );
  dp_1 \ANSWER/mem_reg[8][8][2]  ( .ip(n3546), .ck(clk), .q(
        \ANSWER/mem[8][8][2] ) );
  dp_1 \ANSWER/mem_reg[8][9][2]  ( .ip(n3545), .ck(clk), .q(
        \ANSWER/mem[8][9][2] ) );
  dp_1 \ANSWER/mem_reg[9][0][2]  ( .ip(n3544), .ck(clk), .q(
        \ANSWER/mem[9][0][2] ) );
  dp_1 \ANSWER/mem_reg[9][1][2]  ( .ip(n3543), .ck(clk), .q(
        \ANSWER/mem[9][1][2] ) );
  dp_1 \ANSWER/mem_reg[9][2][2]  ( .ip(n3542), .ck(clk), .q(
        \ANSWER/mem[9][2][2] ) );
  dp_1 \ANSWER/mem_reg[9][3][2]  ( .ip(n3541), .ck(clk), .q(
        \ANSWER/mem[9][3][2] ) );
  dp_1 \ANSWER/mem_reg[9][4][2]  ( .ip(n3540), .ck(clk), .q(
        \ANSWER/mem[9][4][2] ) );
  dp_1 \ANSWER/mem_reg[9][5][2]  ( .ip(n3539), .ck(clk), .q(
        \ANSWER/mem[9][5][2] ) );
  dp_1 \ANSWER/mem_reg[9][6][2]  ( .ip(n3538), .ck(clk), .q(
        \ANSWER/mem[9][6][2] ) );
  dp_1 \ANSWER/mem_reg[9][7][2]  ( .ip(n3537), .ck(clk), .q(
        \ANSWER/mem[9][7][2] ) );
  dp_1 \ANSWER/mem_reg[9][8][2]  ( .ip(n3536), .ck(clk), .q(
        \ANSWER/mem[9][8][2] ) );
  dp_1 \ANSWER/mem_reg[9][9][2]  ( .ip(n3535), .ck(clk), .q(
        \ANSWER/mem[9][9][2] ) );
  dp_1 \SIGMOID/lut_out_reg[3]  ( .ip(n3839), .ck(clk), .q(
        \SIGMOID/lut_out [3]) );
  dp_1 \ANSWER/mem_reg[0][0][3]  ( .ip(n3534), .ck(clk), .q(
        \ANSWER/mem[0][0][3] ) );
  dp_1 \ANSWER/mem_reg[0][1][3]  ( .ip(n3533), .ck(clk), .q(
        \ANSWER/mem[0][1][3] ) );
  dp_1 \ANSWER/mem_reg[0][2][3]  ( .ip(n3532), .ck(clk), .q(
        \ANSWER/mem[0][2][3] ) );
  dp_1 \ANSWER/mem_reg[0][3][3]  ( .ip(n3531), .ck(clk), .q(
        \ANSWER/mem[0][3][3] ) );
  dp_1 \ANSWER/mem_reg[0][4][3]  ( .ip(n3530), .ck(clk), .q(
        \ANSWER/mem[0][4][3] ) );
  dp_1 \ANSWER/mem_reg[0][5][3]  ( .ip(n3529), .ck(clk), .q(
        \ANSWER/mem[0][5][3] ) );
  dp_1 \ANSWER/mem_reg[0][6][3]  ( .ip(n3528), .ck(clk), .q(
        \ANSWER/mem[0][6][3] ) );
  dp_1 \ANSWER/mem_reg[0][7][3]  ( .ip(n3527), .ck(clk), .q(
        \ANSWER/mem[0][7][3] ) );
  dp_1 \ANSWER/mem_reg[0][8][3]  ( .ip(n3526), .ck(clk), .q(
        \ANSWER/mem[0][8][3] ) );
  dp_1 \ANSWER/mem_reg[0][9][3]  ( .ip(n3525), .ck(clk), .q(
        \ANSWER/mem[0][9][3] ) );
  dp_1 \ANSWER/mem_reg[1][0][3]  ( .ip(n3524), .ck(clk), .q(
        \ANSWER/mem[1][0][3] ) );
  dp_1 \ANSWER/mem_reg[1][1][3]  ( .ip(n3523), .ck(clk), .q(
        \ANSWER/mem[1][1][3] ) );
  dp_1 \ANSWER/mem_reg[1][2][3]  ( .ip(n3522), .ck(clk), .q(
        \ANSWER/mem[1][2][3] ) );
  dp_1 \ANSWER/mem_reg[1][3][3]  ( .ip(n3521), .ck(clk), .q(
        \ANSWER/mem[1][3][3] ) );
  dp_1 \ANSWER/mem_reg[1][4][3]  ( .ip(n3520), .ck(clk), .q(
        \ANSWER/mem[1][4][3] ) );
  dp_1 \ANSWER/mem_reg[1][5][3]  ( .ip(n3519), .ck(clk), .q(
        \ANSWER/mem[1][5][3] ) );
  dp_1 \ANSWER/mem_reg[1][6][3]  ( .ip(n3518), .ck(clk), .q(
        \ANSWER/mem[1][6][3] ) );
  dp_1 \ANSWER/mem_reg[1][7][3]  ( .ip(n3517), .ck(clk), .q(
        \ANSWER/mem[1][7][3] ) );
  dp_1 \ANSWER/mem_reg[1][8][3]  ( .ip(n3516), .ck(clk), .q(
        \ANSWER/mem[1][8][3] ) );
  dp_1 \ANSWER/mem_reg[1][9][3]  ( .ip(n3515), .ck(clk), .q(
        \ANSWER/mem[1][9][3] ) );
  dp_1 \ANSWER/mem_reg[2][0][3]  ( .ip(n3514), .ck(clk), .q(
        \ANSWER/mem[2][0][3] ) );
  dp_1 \ANSWER/mem_reg[2][1][3]  ( .ip(n3513), .ck(clk), .q(
        \ANSWER/mem[2][1][3] ) );
  dp_1 \ANSWER/mem_reg[2][2][3]  ( .ip(n3512), .ck(clk), .q(
        \ANSWER/mem[2][2][3] ) );
  dp_1 \ANSWER/mem_reg[2][3][3]  ( .ip(n3511), .ck(clk), .q(
        \ANSWER/mem[2][3][3] ) );
  dp_1 \ANSWER/mem_reg[2][4][3]  ( .ip(n3510), .ck(clk), .q(
        \ANSWER/mem[2][4][3] ) );
  dp_1 \ANSWER/mem_reg[2][5][3]  ( .ip(n3509), .ck(clk), .q(
        \ANSWER/mem[2][5][3] ) );
  dp_1 \ANSWER/mem_reg[2][6][3]  ( .ip(n3508), .ck(clk), .q(
        \ANSWER/mem[2][6][3] ) );
  dp_1 \ANSWER/mem_reg[2][7][3]  ( .ip(n3507), .ck(clk), .q(
        \ANSWER/mem[2][7][3] ) );
  dp_1 \ANSWER/mem_reg[2][8][3]  ( .ip(n3506), .ck(clk), .q(
        \ANSWER/mem[2][8][3] ) );
  dp_1 \ANSWER/mem_reg[2][9][3]  ( .ip(n3505), .ck(clk), .q(
        \ANSWER/mem[2][9][3] ) );
  dp_1 \ANSWER/mem_reg[3][0][3]  ( .ip(n3504), .ck(clk), .q(
        \ANSWER/mem[3][0][3] ) );
  dp_1 \ANSWER/mem_reg[3][1][3]  ( .ip(n3503), .ck(clk), .q(
        \ANSWER/mem[3][1][3] ) );
  dp_1 \ANSWER/mem_reg[3][2][3]  ( .ip(n3502), .ck(clk), .q(
        \ANSWER/mem[3][2][3] ) );
  dp_1 \ANSWER/mem_reg[3][3][3]  ( .ip(n3501), .ck(clk), .q(
        \ANSWER/mem[3][3][3] ) );
  dp_1 \ANSWER/mem_reg[3][4][3]  ( .ip(n3500), .ck(clk), .q(
        \ANSWER/mem[3][4][3] ) );
  dp_1 \ANSWER/mem_reg[3][5][3]  ( .ip(n3499), .ck(clk), .q(
        \ANSWER/mem[3][5][3] ) );
  dp_1 \ANSWER/mem_reg[3][6][3]  ( .ip(n3498), .ck(clk), .q(
        \ANSWER/mem[3][6][3] ) );
  dp_1 \ANSWER/mem_reg[3][7][3]  ( .ip(n3497), .ck(clk), .q(
        \ANSWER/mem[3][7][3] ) );
  dp_1 \ANSWER/mem_reg[3][8][3]  ( .ip(n3496), .ck(clk), .q(
        \ANSWER/mem[3][8][3] ) );
  dp_1 \ANSWER/mem_reg[3][9][3]  ( .ip(n3495), .ck(clk), .q(
        \ANSWER/mem[3][9][3] ) );
  dp_1 \ANSWER/mem_reg[4][0][3]  ( .ip(n3494), .ck(clk), .q(
        \ANSWER/mem[4][0][3] ) );
  dp_1 \ANSWER/mem_reg[4][1][3]  ( .ip(n3493), .ck(clk), .q(
        \ANSWER/mem[4][1][3] ) );
  dp_1 \ANSWER/mem_reg[4][2][3]  ( .ip(n3492), .ck(clk), .q(
        \ANSWER/mem[4][2][3] ) );
  dp_1 \ANSWER/mem_reg[4][3][3]  ( .ip(n3491), .ck(clk), .q(
        \ANSWER/mem[4][3][3] ) );
  dp_1 \ANSWER/mem_reg[4][4][3]  ( .ip(n3490), .ck(clk), .q(
        \ANSWER/mem[4][4][3] ) );
  dp_1 \ANSWER/mem_reg[4][5][3]  ( .ip(n3489), .ck(clk), .q(
        \ANSWER/mem[4][5][3] ) );
  dp_1 \ANSWER/mem_reg[4][6][3]  ( .ip(n3488), .ck(clk), .q(
        \ANSWER/mem[4][6][3] ) );
  dp_1 \ANSWER/mem_reg[4][7][3]  ( .ip(n3487), .ck(clk), .q(
        \ANSWER/mem[4][7][3] ) );
  dp_1 \ANSWER/mem_reg[4][8][3]  ( .ip(n3486), .ck(clk), .q(
        \ANSWER/mem[4][8][3] ) );
  dp_1 \ANSWER/mem_reg[4][9][3]  ( .ip(n3485), .ck(clk), .q(
        \ANSWER/mem[4][9][3] ) );
  dp_1 \ANSWER/mem_reg[5][0][3]  ( .ip(n3484), .ck(clk), .q(
        \ANSWER/mem[5][0][3] ) );
  dp_1 \ANSWER/mem_reg[5][1][3]  ( .ip(n3483), .ck(clk), .q(
        \ANSWER/mem[5][1][3] ) );
  dp_1 \ANSWER/mem_reg[5][2][3]  ( .ip(n3482), .ck(clk), .q(
        \ANSWER/mem[5][2][3] ) );
  dp_1 \ANSWER/mem_reg[5][3][3]  ( .ip(n3481), .ck(clk), .q(
        \ANSWER/mem[5][3][3] ) );
  dp_1 \ANSWER/mem_reg[5][4][3]  ( .ip(n3480), .ck(clk), .q(
        \ANSWER/mem[5][4][3] ) );
  dp_1 \ANSWER/mem_reg[5][5][3]  ( .ip(n3479), .ck(clk), .q(
        \ANSWER/mem[5][5][3] ) );
  dp_1 \ANSWER/mem_reg[5][6][3]  ( .ip(n3478), .ck(clk), .q(
        \ANSWER/mem[5][6][3] ) );
  dp_1 \ANSWER/mem_reg[5][7][3]  ( .ip(n3477), .ck(clk), .q(
        \ANSWER/mem[5][7][3] ) );
  dp_1 \ANSWER/mem_reg[5][8][3]  ( .ip(n3476), .ck(clk), .q(
        \ANSWER/mem[5][8][3] ) );
  dp_1 \ANSWER/mem_reg[5][9][3]  ( .ip(n3475), .ck(clk), .q(
        \ANSWER/mem[5][9][3] ) );
  dp_1 \ANSWER/mem_reg[6][0][3]  ( .ip(n3474), .ck(clk), .q(
        \ANSWER/mem[6][0][3] ) );
  dp_1 \ANSWER/mem_reg[6][1][3]  ( .ip(n3473), .ck(clk), .q(
        \ANSWER/mem[6][1][3] ) );
  dp_1 \ANSWER/mem_reg[6][2][3]  ( .ip(n3472), .ck(clk), .q(
        \ANSWER/mem[6][2][3] ) );
  dp_1 \ANSWER/mem_reg[6][3][3]  ( .ip(n3471), .ck(clk), .q(
        \ANSWER/mem[6][3][3] ) );
  dp_1 \ANSWER/mem_reg[6][4][3]  ( .ip(n3470), .ck(clk), .q(
        \ANSWER/mem[6][4][3] ) );
  dp_1 \ANSWER/mem_reg[6][5][3]  ( .ip(n3469), .ck(clk), .q(
        \ANSWER/mem[6][5][3] ) );
  dp_1 \ANSWER/mem_reg[6][6][3]  ( .ip(n3468), .ck(clk), .q(
        \ANSWER/mem[6][6][3] ) );
  dp_1 \ANSWER/mem_reg[6][7][3]  ( .ip(n3467), .ck(clk), .q(
        \ANSWER/mem[6][7][3] ) );
  dp_1 \ANSWER/mem_reg[6][8][3]  ( .ip(n3466), .ck(clk), .q(
        \ANSWER/mem[6][8][3] ) );
  dp_1 \ANSWER/mem_reg[6][9][3]  ( .ip(n3465), .ck(clk), .q(
        \ANSWER/mem[6][9][3] ) );
  dp_1 \ANSWER/mem_reg[7][0][3]  ( .ip(n3464), .ck(clk), .q(
        \ANSWER/mem[7][0][3] ) );
  dp_1 \ANSWER/mem_reg[7][1][3]  ( .ip(n3463), .ck(clk), .q(
        \ANSWER/mem[7][1][3] ) );
  dp_1 \ANSWER/mem_reg[7][2][3]  ( .ip(n3462), .ck(clk), .q(
        \ANSWER/mem[7][2][3] ) );
  dp_1 \ANSWER/mem_reg[7][3][3]  ( .ip(n3461), .ck(clk), .q(
        \ANSWER/mem[7][3][3] ) );
  dp_1 \ANSWER/mem_reg[7][4][3]  ( .ip(n3460), .ck(clk), .q(
        \ANSWER/mem[7][4][3] ) );
  dp_1 \ANSWER/mem_reg[7][5][3]  ( .ip(n3459), .ck(clk), .q(
        \ANSWER/mem[7][5][3] ) );
  dp_1 \ANSWER/mem_reg[7][6][3]  ( .ip(n3458), .ck(clk), .q(
        \ANSWER/mem[7][6][3] ) );
  dp_1 \ANSWER/mem_reg[7][7][3]  ( .ip(n3457), .ck(clk), .q(
        \ANSWER/mem[7][7][3] ) );
  dp_1 \ANSWER/mem_reg[7][8][3]  ( .ip(n3456), .ck(clk), .q(
        \ANSWER/mem[7][8][3] ) );
  dp_1 \ANSWER/mem_reg[7][9][3]  ( .ip(n3455), .ck(clk), .q(
        \ANSWER/mem[7][9][3] ) );
  dp_1 \ANSWER/mem_reg[8][0][3]  ( .ip(n3454), .ck(clk), .q(
        \ANSWER/mem[8][0][3] ) );
  dp_1 \ANSWER/mem_reg[8][1][3]  ( .ip(n3453), .ck(clk), .q(
        \ANSWER/mem[8][1][3] ) );
  dp_1 \ANSWER/mem_reg[8][2][3]  ( .ip(n3452), .ck(clk), .q(
        \ANSWER/mem[8][2][3] ) );
  dp_1 \ANSWER/mem_reg[8][3][3]  ( .ip(n3451), .ck(clk), .q(
        \ANSWER/mem[8][3][3] ) );
  dp_1 \ANSWER/mem_reg[8][4][3]  ( .ip(n3450), .ck(clk), .q(
        \ANSWER/mem[8][4][3] ) );
  dp_1 \ANSWER/mem_reg[8][5][3]  ( .ip(n3449), .ck(clk), .q(
        \ANSWER/mem[8][5][3] ) );
  dp_1 \ANSWER/mem_reg[8][6][3]  ( .ip(n3448), .ck(clk), .q(
        \ANSWER/mem[8][6][3] ) );
  dp_1 \ANSWER/mem_reg[8][7][3]  ( .ip(n3447), .ck(clk), .q(
        \ANSWER/mem[8][7][3] ) );
  dp_1 \ANSWER/mem_reg[8][8][3]  ( .ip(n3446), .ck(clk), .q(
        \ANSWER/mem[8][8][3] ) );
  dp_1 \ANSWER/mem_reg[8][9][3]  ( .ip(n3445), .ck(clk), .q(
        \ANSWER/mem[8][9][3] ) );
  dp_1 \ANSWER/mem_reg[9][0][3]  ( .ip(n3444), .ck(clk), .q(
        \ANSWER/mem[9][0][3] ) );
  dp_1 \ANSWER/mem_reg[9][1][3]  ( .ip(n3443), .ck(clk), .q(
        \ANSWER/mem[9][1][3] ) );
  dp_1 \ANSWER/mem_reg[9][2][3]  ( .ip(n3442), .ck(clk), .q(
        \ANSWER/mem[9][2][3] ) );
  dp_1 \ANSWER/mem_reg[9][3][3]  ( .ip(n3441), .ck(clk), .q(
        \ANSWER/mem[9][3][3] ) );
  dp_1 \ANSWER/mem_reg[9][4][3]  ( .ip(n3440), .ck(clk), .q(
        \ANSWER/mem[9][4][3] ) );
  dp_1 \ANSWER/mem_reg[9][5][3]  ( .ip(n3439), .ck(clk), .q(
        \ANSWER/mem[9][5][3] ) );
  dp_1 \ANSWER/mem_reg[9][6][3]  ( .ip(n3438), .ck(clk), .q(
        \ANSWER/mem[9][6][3] ) );
  dp_1 \ANSWER/mem_reg[9][7][3]  ( .ip(n3437), .ck(clk), .q(
        \ANSWER/mem[9][7][3] ) );
  dp_1 \ANSWER/mem_reg[9][8][3]  ( .ip(n3436), .ck(clk), .q(
        \ANSWER/mem[9][8][3] ) );
  dp_1 \ANSWER/mem_reg[9][9][3]  ( .ip(n3435), .ck(clk), .q(
        \ANSWER/mem[9][9][3] ) );
  dp_1 \SIGMOID/lut_out_reg[4]  ( .ip(n3838), .ck(clk), .q(
        \SIGMOID/lut_out [4]) );
  dp_1 \ANSWER/mem_reg[0][0][4]  ( .ip(n3434), .ck(clk), .q(
        \ANSWER/mem[0][0][4] ) );
  dp_1 \ANSWER/mem_reg[0][1][4]  ( .ip(n3433), .ck(clk), .q(
        \ANSWER/mem[0][1][4] ) );
  dp_1 \ANSWER/mem_reg[0][2][4]  ( .ip(n3432), .ck(clk), .q(
        \ANSWER/mem[0][2][4] ) );
  dp_1 \ANSWER/mem_reg[0][3][4]  ( .ip(n3431), .ck(clk), .q(
        \ANSWER/mem[0][3][4] ) );
  dp_1 \ANSWER/mem_reg[0][4][4]  ( .ip(n3430), .ck(clk), .q(
        \ANSWER/mem[0][4][4] ) );
  dp_1 \ANSWER/mem_reg[0][5][4]  ( .ip(n3429), .ck(clk), .q(
        \ANSWER/mem[0][5][4] ) );
  dp_1 \ANSWER/mem_reg[0][6][4]  ( .ip(n3428), .ck(clk), .q(
        \ANSWER/mem[0][6][4] ) );
  dp_1 \ANSWER/mem_reg[0][7][4]  ( .ip(n3427), .ck(clk), .q(
        \ANSWER/mem[0][7][4] ) );
  dp_1 \ANSWER/mem_reg[0][8][4]  ( .ip(n3426), .ck(clk), .q(
        \ANSWER/mem[0][8][4] ) );
  dp_1 \ANSWER/mem_reg[0][9][4]  ( .ip(n3425), .ck(clk), .q(
        \ANSWER/mem[0][9][4] ) );
  dp_1 \ANSWER/mem_reg[1][0][4]  ( .ip(n3424), .ck(clk), .q(
        \ANSWER/mem[1][0][4] ) );
  dp_1 \ANSWER/mem_reg[1][1][4]  ( .ip(n3423), .ck(clk), .q(
        \ANSWER/mem[1][1][4] ) );
  dp_1 \ANSWER/mem_reg[1][2][4]  ( .ip(n3422), .ck(clk), .q(
        \ANSWER/mem[1][2][4] ) );
  dp_1 \ANSWER/mem_reg[1][3][4]  ( .ip(n3421), .ck(clk), .q(
        \ANSWER/mem[1][3][4] ) );
  dp_1 \ANSWER/mem_reg[1][4][4]  ( .ip(n3420), .ck(clk), .q(
        \ANSWER/mem[1][4][4] ) );
  dp_1 \ANSWER/mem_reg[1][5][4]  ( .ip(n3419), .ck(clk), .q(
        \ANSWER/mem[1][5][4] ) );
  dp_1 \ANSWER/mem_reg[1][6][4]  ( .ip(n3418), .ck(clk), .q(
        \ANSWER/mem[1][6][4] ) );
  dp_1 \ANSWER/mem_reg[1][7][4]  ( .ip(n3417), .ck(clk), .q(
        \ANSWER/mem[1][7][4] ) );
  dp_1 \ANSWER/mem_reg[1][8][4]  ( .ip(n3416), .ck(clk), .q(
        \ANSWER/mem[1][8][4] ) );
  dp_1 \ANSWER/mem_reg[1][9][4]  ( .ip(n3415), .ck(clk), .q(
        \ANSWER/mem[1][9][4] ) );
  dp_1 \ANSWER/mem_reg[2][0][4]  ( .ip(n3414), .ck(clk), .q(
        \ANSWER/mem[2][0][4] ) );
  dp_1 \ANSWER/mem_reg[2][1][4]  ( .ip(n3413), .ck(clk), .q(
        \ANSWER/mem[2][1][4] ) );
  dp_1 \ANSWER/mem_reg[2][2][4]  ( .ip(n3412), .ck(clk), .q(
        \ANSWER/mem[2][2][4] ) );
  dp_1 \ANSWER/mem_reg[2][3][4]  ( .ip(n3411), .ck(clk), .q(
        \ANSWER/mem[2][3][4] ) );
  dp_1 \ANSWER/mem_reg[2][4][4]  ( .ip(n3410), .ck(clk), .q(
        \ANSWER/mem[2][4][4] ) );
  dp_1 \ANSWER/mem_reg[2][5][4]  ( .ip(n3409), .ck(clk), .q(
        \ANSWER/mem[2][5][4] ) );
  dp_1 \ANSWER/mem_reg[2][6][4]  ( .ip(n3408), .ck(clk), .q(
        \ANSWER/mem[2][6][4] ) );
  dp_1 \ANSWER/mem_reg[2][7][4]  ( .ip(n3407), .ck(clk), .q(
        \ANSWER/mem[2][7][4] ) );
  dp_1 \ANSWER/mem_reg[2][8][4]  ( .ip(n3406), .ck(clk), .q(
        \ANSWER/mem[2][8][4] ) );
  dp_1 \ANSWER/mem_reg[2][9][4]  ( .ip(n3405), .ck(clk), .q(
        \ANSWER/mem[2][9][4] ) );
  dp_1 \ANSWER/mem_reg[3][0][4]  ( .ip(n3404), .ck(clk), .q(
        \ANSWER/mem[3][0][4] ) );
  dp_1 \ANSWER/mem_reg[3][1][4]  ( .ip(n3403), .ck(clk), .q(
        \ANSWER/mem[3][1][4] ) );
  dp_1 \ANSWER/mem_reg[3][2][4]  ( .ip(n3402), .ck(clk), .q(
        \ANSWER/mem[3][2][4] ) );
  dp_1 \ANSWER/mem_reg[3][3][4]  ( .ip(n3401), .ck(clk), .q(
        \ANSWER/mem[3][3][4] ) );
  dp_1 \ANSWER/mem_reg[3][4][4]  ( .ip(n3400), .ck(clk), .q(
        \ANSWER/mem[3][4][4] ) );
  dp_1 \ANSWER/mem_reg[3][5][4]  ( .ip(n3399), .ck(clk), .q(
        \ANSWER/mem[3][5][4] ) );
  dp_1 \ANSWER/mem_reg[3][6][4]  ( .ip(n3398), .ck(clk), .q(
        \ANSWER/mem[3][6][4] ) );
  dp_1 \ANSWER/mem_reg[3][7][4]  ( .ip(n3397), .ck(clk), .q(
        \ANSWER/mem[3][7][4] ) );
  dp_1 \ANSWER/mem_reg[3][8][4]  ( .ip(n3396), .ck(clk), .q(
        \ANSWER/mem[3][8][4] ) );
  dp_1 \ANSWER/mem_reg[3][9][4]  ( .ip(n3395), .ck(clk), .q(
        \ANSWER/mem[3][9][4] ) );
  dp_1 \ANSWER/mem_reg[4][0][4]  ( .ip(n3394), .ck(clk), .q(
        \ANSWER/mem[4][0][4] ) );
  dp_1 \ANSWER/mem_reg[4][1][4]  ( .ip(n3393), .ck(clk), .q(
        \ANSWER/mem[4][1][4] ) );
  dp_1 \ANSWER/mem_reg[4][2][4]  ( .ip(n3392), .ck(clk), .q(
        \ANSWER/mem[4][2][4] ) );
  dp_1 \ANSWER/mem_reg[4][3][4]  ( .ip(n3391), .ck(clk), .q(
        \ANSWER/mem[4][3][4] ) );
  dp_1 \ANSWER/mem_reg[4][4][4]  ( .ip(n3390), .ck(clk), .q(
        \ANSWER/mem[4][4][4] ) );
  dp_1 \ANSWER/mem_reg[4][5][4]  ( .ip(n3389), .ck(clk), .q(
        \ANSWER/mem[4][5][4] ) );
  dp_1 \ANSWER/mem_reg[4][6][4]  ( .ip(n3388), .ck(clk), .q(
        \ANSWER/mem[4][6][4] ) );
  dp_1 \ANSWER/mem_reg[4][7][4]  ( .ip(n3387), .ck(clk), .q(
        \ANSWER/mem[4][7][4] ) );
  dp_1 \ANSWER/mem_reg[4][8][4]  ( .ip(n3386), .ck(clk), .q(
        \ANSWER/mem[4][8][4] ) );
  dp_1 \ANSWER/mem_reg[4][9][4]  ( .ip(n3385), .ck(clk), .q(
        \ANSWER/mem[4][9][4] ) );
  dp_1 \ANSWER/mem_reg[5][0][4]  ( .ip(n3384), .ck(clk), .q(
        \ANSWER/mem[5][0][4] ) );
  dp_1 \ANSWER/mem_reg[5][1][4]  ( .ip(n3383), .ck(clk), .q(
        \ANSWER/mem[5][1][4] ) );
  dp_1 \ANSWER/mem_reg[5][2][4]  ( .ip(n3382), .ck(clk), .q(
        \ANSWER/mem[5][2][4] ) );
  dp_1 \ANSWER/mem_reg[5][3][4]  ( .ip(n3381), .ck(clk), .q(
        \ANSWER/mem[5][3][4] ) );
  dp_1 \ANSWER/mem_reg[5][4][4]  ( .ip(n3380), .ck(clk), .q(
        \ANSWER/mem[5][4][4] ) );
  dp_1 \ANSWER/mem_reg[5][5][4]  ( .ip(n3379), .ck(clk), .q(
        \ANSWER/mem[5][5][4] ) );
  dp_1 \ANSWER/mem_reg[5][6][4]  ( .ip(n3378), .ck(clk), .q(
        \ANSWER/mem[5][6][4] ) );
  dp_1 \ANSWER/mem_reg[5][7][4]  ( .ip(n3377), .ck(clk), .q(
        \ANSWER/mem[5][7][4] ) );
  dp_1 \ANSWER/mem_reg[5][8][4]  ( .ip(n3376), .ck(clk), .q(
        \ANSWER/mem[5][8][4] ) );
  dp_1 \ANSWER/mem_reg[5][9][4]  ( .ip(n3375), .ck(clk), .q(
        \ANSWER/mem[5][9][4] ) );
  dp_1 \ANSWER/mem_reg[6][0][4]  ( .ip(n3374), .ck(clk), .q(
        \ANSWER/mem[6][0][4] ) );
  dp_1 \ANSWER/mem_reg[6][1][4]  ( .ip(n3373), .ck(clk), .q(
        \ANSWER/mem[6][1][4] ) );
  dp_1 \ANSWER/mem_reg[6][2][4]  ( .ip(n3372), .ck(clk), .q(
        \ANSWER/mem[6][2][4] ) );
  dp_1 \ANSWER/mem_reg[6][3][4]  ( .ip(n3371), .ck(clk), .q(
        \ANSWER/mem[6][3][4] ) );
  dp_1 \ANSWER/mem_reg[6][4][4]  ( .ip(n3370), .ck(clk), .q(
        \ANSWER/mem[6][4][4] ) );
  dp_1 \ANSWER/mem_reg[6][5][4]  ( .ip(n3369), .ck(clk), .q(
        \ANSWER/mem[6][5][4] ) );
  dp_1 \ANSWER/mem_reg[6][6][4]  ( .ip(n3368), .ck(clk), .q(
        \ANSWER/mem[6][6][4] ) );
  dp_1 \ANSWER/mem_reg[6][7][4]  ( .ip(n3367), .ck(clk), .q(
        \ANSWER/mem[6][7][4] ) );
  dp_1 \ANSWER/mem_reg[6][8][4]  ( .ip(n3366), .ck(clk), .q(
        \ANSWER/mem[6][8][4] ) );
  dp_1 \ANSWER/mem_reg[6][9][4]  ( .ip(n3365), .ck(clk), .q(
        \ANSWER/mem[6][9][4] ) );
  dp_1 \ANSWER/mem_reg[7][0][4]  ( .ip(n3364), .ck(clk), .q(
        \ANSWER/mem[7][0][4] ) );
  dp_1 \ANSWER/mem_reg[7][1][4]  ( .ip(n3363), .ck(clk), .q(
        \ANSWER/mem[7][1][4] ) );
  dp_1 \ANSWER/mem_reg[7][2][4]  ( .ip(n3362), .ck(clk), .q(
        \ANSWER/mem[7][2][4] ) );
  dp_1 \ANSWER/mem_reg[7][3][4]  ( .ip(n3361), .ck(clk), .q(
        \ANSWER/mem[7][3][4] ) );
  dp_1 \ANSWER/mem_reg[7][4][4]  ( .ip(n3360), .ck(clk), .q(
        \ANSWER/mem[7][4][4] ) );
  dp_1 \ANSWER/mem_reg[7][5][4]  ( .ip(n3359), .ck(clk), .q(
        \ANSWER/mem[7][5][4] ) );
  dp_1 \ANSWER/mem_reg[7][6][4]  ( .ip(n3358), .ck(clk), .q(
        \ANSWER/mem[7][6][4] ) );
  dp_1 \ANSWER/mem_reg[7][7][4]  ( .ip(n3357), .ck(clk), .q(
        \ANSWER/mem[7][7][4] ) );
  dp_1 \ANSWER/mem_reg[7][8][4]  ( .ip(n3356), .ck(clk), .q(
        \ANSWER/mem[7][8][4] ) );
  dp_1 \ANSWER/mem_reg[7][9][4]  ( .ip(n3355), .ck(clk), .q(
        \ANSWER/mem[7][9][4] ) );
  dp_1 \ANSWER/mem_reg[8][0][4]  ( .ip(n3354), .ck(clk), .q(
        \ANSWER/mem[8][0][4] ) );
  dp_1 \ANSWER/mem_reg[8][1][4]  ( .ip(n3353), .ck(clk), .q(
        \ANSWER/mem[8][1][4] ) );
  dp_1 \ANSWER/mem_reg[8][2][4]  ( .ip(n3352), .ck(clk), .q(
        \ANSWER/mem[8][2][4] ) );
  dp_1 \ANSWER/mem_reg[8][3][4]  ( .ip(n3351), .ck(clk), .q(
        \ANSWER/mem[8][3][4] ) );
  dp_1 \ANSWER/mem_reg[8][4][4]  ( .ip(n3350), .ck(clk), .q(
        \ANSWER/mem[8][4][4] ) );
  dp_1 \ANSWER/mem_reg[8][5][4]  ( .ip(n3349), .ck(clk), .q(
        \ANSWER/mem[8][5][4] ) );
  dp_1 \ANSWER/mem_reg[8][6][4]  ( .ip(n3348), .ck(clk), .q(
        \ANSWER/mem[8][6][4] ) );
  dp_1 \ANSWER/mem_reg[8][7][4]  ( .ip(n3347), .ck(clk), .q(
        \ANSWER/mem[8][7][4] ) );
  dp_1 \ANSWER/mem_reg[8][8][4]  ( .ip(n3346), .ck(clk), .q(
        \ANSWER/mem[8][8][4] ) );
  dp_1 \ANSWER/mem_reg[8][9][4]  ( .ip(n3345), .ck(clk), .q(
        \ANSWER/mem[8][9][4] ) );
  dp_1 \ANSWER/mem_reg[9][0][4]  ( .ip(n3344), .ck(clk), .q(
        \ANSWER/mem[9][0][4] ) );
  dp_1 \ANSWER/mem_reg[9][1][4]  ( .ip(n3343), .ck(clk), .q(
        \ANSWER/mem[9][1][4] ) );
  dp_1 \ANSWER/mem_reg[9][2][4]  ( .ip(n3342), .ck(clk), .q(
        \ANSWER/mem[9][2][4] ) );
  dp_1 \ANSWER/mem_reg[9][3][4]  ( .ip(n3341), .ck(clk), .q(
        \ANSWER/mem[9][3][4] ) );
  dp_1 \ANSWER/mem_reg[9][4][4]  ( .ip(n3340), .ck(clk), .q(
        \ANSWER/mem[9][4][4] ) );
  dp_1 \ANSWER/mem_reg[9][5][4]  ( .ip(n3339), .ck(clk), .q(
        \ANSWER/mem[9][5][4] ) );
  dp_1 \ANSWER/mem_reg[9][6][4]  ( .ip(n3338), .ck(clk), .q(
        \ANSWER/mem[9][6][4] ) );
  dp_1 \ANSWER/mem_reg[9][7][4]  ( .ip(n3337), .ck(clk), .q(
        \ANSWER/mem[9][7][4] ) );
  dp_1 \ANSWER/mem_reg[9][8][4]  ( .ip(n3336), .ck(clk), .q(
        \ANSWER/mem[9][8][4] ) );
  dp_1 \ANSWER/mem_reg[9][9][4]  ( .ip(n3335), .ck(clk), .q(
        \ANSWER/mem[9][9][4] ) );
  dp_1 \SIGMOID/lut_out_reg[5]  ( .ip(n3837), .ck(clk), .q(
        \SIGMOID/lut_out [5]) );
  dp_1 \ANSWER/mem_reg[0][0][5]  ( .ip(n3334), .ck(clk), .q(
        \ANSWER/mem[0][0][5] ) );
  dp_1 \ANSWER/mem_reg[0][1][5]  ( .ip(n3333), .ck(clk), .q(
        \ANSWER/mem[0][1][5] ) );
  dp_1 \ANSWER/mem_reg[0][2][5]  ( .ip(n3332), .ck(clk), .q(
        \ANSWER/mem[0][2][5] ) );
  dp_1 \ANSWER/mem_reg[0][3][5]  ( .ip(n3331), .ck(clk), .q(
        \ANSWER/mem[0][3][5] ) );
  dp_1 \ANSWER/mem_reg[0][4][5]  ( .ip(n3330), .ck(clk), .q(
        \ANSWER/mem[0][4][5] ) );
  dp_1 \ANSWER/mem_reg[0][5][5]  ( .ip(n3329), .ck(clk), .q(
        \ANSWER/mem[0][5][5] ) );
  dp_1 \ANSWER/mem_reg[0][6][5]  ( .ip(n3328), .ck(clk), .q(
        \ANSWER/mem[0][6][5] ) );
  dp_1 \ANSWER/mem_reg[0][7][5]  ( .ip(n3327), .ck(clk), .q(
        \ANSWER/mem[0][7][5] ) );
  dp_1 \ANSWER/mem_reg[0][8][5]  ( .ip(n3326), .ck(clk), .q(
        \ANSWER/mem[0][8][5] ) );
  dp_1 \ANSWER/mem_reg[0][9][5]  ( .ip(n3325), .ck(clk), .q(
        \ANSWER/mem[0][9][5] ) );
  dp_1 \ANSWER/mem_reg[1][0][5]  ( .ip(n3324), .ck(clk), .q(
        \ANSWER/mem[1][0][5] ) );
  dp_1 \ANSWER/mem_reg[1][1][5]  ( .ip(n3323), .ck(clk), .q(
        \ANSWER/mem[1][1][5] ) );
  dp_1 \ANSWER/mem_reg[1][2][5]  ( .ip(n3322), .ck(clk), .q(
        \ANSWER/mem[1][2][5] ) );
  dp_1 \ANSWER/mem_reg[1][3][5]  ( .ip(n3321), .ck(clk), .q(
        \ANSWER/mem[1][3][5] ) );
  dp_1 \ANSWER/mem_reg[1][4][5]  ( .ip(n3320), .ck(clk), .q(
        \ANSWER/mem[1][4][5] ) );
  dp_1 \ANSWER/mem_reg[1][5][5]  ( .ip(n3319), .ck(clk), .q(
        \ANSWER/mem[1][5][5] ) );
  dp_1 \ANSWER/mem_reg[1][6][5]  ( .ip(n3318), .ck(clk), .q(
        \ANSWER/mem[1][6][5] ) );
  dp_1 \ANSWER/mem_reg[1][7][5]  ( .ip(n3317), .ck(clk), .q(
        \ANSWER/mem[1][7][5] ) );
  dp_1 \ANSWER/mem_reg[1][8][5]  ( .ip(n3316), .ck(clk), .q(
        \ANSWER/mem[1][8][5] ) );
  dp_1 \ANSWER/mem_reg[1][9][5]  ( .ip(n3315), .ck(clk), .q(
        \ANSWER/mem[1][9][5] ) );
  dp_1 \ANSWER/mem_reg[2][0][5]  ( .ip(n3314), .ck(clk), .q(
        \ANSWER/mem[2][0][5] ) );
  dp_1 \ANSWER/mem_reg[2][1][5]  ( .ip(n3313), .ck(clk), .q(
        \ANSWER/mem[2][1][5] ) );
  dp_1 \ANSWER/mem_reg[2][2][5]  ( .ip(n3312), .ck(clk), .q(
        \ANSWER/mem[2][2][5] ) );
  dp_1 \ANSWER/mem_reg[2][3][5]  ( .ip(n3311), .ck(clk), .q(
        \ANSWER/mem[2][3][5] ) );
  dp_1 \ANSWER/mem_reg[2][4][5]  ( .ip(n3310), .ck(clk), .q(
        \ANSWER/mem[2][4][5] ) );
  dp_1 \ANSWER/mem_reg[2][5][5]  ( .ip(n3309), .ck(clk), .q(
        \ANSWER/mem[2][5][5] ) );
  dp_1 \ANSWER/mem_reg[2][6][5]  ( .ip(n3308), .ck(clk), .q(
        \ANSWER/mem[2][6][5] ) );
  dp_1 \ANSWER/mem_reg[2][7][5]  ( .ip(n3307), .ck(clk), .q(
        \ANSWER/mem[2][7][5] ) );
  dp_1 \ANSWER/mem_reg[2][8][5]  ( .ip(n3306), .ck(clk), .q(
        \ANSWER/mem[2][8][5] ) );
  dp_1 \ANSWER/mem_reg[2][9][5]  ( .ip(n3305), .ck(clk), .q(
        \ANSWER/mem[2][9][5] ) );
  dp_1 \ANSWER/mem_reg[3][0][5]  ( .ip(n3304), .ck(clk), .q(
        \ANSWER/mem[3][0][5] ) );
  dp_1 \ANSWER/mem_reg[3][1][5]  ( .ip(n3303), .ck(clk), .q(
        \ANSWER/mem[3][1][5] ) );
  dp_1 \ANSWER/mem_reg[3][2][5]  ( .ip(n3302), .ck(clk), .q(
        \ANSWER/mem[3][2][5] ) );
  dp_1 \ANSWER/mem_reg[3][3][5]  ( .ip(n3301), .ck(clk), .q(
        \ANSWER/mem[3][3][5] ) );
  dp_1 \ANSWER/mem_reg[3][4][5]  ( .ip(n3300), .ck(clk), .q(
        \ANSWER/mem[3][4][5] ) );
  dp_1 \ANSWER/mem_reg[3][5][5]  ( .ip(n3299), .ck(clk), .q(
        \ANSWER/mem[3][5][5] ) );
  dp_1 \ANSWER/mem_reg[3][6][5]  ( .ip(n3298), .ck(clk), .q(
        \ANSWER/mem[3][6][5] ) );
  dp_1 \ANSWER/mem_reg[3][7][5]  ( .ip(n3297), .ck(clk), .q(
        \ANSWER/mem[3][7][5] ) );
  dp_1 \ANSWER/mem_reg[3][8][5]  ( .ip(n3296), .ck(clk), .q(
        \ANSWER/mem[3][8][5] ) );
  dp_1 \ANSWER/mem_reg[3][9][5]  ( .ip(n3295), .ck(clk), .q(
        \ANSWER/mem[3][9][5] ) );
  dp_1 \ANSWER/mem_reg[4][0][5]  ( .ip(n3294), .ck(clk), .q(
        \ANSWER/mem[4][0][5] ) );
  dp_1 \ANSWER/mem_reg[4][1][5]  ( .ip(n3293), .ck(clk), .q(
        \ANSWER/mem[4][1][5] ) );
  dp_1 \ANSWER/mem_reg[4][2][5]  ( .ip(n3292), .ck(clk), .q(
        \ANSWER/mem[4][2][5] ) );
  dp_1 \ANSWER/mem_reg[4][3][5]  ( .ip(n3291), .ck(clk), .q(
        \ANSWER/mem[4][3][5] ) );
  dp_1 \ANSWER/mem_reg[4][4][5]  ( .ip(n3290), .ck(clk), .q(
        \ANSWER/mem[4][4][5] ) );
  dp_1 \ANSWER/mem_reg[4][5][5]  ( .ip(n3289), .ck(clk), .q(
        \ANSWER/mem[4][5][5] ) );
  dp_1 \ANSWER/mem_reg[4][6][5]  ( .ip(n3288), .ck(clk), .q(
        \ANSWER/mem[4][6][5] ) );
  dp_1 \ANSWER/mem_reg[4][7][5]  ( .ip(n3287), .ck(clk), .q(
        \ANSWER/mem[4][7][5] ) );
  dp_1 \ANSWER/mem_reg[4][8][5]  ( .ip(n3286), .ck(clk), .q(
        \ANSWER/mem[4][8][5] ) );
  dp_1 \ANSWER/mem_reg[4][9][5]  ( .ip(n3285), .ck(clk), .q(
        \ANSWER/mem[4][9][5] ) );
  dp_1 \ANSWER/mem_reg[5][0][5]  ( .ip(n3284), .ck(clk), .q(
        \ANSWER/mem[5][0][5] ) );
  dp_1 \ANSWER/mem_reg[5][1][5]  ( .ip(n3283), .ck(clk), .q(
        \ANSWER/mem[5][1][5] ) );
  dp_1 \ANSWER/mem_reg[5][2][5]  ( .ip(n3282), .ck(clk), .q(
        \ANSWER/mem[5][2][5] ) );
  dp_1 \ANSWER/mem_reg[5][3][5]  ( .ip(n3281), .ck(clk), .q(
        \ANSWER/mem[5][3][5] ) );
  dp_1 \ANSWER/mem_reg[5][4][5]  ( .ip(n3280), .ck(clk), .q(
        \ANSWER/mem[5][4][5] ) );
  dp_1 \ANSWER/mem_reg[5][5][5]  ( .ip(n3279), .ck(clk), .q(
        \ANSWER/mem[5][5][5] ) );
  dp_1 \ANSWER/mem_reg[5][6][5]  ( .ip(n3278), .ck(clk), .q(
        \ANSWER/mem[5][6][5] ) );
  dp_1 \ANSWER/mem_reg[5][7][5]  ( .ip(n3277), .ck(clk), .q(
        \ANSWER/mem[5][7][5] ) );
  dp_1 \ANSWER/mem_reg[5][8][5]  ( .ip(n3276), .ck(clk), .q(
        \ANSWER/mem[5][8][5] ) );
  dp_1 \ANSWER/mem_reg[5][9][5]  ( .ip(n3275), .ck(clk), .q(
        \ANSWER/mem[5][9][5] ) );
  dp_1 \ANSWER/mem_reg[6][0][5]  ( .ip(n3274), .ck(clk), .q(
        \ANSWER/mem[6][0][5] ) );
  dp_1 \ANSWER/mem_reg[6][1][5]  ( .ip(n3273), .ck(clk), .q(
        \ANSWER/mem[6][1][5] ) );
  dp_1 \ANSWER/mem_reg[6][2][5]  ( .ip(n3272), .ck(clk), .q(
        \ANSWER/mem[6][2][5] ) );
  dp_1 \ANSWER/mem_reg[6][3][5]  ( .ip(n3271), .ck(clk), .q(
        \ANSWER/mem[6][3][5] ) );
  dp_1 \ANSWER/mem_reg[6][4][5]  ( .ip(n3270), .ck(clk), .q(
        \ANSWER/mem[6][4][5] ) );
  dp_1 \ANSWER/mem_reg[6][5][5]  ( .ip(n3269), .ck(clk), .q(
        \ANSWER/mem[6][5][5] ) );
  dp_1 \ANSWER/mem_reg[6][6][5]  ( .ip(n3268), .ck(clk), .q(
        \ANSWER/mem[6][6][5] ) );
  dp_1 \ANSWER/mem_reg[6][7][5]  ( .ip(n3267), .ck(clk), .q(
        \ANSWER/mem[6][7][5] ) );
  dp_1 \ANSWER/mem_reg[6][8][5]  ( .ip(n3266), .ck(clk), .q(
        \ANSWER/mem[6][8][5] ) );
  dp_1 \ANSWER/mem_reg[6][9][5]  ( .ip(n3265), .ck(clk), .q(
        \ANSWER/mem[6][9][5] ) );
  dp_1 \ANSWER/mem_reg[7][0][5]  ( .ip(n3264), .ck(clk), .q(
        \ANSWER/mem[7][0][5] ) );
  dp_1 \ANSWER/mem_reg[7][1][5]  ( .ip(n3263), .ck(clk), .q(
        \ANSWER/mem[7][1][5] ) );
  dp_1 \ANSWER/mem_reg[7][2][5]  ( .ip(n3262), .ck(clk), .q(
        \ANSWER/mem[7][2][5] ) );
  dp_1 \ANSWER/mem_reg[7][3][5]  ( .ip(n3261), .ck(clk), .q(
        \ANSWER/mem[7][3][5] ) );
  dp_1 \ANSWER/mem_reg[7][4][5]  ( .ip(n3260), .ck(clk), .q(
        \ANSWER/mem[7][4][5] ) );
  dp_1 \ANSWER/mem_reg[7][5][5]  ( .ip(n3259), .ck(clk), .q(
        \ANSWER/mem[7][5][5] ) );
  dp_1 \ANSWER/mem_reg[7][6][5]  ( .ip(n3258), .ck(clk), .q(
        \ANSWER/mem[7][6][5] ) );
  dp_1 \ANSWER/mem_reg[7][7][5]  ( .ip(n3257), .ck(clk), .q(
        \ANSWER/mem[7][7][5] ) );
  dp_1 \ANSWER/mem_reg[7][8][5]  ( .ip(n3256), .ck(clk), .q(
        \ANSWER/mem[7][8][5] ) );
  dp_1 \ANSWER/mem_reg[7][9][5]  ( .ip(n3255), .ck(clk), .q(
        \ANSWER/mem[7][9][5] ) );
  dp_1 \ANSWER/mem_reg[8][0][5]  ( .ip(n3254), .ck(clk), .q(
        \ANSWER/mem[8][0][5] ) );
  dp_1 \ANSWER/mem_reg[8][1][5]  ( .ip(n3253), .ck(clk), .q(
        \ANSWER/mem[8][1][5] ) );
  dp_1 \ANSWER/mem_reg[8][2][5]  ( .ip(n3252), .ck(clk), .q(
        \ANSWER/mem[8][2][5] ) );
  dp_1 \ANSWER/mem_reg[8][3][5]  ( .ip(n3251), .ck(clk), .q(
        \ANSWER/mem[8][3][5] ) );
  dp_1 \ANSWER/mem_reg[8][4][5]  ( .ip(n3250), .ck(clk), .q(
        \ANSWER/mem[8][4][5] ) );
  dp_1 \ANSWER/mem_reg[8][5][5]  ( .ip(n3249), .ck(clk), .q(
        \ANSWER/mem[8][5][5] ) );
  dp_1 \ANSWER/mem_reg[8][6][5]  ( .ip(n3248), .ck(clk), .q(
        \ANSWER/mem[8][6][5] ) );
  dp_1 \ANSWER/mem_reg[8][7][5]  ( .ip(n3247), .ck(clk), .q(
        \ANSWER/mem[8][7][5] ) );
  dp_1 \ANSWER/mem_reg[8][8][5]  ( .ip(n3246), .ck(clk), .q(
        \ANSWER/mem[8][8][5] ) );
  dp_1 \ANSWER/mem_reg[8][9][5]  ( .ip(n3245), .ck(clk), .q(
        \ANSWER/mem[8][9][5] ) );
  dp_1 \ANSWER/mem_reg[9][0][5]  ( .ip(n3244), .ck(clk), .q(
        \ANSWER/mem[9][0][5] ) );
  dp_1 \ANSWER/mem_reg[9][1][5]  ( .ip(n3243), .ck(clk), .q(
        \ANSWER/mem[9][1][5] ) );
  dp_1 \ANSWER/mem_reg[9][2][5]  ( .ip(n3242), .ck(clk), .q(
        \ANSWER/mem[9][2][5] ) );
  dp_1 \ANSWER/mem_reg[9][3][5]  ( .ip(n3241), .ck(clk), .q(
        \ANSWER/mem[9][3][5] ) );
  dp_1 \ANSWER/mem_reg[9][4][5]  ( .ip(n3240), .ck(clk), .q(
        \ANSWER/mem[9][4][5] ) );
  dp_1 \ANSWER/mem_reg[9][5][5]  ( .ip(n3239), .ck(clk), .q(
        \ANSWER/mem[9][5][5] ) );
  dp_1 \ANSWER/mem_reg[9][6][5]  ( .ip(n3238), .ck(clk), .q(
        \ANSWER/mem[9][6][5] ) );
  dp_1 \ANSWER/mem_reg[9][7][5]  ( .ip(n3237), .ck(clk), .q(
        \ANSWER/mem[9][7][5] ) );
  dp_1 \ANSWER/mem_reg[9][8][5]  ( .ip(n3236), .ck(clk), .q(
        \ANSWER/mem[9][8][5] ) );
  dp_1 \ANSWER/mem_reg[9][9][5]  ( .ip(n3235), .ck(clk), .q(
        \ANSWER/mem[9][9][5] ) );
  dp_1 \SIGMOID/lut_out_reg[6]  ( .ip(n3836), .ck(clk), .q(
        \SIGMOID/lut_out [6]) );
  dp_1 \ANSWER/mem_reg[0][0][6]  ( .ip(n3234), .ck(clk), .q(
        \ANSWER/mem[0][0][6] ) );
  dp_1 \ANSWER/mem_reg[0][1][6]  ( .ip(n3233), .ck(clk), .q(
        \ANSWER/mem[0][1][6] ) );
  dp_1 \ANSWER/mem_reg[0][2][6]  ( .ip(n3232), .ck(clk), .q(
        \ANSWER/mem[0][2][6] ) );
  dp_1 \ANSWER/mem_reg[0][3][6]  ( .ip(n3231), .ck(clk), .q(
        \ANSWER/mem[0][3][6] ) );
  dp_1 \ANSWER/mem_reg[0][4][6]  ( .ip(n3230), .ck(clk), .q(
        \ANSWER/mem[0][4][6] ) );
  dp_1 \ANSWER/mem_reg[0][5][6]  ( .ip(n3229), .ck(clk), .q(
        \ANSWER/mem[0][5][6] ) );
  dp_1 \ANSWER/mem_reg[0][6][6]  ( .ip(n3228), .ck(clk), .q(
        \ANSWER/mem[0][6][6] ) );
  dp_1 \ANSWER/mem_reg[0][7][6]  ( .ip(n3227), .ck(clk), .q(
        \ANSWER/mem[0][7][6] ) );
  dp_1 \ANSWER/mem_reg[0][8][6]  ( .ip(n3226), .ck(clk), .q(
        \ANSWER/mem[0][8][6] ) );
  dp_1 \ANSWER/mem_reg[0][9][6]  ( .ip(n3225), .ck(clk), .q(
        \ANSWER/mem[0][9][6] ) );
  dp_1 \ANSWER/mem_reg[1][0][6]  ( .ip(n3224), .ck(clk), .q(
        \ANSWER/mem[1][0][6] ) );
  dp_1 \ANSWER/mem_reg[1][1][6]  ( .ip(n3223), .ck(clk), .q(
        \ANSWER/mem[1][1][6] ) );
  dp_1 \ANSWER/mem_reg[1][2][6]  ( .ip(n3222), .ck(clk), .q(
        \ANSWER/mem[1][2][6] ) );
  dp_1 \ANSWER/mem_reg[1][3][6]  ( .ip(n3221), .ck(clk), .q(
        \ANSWER/mem[1][3][6] ) );
  dp_1 \ANSWER/mem_reg[1][4][6]  ( .ip(n3220), .ck(clk), .q(
        \ANSWER/mem[1][4][6] ) );
  dp_1 \ANSWER/mem_reg[1][5][6]  ( .ip(n3219), .ck(clk), .q(
        \ANSWER/mem[1][5][6] ) );
  dp_1 \ANSWER/mem_reg[1][6][6]  ( .ip(n3218), .ck(clk), .q(
        \ANSWER/mem[1][6][6] ) );
  dp_1 \ANSWER/mem_reg[1][7][6]  ( .ip(n3217), .ck(clk), .q(
        \ANSWER/mem[1][7][6] ) );
  dp_1 \ANSWER/mem_reg[1][8][6]  ( .ip(n3216), .ck(clk), .q(
        \ANSWER/mem[1][8][6] ) );
  dp_1 \ANSWER/mem_reg[1][9][6]  ( .ip(n3215), .ck(clk), .q(
        \ANSWER/mem[1][9][6] ) );
  dp_1 \ANSWER/mem_reg[2][0][6]  ( .ip(n3214), .ck(clk), .q(
        \ANSWER/mem[2][0][6] ) );
  dp_1 \ANSWER/mem_reg[2][1][6]  ( .ip(n3213), .ck(clk), .q(
        \ANSWER/mem[2][1][6] ) );
  dp_1 \ANSWER/mem_reg[2][2][6]  ( .ip(n3212), .ck(clk), .q(
        \ANSWER/mem[2][2][6] ) );
  dp_1 \ANSWER/mem_reg[2][3][6]  ( .ip(n3211), .ck(clk), .q(
        \ANSWER/mem[2][3][6] ) );
  dp_1 \ANSWER/mem_reg[2][4][6]  ( .ip(n3210), .ck(clk), .q(
        \ANSWER/mem[2][4][6] ) );
  dp_1 \ANSWER/mem_reg[2][5][6]  ( .ip(n3209), .ck(clk), .q(
        \ANSWER/mem[2][5][6] ) );
  dp_1 \ANSWER/mem_reg[2][6][6]  ( .ip(n3208), .ck(clk), .q(
        \ANSWER/mem[2][6][6] ) );
  dp_1 \ANSWER/mem_reg[2][7][6]  ( .ip(n3207), .ck(clk), .q(
        \ANSWER/mem[2][7][6] ) );
  dp_1 \ANSWER/mem_reg[2][8][6]  ( .ip(n3206), .ck(clk), .q(
        \ANSWER/mem[2][8][6] ) );
  dp_1 \ANSWER/mem_reg[2][9][6]  ( .ip(n3205), .ck(clk), .q(
        \ANSWER/mem[2][9][6] ) );
  dp_1 \ANSWER/mem_reg[3][0][6]  ( .ip(n3204), .ck(clk), .q(
        \ANSWER/mem[3][0][6] ) );
  dp_1 \ANSWER/mem_reg[3][1][6]  ( .ip(n3203), .ck(clk), .q(
        \ANSWER/mem[3][1][6] ) );
  dp_1 \ANSWER/mem_reg[3][2][6]  ( .ip(n3202), .ck(clk), .q(
        \ANSWER/mem[3][2][6] ) );
  dp_1 \ANSWER/mem_reg[3][3][6]  ( .ip(n3201), .ck(clk), .q(
        \ANSWER/mem[3][3][6] ) );
  dp_1 \ANSWER/mem_reg[3][4][6]  ( .ip(n3200), .ck(clk), .q(
        \ANSWER/mem[3][4][6] ) );
  dp_1 \ANSWER/mem_reg[3][5][6]  ( .ip(n3199), .ck(clk), .q(
        \ANSWER/mem[3][5][6] ) );
  dp_1 \ANSWER/mem_reg[3][6][6]  ( .ip(n3198), .ck(clk), .q(
        \ANSWER/mem[3][6][6] ) );
  dp_1 \ANSWER/mem_reg[3][7][6]  ( .ip(n3197), .ck(clk), .q(
        \ANSWER/mem[3][7][6] ) );
  dp_1 \ANSWER/mem_reg[3][8][6]  ( .ip(n3196), .ck(clk), .q(
        \ANSWER/mem[3][8][6] ) );
  dp_1 \ANSWER/mem_reg[3][9][6]  ( .ip(n3195), .ck(clk), .q(
        \ANSWER/mem[3][9][6] ) );
  dp_1 \ANSWER/mem_reg[4][0][6]  ( .ip(n3194), .ck(clk), .q(
        \ANSWER/mem[4][0][6] ) );
  dp_1 \ANSWER/mem_reg[4][1][6]  ( .ip(n3193), .ck(clk), .q(
        \ANSWER/mem[4][1][6] ) );
  dp_1 \ANSWER/mem_reg[4][2][6]  ( .ip(n3192), .ck(clk), .q(
        \ANSWER/mem[4][2][6] ) );
  dp_1 \ANSWER/mem_reg[4][3][6]  ( .ip(n3191), .ck(clk), .q(
        \ANSWER/mem[4][3][6] ) );
  dp_1 \ANSWER/mem_reg[4][4][6]  ( .ip(n3190), .ck(clk), .q(
        \ANSWER/mem[4][4][6] ) );
  dp_1 \ANSWER/mem_reg[4][5][6]  ( .ip(n3189), .ck(clk), .q(
        \ANSWER/mem[4][5][6] ) );
  dp_1 \ANSWER/mem_reg[4][6][6]  ( .ip(n3188), .ck(clk), .q(
        \ANSWER/mem[4][6][6] ) );
  dp_1 \ANSWER/mem_reg[4][7][6]  ( .ip(n3187), .ck(clk), .q(
        \ANSWER/mem[4][7][6] ) );
  dp_1 \ANSWER/mem_reg[4][8][6]  ( .ip(n3186), .ck(clk), .q(
        \ANSWER/mem[4][8][6] ) );
  dp_1 \ANSWER/mem_reg[4][9][6]  ( .ip(n3185), .ck(clk), .q(
        \ANSWER/mem[4][9][6] ) );
  dp_1 \ANSWER/mem_reg[5][0][6]  ( .ip(n3184), .ck(clk), .q(
        \ANSWER/mem[5][0][6] ) );
  dp_1 \ANSWER/mem_reg[5][1][6]  ( .ip(n3183), .ck(clk), .q(
        \ANSWER/mem[5][1][6] ) );
  dp_1 \ANSWER/mem_reg[5][2][6]  ( .ip(n3182), .ck(clk), .q(
        \ANSWER/mem[5][2][6] ) );
  dp_1 \ANSWER/mem_reg[5][3][6]  ( .ip(n3181), .ck(clk), .q(
        \ANSWER/mem[5][3][6] ) );
  dp_1 \ANSWER/mem_reg[5][4][6]  ( .ip(n3180), .ck(clk), .q(
        \ANSWER/mem[5][4][6] ) );
  dp_1 \ANSWER/mem_reg[5][5][6]  ( .ip(n3179), .ck(clk), .q(
        \ANSWER/mem[5][5][6] ) );
  dp_1 \ANSWER/mem_reg[5][6][6]  ( .ip(n3178), .ck(clk), .q(
        \ANSWER/mem[5][6][6] ) );
  dp_1 \ANSWER/mem_reg[5][7][6]  ( .ip(n3177), .ck(clk), .q(
        \ANSWER/mem[5][7][6] ) );
  dp_1 \ANSWER/mem_reg[5][8][6]  ( .ip(n3176), .ck(clk), .q(
        \ANSWER/mem[5][8][6] ) );
  dp_1 \ANSWER/mem_reg[5][9][6]  ( .ip(n3175), .ck(clk), .q(
        \ANSWER/mem[5][9][6] ) );
  dp_1 \ANSWER/mem_reg[6][0][6]  ( .ip(n3174), .ck(clk), .q(
        \ANSWER/mem[6][0][6] ) );
  dp_1 \ANSWER/mem_reg[6][1][6]  ( .ip(n3173), .ck(clk), .q(
        \ANSWER/mem[6][1][6] ) );
  dp_1 \ANSWER/mem_reg[6][2][6]  ( .ip(n3172), .ck(clk), .q(
        \ANSWER/mem[6][2][6] ) );
  dp_1 \ANSWER/mem_reg[6][3][6]  ( .ip(n3171), .ck(clk), .q(
        \ANSWER/mem[6][3][6] ) );
  dp_1 \ANSWER/mem_reg[6][4][6]  ( .ip(n3170), .ck(clk), .q(
        \ANSWER/mem[6][4][6] ) );
  dp_1 \ANSWER/mem_reg[6][5][6]  ( .ip(n3169), .ck(clk), .q(
        \ANSWER/mem[6][5][6] ) );
  dp_1 \ANSWER/mem_reg[6][6][6]  ( .ip(n3168), .ck(clk), .q(
        \ANSWER/mem[6][6][6] ) );
  dp_1 \ANSWER/mem_reg[6][7][6]  ( .ip(n3167), .ck(clk), .q(
        \ANSWER/mem[6][7][6] ) );
  dp_1 \ANSWER/mem_reg[6][8][6]  ( .ip(n3166), .ck(clk), .q(
        \ANSWER/mem[6][8][6] ) );
  dp_1 \ANSWER/mem_reg[6][9][6]  ( .ip(n3165), .ck(clk), .q(
        \ANSWER/mem[6][9][6] ) );
  dp_1 \ANSWER/mem_reg[7][0][6]  ( .ip(n3164), .ck(clk), .q(
        \ANSWER/mem[7][0][6] ) );
  dp_1 \ANSWER/mem_reg[7][1][6]  ( .ip(n3163), .ck(clk), .q(
        \ANSWER/mem[7][1][6] ) );
  dp_1 \ANSWER/mem_reg[7][2][6]  ( .ip(n3162), .ck(clk), .q(
        \ANSWER/mem[7][2][6] ) );
  dp_1 \ANSWER/mem_reg[7][3][6]  ( .ip(n3161), .ck(clk), .q(
        \ANSWER/mem[7][3][6] ) );
  dp_1 \ANSWER/mem_reg[7][4][6]  ( .ip(n3160), .ck(clk), .q(
        \ANSWER/mem[7][4][6] ) );
  dp_1 \ANSWER/mem_reg[7][5][6]  ( .ip(n3159), .ck(clk), .q(
        \ANSWER/mem[7][5][6] ) );
  dp_1 \ANSWER/mem_reg[7][6][6]  ( .ip(n3158), .ck(clk), .q(
        \ANSWER/mem[7][6][6] ) );
  dp_1 \ANSWER/mem_reg[7][7][6]  ( .ip(n3157), .ck(clk), .q(
        \ANSWER/mem[7][7][6] ) );
  dp_1 \ANSWER/mem_reg[7][8][6]  ( .ip(n3156), .ck(clk), .q(
        \ANSWER/mem[7][8][6] ) );
  dp_1 \ANSWER/mem_reg[7][9][6]  ( .ip(n3155), .ck(clk), .q(
        \ANSWER/mem[7][9][6] ) );
  dp_1 \ANSWER/mem_reg[8][0][6]  ( .ip(n3154), .ck(clk), .q(
        \ANSWER/mem[8][0][6] ) );
  dp_1 \ANSWER/mem_reg[8][1][6]  ( .ip(n3153), .ck(clk), .q(
        \ANSWER/mem[8][1][6] ) );
  dp_1 \ANSWER/mem_reg[8][2][6]  ( .ip(n3152), .ck(clk), .q(
        \ANSWER/mem[8][2][6] ) );
  dp_1 \ANSWER/mem_reg[8][3][6]  ( .ip(n3151), .ck(clk), .q(
        \ANSWER/mem[8][3][6] ) );
  dp_1 \ANSWER/mem_reg[8][4][6]  ( .ip(n3150), .ck(clk), .q(
        \ANSWER/mem[8][4][6] ) );
  dp_1 \ANSWER/mem_reg[8][5][6]  ( .ip(n3149), .ck(clk), .q(
        \ANSWER/mem[8][5][6] ) );
  dp_1 \ANSWER/mem_reg[8][6][6]  ( .ip(n3148), .ck(clk), .q(
        \ANSWER/mem[8][6][6] ) );
  dp_1 \ANSWER/mem_reg[8][7][6]  ( .ip(n3147), .ck(clk), .q(
        \ANSWER/mem[8][7][6] ) );
  dp_1 \ANSWER/mem_reg[8][8][6]  ( .ip(n3146), .ck(clk), .q(
        \ANSWER/mem[8][8][6] ) );
  dp_1 \ANSWER/mem_reg[8][9][6]  ( .ip(n3145), .ck(clk), .q(
        \ANSWER/mem[8][9][6] ) );
  dp_1 \ANSWER/mem_reg[9][0][6]  ( .ip(n3144), .ck(clk), .q(
        \ANSWER/mem[9][0][6] ) );
  dp_1 \ANSWER/mem_reg[9][1][6]  ( .ip(n3143), .ck(clk), .q(
        \ANSWER/mem[9][1][6] ) );
  dp_1 \ANSWER/mem_reg[9][2][6]  ( .ip(n3142), .ck(clk), .q(
        \ANSWER/mem[9][2][6] ) );
  dp_1 \ANSWER/mem_reg[9][3][6]  ( .ip(n3141), .ck(clk), .q(
        \ANSWER/mem[9][3][6] ) );
  dp_1 \ANSWER/mem_reg[9][4][6]  ( .ip(n3140), .ck(clk), .q(
        \ANSWER/mem[9][4][6] ) );
  dp_1 \ANSWER/mem_reg[9][5][6]  ( .ip(n3139), .ck(clk), .q(
        \ANSWER/mem[9][5][6] ) );
  dp_1 \ANSWER/mem_reg[9][6][6]  ( .ip(n3138), .ck(clk), .q(
        \ANSWER/mem[9][6][6] ) );
  dp_1 \ANSWER/mem_reg[9][7][6]  ( .ip(n3137), .ck(clk), .q(
        \ANSWER/mem[9][7][6] ) );
  dp_1 \ANSWER/mem_reg[9][8][6]  ( .ip(n3136), .ck(clk), .q(
        \ANSWER/mem[9][8][6] ) );
  dp_1 \ANSWER/mem_reg[9][9][6]  ( .ip(n3135), .ck(clk), .q(
        \ANSWER/mem[9][9][6] ) );
  dp_1 \SIGMOID/lut_out_reg[7]  ( .ip(n3835), .ck(clk), .q(
        \SIGMOID/lut_out [7]) );
  dp_1 \ANSWER/mem_reg[0][0][7]  ( .ip(n3134), .ck(clk), .q(
        \ANSWER/mem[0][0][7] ) );
  dp_1 \ANSWER/mem_reg[0][1][7]  ( .ip(n3133), .ck(clk), .q(
        \ANSWER/mem[0][1][7] ) );
  dp_1 \ANSWER/mem_reg[0][2][7]  ( .ip(n3132), .ck(clk), .q(
        \ANSWER/mem[0][2][7] ) );
  dp_1 \ANSWER/mem_reg[0][3][7]  ( .ip(n3131), .ck(clk), .q(
        \ANSWER/mem[0][3][7] ) );
  dp_1 \ANSWER/mem_reg[0][4][7]  ( .ip(n3130), .ck(clk), .q(
        \ANSWER/mem[0][4][7] ) );
  dp_1 \ANSWER/mem_reg[0][5][7]  ( .ip(n3129), .ck(clk), .q(
        \ANSWER/mem[0][5][7] ) );
  dp_1 \ANSWER/mem_reg[0][6][7]  ( .ip(n3128), .ck(clk), .q(
        \ANSWER/mem[0][6][7] ) );
  dp_1 \ANSWER/mem_reg[0][7][7]  ( .ip(n3127), .ck(clk), .q(
        \ANSWER/mem[0][7][7] ) );
  dp_1 \ANSWER/mem_reg[0][8][7]  ( .ip(n3126), .ck(clk), .q(
        \ANSWER/mem[0][8][7] ) );
  dp_1 \ANSWER/mem_reg[0][9][7]  ( .ip(n3125), .ck(clk), .q(
        \ANSWER/mem[0][9][7] ) );
  dp_1 \ANSWER/mem_reg[1][0][7]  ( .ip(n3124), .ck(clk), .q(
        \ANSWER/mem[1][0][7] ) );
  dp_1 \ANSWER/mem_reg[1][1][7]  ( .ip(n3123), .ck(clk), .q(
        \ANSWER/mem[1][1][7] ) );
  dp_1 \ANSWER/mem_reg[1][2][7]  ( .ip(n3122), .ck(clk), .q(
        \ANSWER/mem[1][2][7] ) );
  dp_1 \ANSWER/mem_reg[1][3][7]  ( .ip(n3121), .ck(clk), .q(
        \ANSWER/mem[1][3][7] ) );
  dp_1 \ANSWER/mem_reg[1][4][7]  ( .ip(n3120), .ck(clk), .q(
        \ANSWER/mem[1][4][7] ) );
  dp_1 \ANSWER/mem_reg[1][5][7]  ( .ip(n3119), .ck(clk), .q(
        \ANSWER/mem[1][5][7] ) );
  dp_1 \ANSWER/mem_reg[1][6][7]  ( .ip(n3118), .ck(clk), .q(
        \ANSWER/mem[1][6][7] ) );
  dp_1 \ANSWER/mem_reg[1][7][7]  ( .ip(n3117), .ck(clk), .q(
        \ANSWER/mem[1][7][7] ) );
  dp_1 \ANSWER/mem_reg[1][8][7]  ( .ip(n3116), .ck(clk), .q(
        \ANSWER/mem[1][8][7] ) );
  dp_1 \ANSWER/mem_reg[1][9][7]  ( .ip(n3115), .ck(clk), .q(
        \ANSWER/mem[1][9][7] ) );
  dp_1 \ANSWER/mem_reg[2][0][7]  ( .ip(n3114), .ck(clk), .q(
        \ANSWER/mem[2][0][7] ) );
  dp_1 \ANSWER/mem_reg[2][1][7]  ( .ip(n3113), .ck(clk), .q(
        \ANSWER/mem[2][1][7] ) );
  dp_1 \ANSWER/mem_reg[2][2][7]  ( .ip(n3112), .ck(clk), .q(
        \ANSWER/mem[2][2][7] ) );
  dp_1 \ANSWER/mem_reg[2][3][7]  ( .ip(n3111), .ck(clk), .q(
        \ANSWER/mem[2][3][7] ) );
  dp_1 \ANSWER/mem_reg[2][4][7]  ( .ip(n3110), .ck(clk), .q(
        \ANSWER/mem[2][4][7] ) );
  dp_1 \ANSWER/mem_reg[2][5][7]  ( .ip(n3109), .ck(clk), .q(
        \ANSWER/mem[2][5][7] ) );
  dp_1 \ANSWER/mem_reg[2][6][7]  ( .ip(n3108), .ck(clk), .q(
        \ANSWER/mem[2][6][7] ) );
  dp_1 \ANSWER/mem_reg[2][7][7]  ( .ip(n3107), .ck(clk), .q(
        \ANSWER/mem[2][7][7] ) );
  dp_1 \ANSWER/mem_reg[2][8][7]  ( .ip(n3106), .ck(clk), .q(
        \ANSWER/mem[2][8][7] ) );
  dp_1 \ANSWER/mem_reg[2][9][7]  ( .ip(n3105), .ck(clk), .q(
        \ANSWER/mem[2][9][7] ) );
  dp_1 \ANSWER/mem_reg[3][0][7]  ( .ip(n3104), .ck(clk), .q(
        \ANSWER/mem[3][0][7] ) );
  dp_1 \ANSWER/mem_reg[3][1][7]  ( .ip(n3103), .ck(clk), .q(
        \ANSWER/mem[3][1][7] ) );
  dp_1 \ANSWER/mem_reg[3][2][7]  ( .ip(n3102), .ck(clk), .q(
        \ANSWER/mem[3][2][7] ) );
  dp_1 \ANSWER/mem_reg[3][3][7]  ( .ip(n3101), .ck(clk), .q(
        \ANSWER/mem[3][3][7] ) );
  dp_1 \ANSWER/mem_reg[3][4][7]  ( .ip(n3100), .ck(clk), .q(
        \ANSWER/mem[3][4][7] ) );
  dp_1 \ANSWER/mem_reg[3][5][7]  ( .ip(n3099), .ck(clk), .q(
        \ANSWER/mem[3][5][7] ) );
  dp_1 \ANSWER/mem_reg[3][6][7]  ( .ip(n3098), .ck(clk), .q(
        \ANSWER/mem[3][6][7] ) );
  dp_1 \ANSWER/mem_reg[3][7][7]  ( .ip(n3097), .ck(clk), .q(
        \ANSWER/mem[3][7][7] ) );
  dp_1 \ANSWER/mem_reg[3][8][7]  ( .ip(n3096), .ck(clk), .q(
        \ANSWER/mem[3][8][7] ) );
  dp_1 \ANSWER/mem_reg[3][9][7]  ( .ip(n3095), .ck(clk), .q(
        \ANSWER/mem[3][9][7] ) );
  dp_1 \ANSWER/mem_reg[4][0][7]  ( .ip(n3094), .ck(clk), .q(
        \ANSWER/mem[4][0][7] ) );
  dp_1 \ANSWER/mem_reg[4][1][7]  ( .ip(n3093), .ck(clk), .q(
        \ANSWER/mem[4][1][7] ) );
  dp_1 \ANSWER/mem_reg[4][2][7]  ( .ip(n3092), .ck(clk), .q(
        \ANSWER/mem[4][2][7] ) );
  dp_1 \ANSWER/mem_reg[4][3][7]  ( .ip(n3091), .ck(clk), .q(
        \ANSWER/mem[4][3][7] ) );
  dp_1 \ANSWER/mem_reg[4][4][7]  ( .ip(n3090), .ck(clk), .q(
        \ANSWER/mem[4][4][7] ) );
  dp_1 \ANSWER/mem_reg[4][5][7]  ( .ip(n3089), .ck(clk), .q(
        \ANSWER/mem[4][5][7] ) );
  dp_1 \ANSWER/mem_reg[4][6][7]  ( .ip(n3088), .ck(clk), .q(
        \ANSWER/mem[4][6][7] ) );
  dp_1 \ANSWER/mem_reg[4][7][7]  ( .ip(n3087), .ck(clk), .q(
        \ANSWER/mem[4][7][7] ) );
  dp_1 \ANSWER/mem_reg[4][8][7]  ( .ip(n3086), .ck(clk), .q(
        \ANSWER/mem[4][8][7] ) );
  dp_1 \ANSWER/mem_reg[4][9][7]  ( .ip(n3085), .ck(clk), .q(
        \ANSWER/mem[4][9][7] ) );
  dp_1 \ANSWER/mem_reg[5][0][7]  ( .ip(n3084), .ck(clk), .q(
        \ANSWER/mem[5][0][7] ) );
  dp_1 \ANSWER/mem_reg[5][1][7]  ( .ip(n3083), .ck(clk), .q(
        \ANSWER/mem[5][1][7] ) );
  dp_1 \ANSWER/mem_reg[5][2][7]  ( .ip(n3082), .ck(clk), .q(
        \ANSWER/mem[5][2][7] ) );
  dp_1 \ANSWER/mem_reg[5][3][7]  ( .ip(n3081), .ck(clk), .q(
        \ANSWER/mem[5][3][7] ) );
  dp_1 \ANSWER/mem_reg[5][4][7]  ( .ip(n3080), .ck(clk), .q(
        \ANSWER/mem[5][4][7] ) );
  dp_1 \ANSWER/mem_reg[5][5][7]  ( .ip(n3079), .ck(clk), .q(
        \ANSWER/mem[5][5][7] ) );
  dp_1 \ANSWER/mem_reg[5][6][7]  ( .ip(n3078), .ck(clk), .q(
        \ANSWER/mem[5][6][7] ) );
  dp_1 \ANSWER/mem_reg[5][7][7]  ( .ip(n3077), .ck(clk), .q(
        \ANSWER/mem[5][7][7] ) );
  dp_1 \ANSWER/mem_reg[5][8][7]  ( .ip(n3076), .ck(clk), .q(
        \ANSWER/mem[5][8][7] ) );
  dp_1 \ANSWER/mem_reg[5][9][7]  ( .ip(n3075), .ck(clk), .q(
        \ANSWER/mem[5][9][7] ) );
  dp_1 \ANSWER/mem_reg[6][0][7]  ( .ip(n3074), .ck(clk), .q(
        \ANSWER/mem[6][0][7] ) );
  dp_1 \ANSWER/mem_reg[6][1][7]  ( .ip(n3073), .ck(clk), .q(
        \ANSWER/mem[6][1][7] ) );
  dp_1 \ANSWER/mem_reg[6][2][7]  ( .ip(n3072), .ck(clk), .q(
        \ANSWER/mem[6][2][7] ) );
  dp_1 \ANSWER/mem_reg[6][3][7]  ( .ip(n3071), .ck(clk), .q(
        \ANSWER/mem[6][3][7] ) );
  dp_1 \ANSWER/mem_reg[6][4][7]  ( .ip(n3070), .ck(clk), .q(
        \ANSWER/mem[6][4][7] ) );
  dp_1 \ANSWER/mem_reg[6][5][7]  ( .ip(n3069), .ck(clk), .q(
        \ANSWER/mem[6][5][7] ) );
  dp_1 \ANSWER/mem_reg[6][6][7]  ( .ip(n3068), .ck(clk), .q(
        \ANSWER/mem[6][6][7] ) );
  dp_1 \ANSWER/mem_reg[6][7][7]  ( .ip(n3067), .ck(clk), .q(
        \ANSWER/mem[6][7][7] ) );
  dp_1 \ANSWER/mem_reg[6][8][7]  ( .ip(n3066), .ck(clk), .q(
        \ANSWER/mem[6][8][7] ) );
  dp_1 \ANSWER/mem_reg[6][9][7]  ( .ip(n3065), .ck(clk), .q(
        \ANSWER/mem[6][9][7] ) );
  dp_1 \ANSWER/mem_reg[7][0][7]  ( .ip(n3064), .ck(clk), .q(
        \ANSWER/mem[7][0][7] ) );
  dp_1 \ANSWER/mem_reg[7][1][7]  ( .ip(n3063), .ck(clk), .q(
        \ANSWER/mem[7][1][7] ) );
  dp_1 \ANSWER/mem_reg[7][2][7]  ( .ip(n3062), .ck(clk), .q(
        \ANSWER/mem[7][2][7] ) );
  dp_1 \ANSWER/mem_reg[7][3][7]  ( .ip(n3061), .ck(clk), .q(
        \ANSWER/mem[7][3][7] ) );
  dp_1 \ANSWER/mem_reg[7][4][7]  ( .ip(n3060), .ck(clk), .q(
        \ANSWER/mem[7][4][7] ) );
  dp_1 \ANSWER/mem_reg[7][5][7]  ( .ip(n3059), .ck(clk), .q(
        \ANSWER/mem[7][5][7] ) );
  dp_1 \ANSWER/mem_reg[7][6][7]  ( .ip(n3058), .ck(clk), .q(
        \ANSWER/mem[7][6][7] ) );
  dp_1 \ANSWER/mem_reg[7][7][7]  ( .ip(n3057), .ck(clk), .q(
        \ANSWER/mem[7][7][7] ) );
  dp_1 \ANSWER/mem_reg[7][8][7]  ( .ip(n3056), .ck(clk), .q(
        \ANSWER/mem[7][8][7] ) );
  dp_1 \ANSWER/mem_reg[7][9][7]  ( .ip(n3055), .ck(clk), .q(
        \ANSWER/mem[7][9][7] ) );
  dp_1 \ANSWER/mem_reg[8][0][7]  ( .ip(n3054), .ck(clk), .q(
        \ANSWER/mem[8][0][7] ) );
  dp_1 \ANSWER/mem_reg[8][1][7]  ( .ip(n3053), .ck(clk), .q(
        \ANSWER/mem[8][1][7] ) );
  dp_1 \ANSWER/mem_reg[8][2][7]  ( .ip(n3052), .ck(clk), .q(
        \ANSWER/mem[8][2][7] ) );
  dp_1 \ANSWER/mem_reg[8][3][7]  ( .ip(n3051), .ck(clk), .q(
        \ANSWER/mem[8][3][7] ) );
  dp_1 \ANSWER/mem_reg[8][4][7]  ( .ip(n3050), .ck(clk), .q(
        \ANSWER/mem[8][4][7] ) );
  dp_1 \ANSWER/mem_reg[8][5][7]  ( .ip(n3049), .ck(clk), .q(
        \ANSWER/mem[8][5][7] ) );
  dp_1 \ANSWER/mem_reg[8][6][7]  ( .ip(n3048), .ck(clk), .q(
        \ANSWER/mem[8][6][7] ) );
  dp_1 \ANSWER/mem_reg[8][7][7]  ( .ip(n3047), .ck(clk), .q(
        \ANSWER/mem[8][7][7] ) );
  dp_1 \ANSWER/mem_reg[8][8][7]  ( .ip(n3046), .ck(clk), .q(
        \ANSWER/mem[8][8][7] ) );
  dp_1 \ANSWER/mem_reg[8][9][7]  ( .ip(n3045), .ck(clk), .q(
        \ANSWER/mem[8][9][7] ) );
  dp_1 \ANSWER/mem_reg[9][0][7]  ( .ip(n3044), .ck(clk), .q(
        \ANSWER/mem[9][0][7] ) );
  dp_1 \ANSWER/mem_reg[9][1][7]  ( .ip(n3043), .ck(clk), .q(
        \ANSWER/mem[9][1][7] ) );
  dp_1 \ANSWER/mem_reg[9][2][7]  ( .ip(n3042), .ck(clk), .q(
        \ANSWER/mem[9][2][7] ) );
  dp_1 \ANSWER/mem_reg[9][3][7]  ( .ip(n3041), .ck(clk), .q(
        \ANSWER/mem[9][3][7] ) );
  dp_1 \ANSWER/mem_reg[9][4][7]  ( .ip(n3040), .ck(clk), .q(
        \ANSWER/mem[9][4][7] ) );
  dp_1 \ANSWER/mem_reg[9][5][7]  ( .ip(n3039), .ck(clk), .q(
        \ANSWER/mem[9][5][7] ) );
  dp_1 \ANSWER/mem_reg[9][6][7]  ( .ip(n3038), .ck(clk), .q(
        \ANSWER/mem[9][6][7] ) );
  dp_1 \ANSWER/mem_reg[9][7][7]  ( .ip(n3037), .ck(clk), .q(
        \ANSWER/mem[9][7][7] ) );
  dp_1 \ANSWER/mem_reg[9][8][7]  ( .ip(n3036), .ck(clk), .q(
        \ANSWER/mem[9][8][7] ) );
  dp_1 \ANSWER/mem_reg[9][9][7]  ( .ip(n3035), .ck(clk), .q(
        \ANSWER/mem[9][9][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][0]  ( .ip(n2234), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][0] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][1]  ( .ip(n2233), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][1] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][2]  ( .ip(n2232), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][2] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][3]  ( .ip(n2231), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][3] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][4]  ( .ip(n2230), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][4] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][5]  ( .ip(n2229), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][5] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][6]  ( .ip(n2228), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][6] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][7]  ( .ip(n2227), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][8]  ( .ip(n2226), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][8] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][0]  ( .ip(n2225), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][0] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][1]  ( .ip(n2224), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][1] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][2]  ( .ip(n2223), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][2] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][3]  ( .ip(n2222), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][3] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][4]  ( .ip(n2221), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][4] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][5]  ( .ip(n2220), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][5] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][6]  ( .ip(n2219), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][6] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][7]  ( .ip(n2218), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][8]  ( .ip(n2217), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][8] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][0]  ( .ip(n2216), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][0] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][1]  ( .ip(n2215), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][1] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][2]  ( .ip(n2214), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][2] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][3]  ( .ip(n2213), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][3] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][4]  ( .ip(n2212), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][4] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][5]  ( .ip(n2211), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][5] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][6]  ( .ip(n2210), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][6] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][7]  ( .ip(n2209), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][8]  ( .ip(n2208), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][8] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][0]  ( .ip(n2207), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][0] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][1]  ( .ip(n2206), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][1] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][2]  ( .ip(n2205), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][2] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][3]  ( .ip(n2204), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][3] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][4]  ( .ip(n2203), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][4] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][5]  ( .ip(n2202), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][5] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][6]  ( .ip(n2201), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][6] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][7]  ( .ip(n2200), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][8]  ( .ip(n2199), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][8] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][0]  ( .ip(n2198), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][0] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][1]  ( .ip(n2197), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][1] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][2]  ( .ip(n2196), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][2] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][3]  ( .ip(n2195), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][3] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][4]  ( .ip(n2194), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][4] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][5]  ( .ip(n2193), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][5] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][6]  ( .ip(n2192), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][6] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][7]  ( .ip(n2191), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][8]  ( .ip(n2190), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][8] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][0]  ( .ip(n2189), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][0] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][1]  ( .ip(n2188), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][1] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][2]  ( .ip(n2187), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][2] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][3]  ( .ip(n2186), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][3] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][4]  ( .ip(n2185), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][4] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][5]  ( .ip(n2184), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][5] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][6]  ( .ip(n2183), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][6] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][7]  ( .ip(n2182), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][8]  ( .ip(n2181), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][8] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][0]  ( .ip(n2180), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][0] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][1]  ( .ip(n2179), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][1] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][2]  ( .ip(n2178), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][2] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][3]  ( .ip(n2177), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][3] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][4]  ( .ip(n2176), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][4] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][5]  ( .ip(n2175), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][5] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][6]  ( .ip(n2174), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][6] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][7]  ( .ip(n2173), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][8]  ( .ip(n2172), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][8] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][0]  ( .ip(n2171), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][0] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][1]  ( .ip(n2170), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][1] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][2]  ( .ip(n2169), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][2] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][3]  ( .ip(n2168), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][3] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][4]  ( .ip(n2167), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][4] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][5]  ( .ip(n2166), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][5] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][6]  ( .ip(n2165), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][6] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][7]  ( .ip(n2164), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][8]  ( .ip(n2163), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][8] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][0]  ( .ip(n2162), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][0] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][1]  ( .ip(n2161), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][1] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][2]  ( .ip(n2160), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][2] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][3]  ( .ip(n2159), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][3] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][4]  ( .ip(n2158), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][4] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][5]  ( .ip(n2157), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][5] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][6]  ( .ip(n2156), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][6] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][7]  ( .ip(n2155), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][8]  ( .ip(n2154), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][8] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][0]  ( .ip(n2153), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][0] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][1]  ( .ip(n2152), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][1] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][2]  ( .ip(n2151), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][2] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][3]  ( .ip(n2150), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][3] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][4]  ( .ip(n2149), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][4] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][5]  ( .ip(n2148), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][5] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][6]  ( .ip(n2147), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][6] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][7]  ( .ip(n2146), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][8]  ( .ip(n2145), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][8] ) );
  dp_1 \WEIGHT_2/q_reg[1]  ( .ip(n2143), .ck(clk), .q(q_w2[1]) );
  dp_1 \WEIGHT_2/q_reg[15]  ( .ip(n2129), .ck(clk), .q(q_w2[15]) );
  dp_1 \ROUTEDATA/regData_reg[8]  ( .ip(n2128), .ck(clk), .q(
        \ROUTEDATA/regData [8]) );
  dp_1 \ROUTEDATA/regData_reg[24]  ( .ip(n2127), .ck(clk), .q(
        \ROUTEDATA/regData [24]) );
  dp_1 \ROUTEDATA/regData_reg[40]  ( .ip(n2126), .ck(clk), .q(
        \ROUTEDATA/regData [40]) );
  dp_1 \ROUTEDATA/regData_reg[56]  ( .ip(n2125), .ck(clk), .q(
        \ROUTEDATA/regData [56]) );
  dp_1 \ROUTEDATA/regData_reg[72]  ( .ip(n2124), .ck(clk), .q(
        \ROUTEDATA/regData [72]) );
  dp_1 \ROUTEDATA/regData_reg[88]  ( .ip(n2123), .ck(clk), .q(
        \ROUTEDATA/regData [88]) );
  dp_1 \ROUTEDATA/regData_reg[104]  ( .ip(n2122), .ck(clk), .q(
        \ROUTEDATA/regData [104]) );
  dp_1 \ROUTEDATA/regData_reg[120]  ( .ip(n2121), .ck(clk), .q(
        \ROUTEDATA/regData [120]) );
  dp_1 \ROUTEDATA/regData_reg[136]  ( .ip(n2120), .ck(clk), .q(
        \ROUTEDATA/regData [136]) );
  dp_1 \ROUTEDATA/regData_reg[152]  ( .ip(n2119), .ck(clk), .q(
        \ROUTEDATA/regData [152]) );
  dp_1 \ROUTEDATA/regData_reg[9]  ( .ip(n2118), .ck(clk), .q(
        \ROUTEDATA/regData [9]) );
  dp_1 \ROUTEDATA/regData_reg[25]  ( .ip(n2117), .ck(clk), .q(
        \ROUTEDATA/regData [25]) );
  dp_1 \ROUTEDATA/regData_reg[41]  ( .ip(n2116), .ck(clk), .q(
        \ROUTEDATA/regData [41]) );
  dp_1 \ROUTEDATA/regData_reg[57]  ( .ip(n2115), .ck(clk), .q(
        \ROUTEDATA/regData [57]) );
  dp_1 \ROUTEDATA/regData_reg[73]  ( .ip(n2114), .ck(clk), .q(
        \ROUTEDATA/regData [73]) );
  dp_1 \ROUTEDATA/regData_reg[89]  ( .ip(n2113), .ck(clk), .q(
        \ROUTEDATA/regData [89]) );
  dp_1 \ROUTEDATA/regData_reg[105]  ( .ip(n2112), .ck(clk), .q(
        \ROUTEDATA/regData [105]) );
  dp_1 \ROUTEDATA/regData_reg[121]  ( .ip(n2111), .ck(clk), .q(
        \ROUTEDATA/regData [121]) );
  dp_1 \ROUTEDATA/regData_reg[137]  ( .ip(n2110), .ck(clk), .q(
        \ROUTEDATA/regData [137]) );
  dp_1 \ROUTEDATA/regData_reg[153]  ( .ip(n2109), .ck(clk), .q(
        \ROUTEDATA/regData [153]) );
  dp_1 \ROUTEDATA/regData_reg[10]  ( .ip(n2108), .ck(clk), .q(
        \ROUTEDATA/regData [10]) );
  dp_1 \ROUTEDATA/regData_reg[26]  ( .ip(n2107), .ck(clk), .q(
        \ROUTEDATA/regData [26]) );
  dp_1 \ROUTEDATA/regData_reg[42]  ( .ip(n2106), .ck(clk), .q(
        \ROUTEDATA/regData [42]) );
  dp_1 \ROUTEDATA/regData_reg[58]  ( .ip(n2105), .ck(clk), .q(
        \ROUTEDATA/regData [58]) );
  dp_1 \ROUTEDATA/regData_reg[74]  ( .ip(n2104), .ck(clk), .q(
        \ROUTEDATA/regData [74]) );
  dp_1 \ROUTEDATA/regData_reg[90]  ( .ip(n2103), .ck(clk), .q(
        \ROUTEDATA/regData [90]) );
  dp_1 \ROUTEDATA/regData_reg[106]  ( .ip(n2102), .ck(clk), .q(
        \ROUTEDATA/regData [106]) );
  dp_1 \ROUTEDATA/regData_reg[122]  ( .ip(n2101), .ck(clk), .q(
        \ROUTEDATA/regData [122]) );
  dp_1 \ROUTEDATA/regData_reg[138]  ( .ip(n2100), .ck(clk), .q(
        \ROUTEDATA/regData [138]) );
  dp_1 \ROUTEDATA/regData_reg[154]  ( .ip(n2099), .ck(clk), .q(
        \ROUTEDATA/regData [154]) );
  dp_1 \ROUTEDATA/regData_reg[11]  ( .ip(n2098), .ck(clk), .q(
        \ROUTEDATA/regData [11]) );
  dp_1 \ROUTEDATA/regData_reg[27]  ( .ip(n2097), .ck(clk), .q(
        \ROUTEDATA/regData [27]) );
  dp_1 \ROUTEDATA/regData_reg[43]  ( .ip(n2096), .ck(clk), .q(
        \ROUTEDATA/regData [43]) );
  dp_1 \ROUTEDATA/regData_reg[59]  ( .ip(n2095), .ck(clk), .q(
        \ROUTEDATA/regData [59]) );
  dp_1 \ROUTEDATA/regData_reg[75]  ( .ip(n2094), .ck(clk), .q(
        \ROUTEDATA/regData [75]) );
  dp_1 \ROUTEDATA/regData_reg[91]  ( .ip(n2093), .ck(clk), .q(
        \ROUTEDATA/regData [91]) );
  dp_1 \ROUTEDATA/regData_reg[107]  ( .ip(n2092), .ck(clk), .q(
        \ROUTEDATA/regData [107]) );
  dp_1 \ROUTEDATA/regData_reg[123]  ( .ip(n2091), .ck(clk), .q(
        \ROUTEDATA/regData [123]) );
  dp_1 \ROUTEDATA/regData_reg[139]  ( .ip(n2090), .ck(clk), .q(
        \ROUTEDATA/regData [139]) );
  dp_1 \ROUTEDATA/regData_reg[155]  ( .ip(n2089), .ck(clk), .q(
        \ROUTEDATA/regData [155]) );
  dp_1 \ROUTEDATA/regData_reg[12]  ( .ip(n2088), .ck(clk), .q(
        \ROUTEDATA/regData [12]) );
  dp_1 \ROUTEDATA/regData_reg[28]  ( .ip(n2087), .ck(clk), .q(
        \ROUTEDATA/regData [28]) );
  dp_1 \ROUTEDATA/regData_reg[44]  ( .ip(n2086), .ck(clk), .q(
        \ROUTEDATA/regData [44]) );
  dp_1 \ROUTEDATA/regData_reg[60]  ( .ip(n2085), .ck(clk), .q(
        \ROUTEDATA/regData [60]) );
  dp_1 \ROUTEDATA/regData_reg[76]  ( .ip(n2084), .ck(clk), .q(
        \ROUTEDATA/regData [76]) );
  dp_1 \ROUTEDATA/regData_reg[92]  ( .ip(n2083), .ck(clk), .q(
        \ROUTEDATA/regData [92]) );
  dp_1 \ROUTEDATA/regData_reg[108]  ( .ip(n2082), .ck(clk), .q(
        \ROUTEDATA/regData [108]) );
  dp_1 \ROUTEDATA/regData_reg[124]  ( .ip(n2081), .ck(clk), .q(
        \ROUTEDATA/regData [124]) );
  dp_1 \ROUTEDATA/regData_reg[140]  ( .ip(n2080), .ck(clk), .q(
        \ROUTEDATA/regData [140]) );
  dp_1 \ROUTEDATA/regData_reg[156]  ( .ip(n2079), .ck(clk), .q(
        \ROUTEDATA/regData [156]) );
  dp_1 \ROUTEDATA/regData_reg[13]  ( .ip(n2078), .ck(clk), .q(
        \ROUTEDATA/regData [13]) );
  dp_1 \ROUTEDATA/regData_reg[29]  ( .ip(n2077), .ck(clk), .q(
        \ROUTEDATA/regData [29]) );
  dp_1 \ROUTEDATA/regData_reg[45]  ( .ip(n2076), .ck(clk), .q(
        \ROUTEDATA/regData [45]) );
  dp_1 \ROUTEDATA/regData_reg[61]  ( .ip(n2075), .ck(clk), .q(
        \ROUTEDATA/regData [61]) );
  dp_1 \ROUTEDATA/regData_reg[77]  ( .ip(n2074), .ck(clk), .q(
        \ROUTEDATA/regData [77]) );
  dp_1 \ROUTEDATA/regData_reg[93]  ( .ip(n2073), .ck(clk), .q(
        \ROUTEDATA/regData [93]) );
  dp_1 \ROUTEDATA/regData_reg[109]  ( .ip(n2072), .ck(clk), .q(
        \ROUTEDATA/regData [109]) );
  dp_1 \ROUTEDATA/regData_reg[125]  ( .ip(n2071), .ck(clk), .q(
        \ROUTEDATA/regData [125]) );
  dp_1 \ROUTEDATA/regData_reg[141]  ( .ip(n2070), .ck(clk), .q(
        \ROUTEDATA/regData [141]) );
  dp_1 \ROUTEDATA/regData_reg[157]  ( .ip(n2069), .ck(clk), .q(
        \ROUTEDATA/regData [157]) );
  dp_1 \ROUTEDATA/regData_reg[14]  ( .ip(n2068), .ck(clk), .q(
        \ROUTEDATA/regData [14]) );
  dp_1 \ROUTEDATA/regData_reg[30]  ( .ip(n2067), .ck(clk), .q(
        \ROUTEDATA/regData [30]) );
  dp_1 \ROUTEDATA/regData_reg[46]  ( .ip(n2066), .ck(clk), .q(
        \ROUTEDATA/regData [46]) );
  dp_1 \ROUTEDATA/regData_reg[62]  ( .ip(n2065), .ck(clk), .q(
        \ROUTEDATA/regData [62]) );
  dp_1 \ROUTEDATA/regData_reg[78]  ( .ip(n2064), .ck(clk), .q(
        \ROUTEDATA/regData [78]) );
  dp_1 \ROUTEDATA/regData_reg[94]  ( .ip(n2063), .ck(clk), .q(
        \ROUTEDATA/regData [94]) );
  dp_1 \ROUTEDATA/regData_reg[110]  ( .ip(n2062), .ck(clk), .q(
        \ROUTEDATA/regData [110]) );
  dp_1 \ROUTEDATA/regData_reg[126]  ( .ip(n2061), .ck(clk), .q(
        \ROUTEDATA/regData [126]) );
  dp_1 \ROUTEDATA/regData_reg[142]  ( .ip(n2060), .ck(clk), .q(
        \ROUTEDATA/regData [142]) );
  dp_1 \ROUTEDATA/regData_reg[158]  ( .ip(n2059), .ck(clk), .q(
        \ROUTEDATA/regData [158]) );
  dp_1 \ROUTEDATA/regData_reg[15]  ( .ip(n2058), .ck(clk), .q(
        \ROUTEDATA/regData [15]) );
  dp_1 \ROUTEDATA/regData_reg[31]  ( .ip(n2057), .ck(clk), .q(
        \ROUTEDATA/regData [31]) );
  dp_1 \ROUTEDATA/regData_reg[47]  ( .ip(n2056), .ck(clk), .q(
        \ROUTEDATA/regData [47]) );
  dp_1 \ROUTEDATA/regData_reg[63]  ( .ip(n2055), .ck(clk), .q(
        \ROUTEDATA/regData [63]) );
  dp_1 \ROUTEDATA/regData_reg[79]  ( .ip(n2054), .ck(clk), .q(
        \ROUTEDATA/regData [79]) );
  dp_1 \ROUTEDATA/regData_reg[95]  ( .ip(n2053), .ck(clk), .q(
        \ROUTEDATA/regData [95]) );
  dp_1 \ROUTEDATA/regData_reg[111]  ( .ip(n2052), .ck(clk), .q(
        \ROUTEDATA/regData [111]) );
  dp_1 \ROUTEDATA/regData_reg[127]  ( .ip(n2051), .ck(clk), .q(
        \ROUTEDATA/regData [127]) );
  dp_1 \ROUTEDATA/regData_reg[143]  ( .ip(n2050), .ck(clk), .q(
        \ROUTEDATA/regData [143]) );
  dp_1 \ROUTEDATA/regData_reg[159]  ( .ip(n2049), .ck(clk), .q(
        \ROUTEDATA/regData [159]) );
  dp_1 \ROUTEDATA/regData_reg[0]  ( .ip(n2048), .ck(clk), .q(
        \ROUTEDATA/regData [0]) );
  dp_1 \ROUTEDATA/regData_reg[16]  ( .ip(n2047), .ck(clk), .q(
        \ROUTEDATA/regData [16]) );
  dp_1 \ROUTEDATA/regData_reg[32]  ( .ip(n2046), .ck(clk), .q(
        \ROUTEDATA/regData [32]) );
  dp_1 \ROUTEDATA/regData_reg[48]  ( .ip(n2045), .ck(clk), .q(
        \ROUTEDATA/regData [48]) );
  dp_1 \ROUTEDATA/regData_reg[64]  ( .ip(n2044), .ck(clk), .q(
        \ROUTEDATA/regData [64]) );
  dp_1 \ROUTEDATA/regData_reg[80]  ( .ip(n2043), .ck(clk), .q(
        \ROUTEDATA/regData [80]) );
  dp_1 \ROUTEDATA/regData_reg[96]  ( .ip(n2042), .ck(clk), .q(
        \ROUTEDATA/regData [96]) );
  dp_1 \ROUTEDATA/regData_reg[112]  ( .ip(n2041), .ck(clk), .q(
        \ROUTEDATA/regData [112]) );
  dp_1 \ROUTEDATA/regData_reg[128]  ( .ip(n2040), .ck(clk), .q(
        \ROUTEDATA/regData [128]) );
  dp_1 \ROUTEDATA/regData_reg[144]  ( .ip(n2039), .ck(clk), .q(
        \ROUTEDATA/regData [144]) );
  dp_1 \ROUTEDATA/regData_reg[1]  ( .ip(n2038), .ck(clk), .q(
        \ROUTEDATA/regData [1]) );
  dp_1 \ROUTEDATA/regData_reg[17]  ( .ip(n2037), .ck(clk), .q(
        \ROUTEDATA/regData [17]) );
  dp_1 \ROUTEDATA/regData_reg[33]  ( .ip(n2036), .ck(clk), .q(
        \ROUTEDATA/regData [33]) );
  dp_1 \ROUTEDATA/regData_reg[49]  ( .ip(n2035), .ck(clk), .q(
        \ROUTEDATA/regData [49]) );
  dp_1 \ROUTEDATA/regData_reg[65]  ( .ip(n2034), .ck(clk), .q(
        \ROUTEDATA/regData [65]) );
  dp_1 \ROUTEDATA/regData_reg[81]  ( .ip(n2033), .ck(clk), .q(
        \ROUTEDATA/regData [81]) );
  dp_1 \ROUTEDATA/regData_reg[97]  ( .ip(n2032), .ck(clk), .q(
        \ROUTEDATA/regData [97]) );
  dp_1 \ROUTEDATA/regData_reg[113]  ( .ip(n2031), .ck(clk), .q(
        \ROUTEDATA/regData [113]) );
  dp_1 \ROUTEDATA/regData_reg[129]  ( .ip(n2030), .ck(clk), .q(
        \ROUTEDATA/regData [129]) );
  dp_1 \ROUTEDATA/regData_reg[145]  ( .ip(n2029), .ck(clk), .q(
        \ROUTEDATA/regData [145]) );
  dp_1 \ROUTEDATA/regData_reg[2]  ( .ip(n2028), .ck(clk), .q(
        \ROUTEDATA/regData [2]) );
  dp_1 \ROUTEDATA/regData_reg[18]  ( .ip(n2027), .ck(clk), .q(
        \ROUTEDATA/regData [18]) );
  dp_1 \ROUTEDATA/regData_reg[34]  ( .ip(n2026), .ck(clk), .q(
        \ROUTEDATA/regData [34]) );
  dp_1 \ROUTEDATA/regData_reg[50]  ( .ip(n2025), .ck(clk), .q(
        \ROUTEDATA/regData [50]) );
  dp_1 \ROUTEDATA/regData_reg[66]  ( .ip(n2024), .ck(clk), .q(
        \ROUTEDATA/regData [66]) );
  dp_1 \ROUTEDATA/regData_reg[82]  ( .ip(n2023), .ck(clk), .q(
        \ROUTEDATA/regData [82]) );
  dp_1 \ROUTEDATA/regData_reg[98]  ( .ip(n2022), .ck(clk), .q(
        \ROUTEDATA/regData [98]) );
  dp_1 \ROUTEDATA/regData_reg[114]  ( .ip(n2021), .ck(clk), .q(
        \ROUTEDATA/regData [114]) );
  dp_1 \ROUTEDATA/regData_reg[130]  ( .ip(n2020), .ck(clk), .q(
        \ROUTEDATA/regData [130]) );
  dp_1 \ROUTEDATA/regData_reg[146]  ( .ip(n2019), .ck(clk), .q(
        \ROUTEDATA/regData [146]) );
  dp_1 \ROUTEDATA/regData_reg[3]  ( .ip(n2018), .ck(clk), .q(
        \ROUTEDATA/regData [3]) );
  dp_1 \ROUTEDATA/regData_reg[19]  ( .ip(n2017), .ck(clk), .q(
        \ROUTEDATA/regData [19]) );
  dp_1 \ROUTEDATA/regData_reg[35]  ( .ip(n2016), .ck(clk), .q(
        \ROUTEDATA/regData [35]) );
  dp_1 \ROUTEDATA/regData_reg[51]  ( .ip(n2015), .ck(clk), .q(
        \ROUTEDATA/regData [51]) );
  dp_1 \ROUTEDATA/regData_reg[67]  ( .ip(n2014), .ck(clk), .q(
        \ROUTEDATA/regData [67]) );
  dp_1 \ROUTEDATA/regData_reg[83]  ( .ip(n2013), .ck(clk), .q(
        \ROUTEDATA/regData [83]) );
  dp_1 \ROUTEDATA/regData_reg[99]  ( .ip(n2012), .ck(clk), .q(
        \ROUTEDATA/regData [99]) );
  dp_1 \ROUTEDATA/regData_reg[115]  ( .ip(n2011), .ck(clk), .q(
        \ROUTEDATA/regData [115]) );
  dp_1 \ROUTEDATA/regData_reg[131]  ( .ip(n2010), .ck(clk), .q(
        \ROUTEDATA/regData [131]) );
  dp_1 \ROUTEDATA/regData_reg[147]  ( .ip(n2009), .ck(clk), .q(
        \ROUTEDATA/regData [147]) );
  dp_1 \ROUTEDATA/regData_reg[4]  ( .ip(n2008), .ck(clk), .q(
        \ROUTEDATA/regData [4]) );
  dp_1 \ROUTEDATA/regData_reg[20]  ( .ip(n2007), .ck(clk), .q(
        \ROUTEDATA/regData [20]) );
  dp_1 \ROUTEDATA/regData_reg[36]  ( .ip(n2006), .ck(clk), .q(
        \ROUTEDATA/regData [36]) );
  dp_1 \ROUTEDATA/regData_reg[52]  ( .ip(n2005), .ck(clk), .q(
        \ROUTEDATA/regData [52]) );
  dp_1 \ROUTEDATA/regData_reg[68]  ( .ip(n2004), .ck(clk), .q(
        \ROUTEDATA/regData [68]) );
  dp_1 \ROUTEDATA/regData_reg[84]  ( .ip(n2003), .ck(clk), .q(
        \ROUTEDATA/regData [84]) );
  dp_1 \ROUTEDATA/regData_reg[100]  ( .ip(n2002), .ck(clk), .q(
        \ROUTEDATA/regData [100]) );
  dp_1 \ROUTEDATA/regData_reg[116]  ( .ip(n2001), .ck(clk), .q(
        \ROUTEDATA/regData [116]) );
  dp_1 \ROUTEDATA/regData_reg[132]  ( .ip(n2000), .ck(clk), .q(
        \ROUTEDATA/regData [132]) );
  dp_1 \ROUTEDATA/regData_reg[148]  ( .ip(n1999), .ck(clk), .q(
        \ROUTEDATA/regData [148]) );
  dp_1 \ROUTEDATA/regData_reg[5]  ( .ip(n1998), .ck(clk), .q(
        \ROUTEDATA/regData [5]) );
  dp_1 \ROUTEDATA/regData_reg[21]  ( .ip(n1997), .ck(clk), .q(
        \ROUTEDATA/regData [21]) );
  dp_1 \ROUTEDATA/regData_reg[37]  ( .ip(n1996), .ck(clk), .q(
        \ROUTEDATA/regData [37]) );
  dp_1 \ROUTEDATA/regData_reg[53]  ( .ip(n1995), .ck(clk), .q(
        \ROUTEDATA/regData [53]) );
  dp_1 \ROUTEDATA/regData_reg[69]  ( .ip(n1994), .ck(clk), .q(
        \ROUTEDATA/regData [69]) );
  dp_1 \ROUTEDATA/regData_reg[85]  ( .ip(n1993), .ck(clk), .q(
        \ROUTEDATA/regData [85]) );
  dp_1 \ROUTEDATA/regData_reg[101]  ( .ip(n1992), .ck(clk), .q(
        \ROUTEDATA/regData [101]) );
  dp_1 \ROUTEDATA/regData_reg[117]  ( .ip(n1991), .ck(clk), .q(
        \ROUTEDATA/regData [117]) );
  dp_1 \ROUTEDATA/regData_reg[133]  ( .ip(n1990), .ck(clk), .q(
        \ROUTEDATA/regData [133]) );
  dp_1 \ROUTEDATA/regData_reg[149]  ( .ip(n1989), .ck(clk), .q(
        \ROUTEDATA/regData [149]) );
  dp_1 \ROUTEDATA/regData_reg[6]  ( .ip(n1988), .ck(clk), .q(
        \ROUTEDATA/regData [6]) );
  dp_1 \ROUTEDATA/regData_reg[22]  ( .ip(n1987), .ck(clk), .q(
        \ROUTEDATA/regData [22]) );
  dp_1 \ROUTEDATA/regData_reg[38]  ( .ip(n1986), .ck(clk), .q(
        \ROUTEDATA/regData [38]) );
  dp_1 \ROUTEDATA/regData_reg[54]  ( .ip(n1985), .ck(clk), .q(
        \ROUTEDATA/regData [54]) );
  dp_1 \ROUTEDATA/regData_reg[70]  ( .ip(n1984), .ck(clk), .q(
        \ROUTEDATA/regData [70]) );
  dp_1 \ROUTEDATA/regData_reg[86]  ( .ip(n1983), .ck(clk), .q(
        \ROUTEDATA/regData [86]) );
  dp_1 \ROUTEDATA/regData_reg[102]  ( .ip(n1982), .ck(clk), .q(
        \ROUTEDATA/regData [102]) );
  dp_1 \ROUTEDATA/regData_reg[118]  ( .ip(n1981), .ck(clk), .q(
        \ROUTEDATA/regData [118]) );
  dp_1 \ROUTEDATA/regData_reg[134]  ( .ip(n1980), .ck(clk), .q(
        \ROUTEDATA/regData [134]) );
  dp_1 \ROUTEDATA/regData_reg[150]  ( .ip(n1979), .ck(clk), .q(
        \ROUTEDATA/regData [150]) );
  dp_1 \ROUTEDATA/regData_reg[7]  ( .ip(n1978), .ck(clk), .q(
        \ROUTEDATA/regData [7]) );
  dp_1 \ROUTEDATA/regData_reg[23]  ( .ip(n1977), .ck(clk), .q(
        \ROUTEDATA/regData [23]) );
  dp_1 \ROUTEDATA/regData_reg[39]  ( .ip(n1976), .ck(clk), .q(
        \ROUTEDATA/regData [39]) );
  dp_1 \ROUTEDATA/regData_reg[55]  ( .ip(n1975), .ck(clk), .q(
        \ROUTEDATA/regData [55]) );
  dp_1 \ROUTEDATA/regData_reg[71]  ( .ip(n1974), .ck(clk), .q(
        \ROUTEDATA/regData [71]) );
  dp_1 \ROUTEDATA/regData_reg[87]  ( .ip(n1973), .ck(clk), .q(
        \ROUTEDATA/regData [87]) );
  dp_1 \ROUTEDATA/regData_reg[103]  ( .ip(n1972), .ck(clk), .q(
        \ROUTEDATA/regData [103]) );
  dp_1 \ROUTEDATA/regData_reg[119]  ( .ip(n1971), .ck(clk), .q(
        \ROUTEDATA/regData [119]) );
  dp_1 \ROUTEDATA/regData_reg[135]  ( .ip(n1970), .ck(clk), .q(
        \ROUTEDATA/regData [135]) );
  dp_1 \ROUTEDATA/regData_reg[151]  ( .ip(n1969), .ck(clk), .q(
        \ROUTEDATA/regData [151]) );
  dp_1 \STAGE_1/weightReg_reg[0]  ( .ip(weight1[0]), .ck(clk), .q(
        \STAGE_1/weightReg [0]) );
  dp_1 \STAGE_1/weightReg_reg[15]  ( .ip(weight1[8]), .ck(clk), .q(
        \STAGE_1/weightReg [15]) );
  dp_1 \STAGE_1/weightReg_reg[7]  ( .ip(weight1[7]), .ck(clk), .q(
        \STAGE_1/weightReg [7]) );
  dp_1 \INPUTSRAM/q_reg[8]  ( .ip(\INPUTSRAM/mem_i[0][8] ), .ck(clk), .q(
        m1Inputs[8]) );
  dp_1 \INPUTSRAM/q_reg[2]  ( .ip(\INPUTSRAM/mem_i[0][2] ), .ck(clk), .q(
        m1Inputs[2]) );
  dp_1 \INPUTSRAM/q_reg[4]  ( .ip(\INPUTSRAM/mem_i[0][4] ), .ck(clk), .q(
        m1Inputs[4]) );
  dp_1 \INPUTSRAM/q_reg[56]  ( .ip(\INPUTSRAM/mem_i[3][8] ), .ck(clk), .q(
        m1Inputs[56]) );
  dp_1 \INPUTSRAM/q_reg[24]  ( .ip(\INPUTSRAM/mem_i[1][8] ), .ck(clk), .q(
        m1Inputs[24]) );
  dp_1 \INPUTSRAM/q_reg[88]  ( .ip(\INPUTSRAM/mem_i[5][8] ), .ck(clk), .q(
        m1Inputs[88]) );
  dp_1 \INPUTSRAM/q_reg[136]  ( .ip(\INPUTSRAM/mem_i[8][8] ), .ck(clk), .q(
        m1Inputs[136]) );
  dp_1 \INPUTSRAM/q_reg[98]  ( .ip(\INPUTSRAM/mem_i[6][2] ), .ck(clk), .q(
        m1Inputs[98]) );
  dp_1 \INPUTSRAM/q_reg[50]  ( .ip(\INPUTSRAM/mem_i[3][2] ), .ck(clk), .q(
        m1Inputs[50]) );
  dp_1 \INPUTSRAM/q_reg[146]  ( .ip(\INPUTSRAM/mem_i[9][2] ), .ck(clk), .q(
        m1Inputs[146]) );
  dp_1 \INPUTSRAM/q_reg[82]  ( .ip(\INPUTSRAM/mem_i[5][2] ), .ck(clk), .q(
        m1Inputs[82]) );
  dp_1 \INPUTSRAM/q_reg[66]  ( .ip(\INPUTSRAM/mem_i[4][2] ), .ck(clk), .q(
        m1Inputs[66]) );
  dp_1 \INPUTSRAM/q_reg[18]  ( .ip(\INPUTSRAM/mem_i[1][2] ), .ck(clk), .q(
        m1Inputs[18]) );
  dp_1 \INPUTSRAM/q_reg[130]  ( .ip(\INPUTSRAM/mem_i[8][2] ), .ck(clk), .q(
        m1Inputs[130]) );
  dp_1 \INPUTSRAM/q_reg[34]  ( .ip(\INPUTSRAM/mem_i[2][2] ), .ck(clk), .q(
        m1Inputs[34]) );
  dp_1 \INPUTSRAM/q_reg[114]  ( .ip(\INPUTSRAM/mem_i[7][2] ), .ck(clk), .q(
        m1Inputs[114]) );
  dp_1 \WEIGHT_2/q_reg[14]  ( .ip(n2130), .ck(clk), .q(q_w2[14]) );
  dp_1 \WEIGHT_2/q_reg[12]  ( .ip(n2132), .ck(clk), .q(q_w2[12]) );
  dp_1 \WEIGHT_2/q_reg[11]  ( .ip(n2133), .ck(clk), .q(q_w2[11]) );
  dp_1 \WEIGHT_2/q_reg[9]  ( .ip(n2135), .ck(clk), .q(q_w2[9]) );
  dp_1 \WEIGHT_2/q_reg[10]  ( .ip(n2134), .ck(clk), .q(q_w2[10]) );
  dp_1 \WEIGHT_2/q_reg[13]  ( .ip(n2131), .ck(clk), .q(q_w2[13]) );
  dp_1 \WEIGHT_2/q_reg[8]  ( .ip(n2136), .ck(clk), .q(q_w2[8]) );
  dp_1 \WEIGHT_2/q_reg[6]  ( .ip(n2138), .ck(clk), .q(q_w2[6]) );
  dp_1 \WEIGHT_2/q_reg[5]  ( .ip(n2139), .ck(clk), .q(q_w2[5]) );
  dp_1 \WEIGHT_2/q_reg[7]  ( .ip(n2137), .ck(clk), .q(q_w2[7]) );
  dp_1 \WEIGHT_2/q_reg[4]  ( .ip(n2140), .ck(clk), .q(q_w2[4]) );
  dp_1 \WEIGHT_2/q_reg[0]  ( .ip(n2144), .ck(clk), .q(q_w2[0]) );
  dp_1 \WEIGHT_2/q_reg[2]  ( .ip(n2142), .ck(clk), .q(q_w2[2]) );
  dp_1 \WEIGHT_2/q_reg[3]  ( .ip(n2141), .ck(clk), .q(q_w2[3]) );
  inv_1 U4268 ( .ip(\CNTRL/currentState [0]), .op(n8195) );
  inv_1 U4269 ( .ip(\CNTRL/currentState [1]), .op(n4405) );
  nand2_1 U4270 ( .ip1(n8195), .ip2(n4405), .op(n4442) );
  inv_1 U4271 ( .ip(n4442), .op(n8810) );
  nand2_1 U4272 ( .ip1(\CNTRL/currentState [2]), .ip2(n8810), .op(n8802) );
  inv_1 U4273 ( .ip(\CNTRL/count_10Q [3]), .op(n8285) );
  nor4_1 U4274 ( .ip1(\CNTRL/count_10Q [0]), .ip2(w2SramWeOffChip), .ip3(n8802), .ip4(n8285), .op(n4266) );
  nand2_1 U4275 ( .ip1(n4266), .ip2(\WEIGHT_2/mem_w2[8][2] ), .op(n4069) );
  nand2_1 U4276 ( .ip1(q_w2[2]), .ip2(w2SramWeOffChip), .op(n4068) );
  inv_1 U4277 ( .ip(n8802), .op(n8793) );
  nand2_1 U4278 ( .ip1(n8793), .ip2(\CNTRL/count_10Q [0]), .op(n8784) );
  nor3_1 U4279 ( .ip1(w2SramWeOffChip), .ip2(n8285), .ip3(n8784), .op(n4267)
         );
  nand2_1 U4280 ( .ip1(n4267), .ip2(\WEIGHT_2/mem_w2[9][2] ), .op(n4067) );
  nor2_1 U4281 ( .ip1(n8802), .ip2(n8285), .op(n8786) );
  nor2_1 U4282 ( .ip1(n8786), .ip2(w2SramWeOffChip), .op(n4278) );
  nor2_1 U4283 ( .ip1(w2SramWeOffChip), .ip2(n8784), .op(n4044) );
  or2_1 U4284 ( .ip1(w2SramWeOffChip), .ip2(n4044), .op(n4046) );
  or2_1 U4285 ( .ip1(weight2AddrOffChip[0]), .ip2(n4044), .op(n4045) );
  nand2_1 U4286 ( .ip1(n4046), .ip2(n4045), .op(n4053) );
  inv_1 U4287 ( .ip(n4053), .op(n4060) );
  inv_1 U4288 ( .ip(\CNTRL/count_10Q [1]), .op(n8280) );
  nor2_1 U4289 ( .ip1(n8802), .ip2(n8280), .op(n8781) );
  mux2_1 U4290 ( .ip1(n8781), .ip2(weight2AddrOffChip[1]), .s(w2SramWeOffChip), 
        .op(n4050) );
  inv_1 U4291 ( .ip(n4050), .op(n4047) );
  inv_1 U4292 ( .ip(\CNTRL/count_10Q [2]), .op(n8282) );
  nor2_1 U4293 ( .ip1(n8802), .ip2(n8282), .op(n8778) );
  mux2_1 U4294 ( .ip1(n8778), .ip2(weight2AddrOffChip[2]), .s(w2SramWeOffChip), 
        .op(n4049) );
  nand2_1 U4295 ( .ip1(n4047), .ip2(n4049), .op(n4051) );
  nor2_1 U4296 ( .ip1(n4060), .ip2(n4051), .op(n8547) );
  nand2_1 U4297 ( .ip1(\WEIGHT_2/mem_w2[4][2] ), .ip2(n8547), .op(n4064) );
  or2_1 U4298 ( .ip1(n4049), .ip2(n4047), .op(n4052) );
  nor2_1 U4299 ( .ip1(n4060), .ip2(n4052), .op(n8541) );
  nor2_1 U4300 ( .ip1(n4050), .ip2(n4049), .op(n4048) );
  nand2_1 U4301 ( .ip1(n4053), .ip2(n4048), .op(n8537) );
  inv_1 U4302 ( .ip(n8537), .op(n8560) );
  and2_1 U4303 ( .ip1(n8560), .ip2(\WEIGHT_2/mem_w2[0][2] ), .op(n4059) );
  nand2_1 U4304 ( .ip1(n4060), .ip2(n4048), .op(n8539) );
  inv_1 U4305 ( .ip(n8539), .op(n8562) );
  nand2_1 U4306 ( .ip1(n8562), .ip2(\WEIGHT_2/mem_w2[1][2] ), .op(n4057) );
  nand2_1 U4307 ( .ip1(n4050), .ip2(n4049), .op(n4061) );
  nor2_1 U4308 ( .ip1(n4053), .ip2(n4061), .op(n8556) );
  nand2_1 U4309 ( .ip1(n8556), .ip2(\WEIGHT_2/mem_w2[7][2] ), .op(n4056) );
  nor2_1 U4310 ( .ip1(n4053), .ip2(n4051), .op(n8550) );
  nand2_1 U4311 ( .ip1(n8550), .ip2(\WEIGHT_2/mem_w2[5][2] ), .op(n4055) );
  nor2_1 U4312 ( .ip1(n4053), .ip2(n4052), .op(n8544) );
  nand2_1 U4313 ( .ip1(n8544), .ip2(\WEIGHT_2/mem_w2[3][2] ), .op(n4054) );
  nand4_1 U4314 ( .ip1(n4057), .ip2(n4056), .ip3(n4055), .ip4(n4054), .op(
        n4058) );
  not_ab_or_c_or_d U4315 ( .ip1(n8541), .ip2(\WEIGHT_2/mem_w2[2][2] ), .ip3(
        n4059), .ip4(n4058), .op(n4063) );
  nor2_1 U4316 ( .ip1(n4061), .ip2(n4060), .op(n8553) );
  nand2_1 U4317 ( .ip1(n8553), .ip2(\WEIGHT_2/mem_w2[6][2] ), .op(n4062) );
  nand3_1 U4318 ( .ip1(n4064), .ip2(n4063), .ip3(n4062), .op(n4065) );
  nand2_1 U4319 ( .ip1(n4278), .ip2(n4065), .op(n4066) );
  nand4_1 U4320 ( .ip1(n4069), .ip2(n4068), .ip3(n4067), .ip4(n4066), .op(
        n2142) );
  nand2_1 U4321 ( .ip1(n4266), .ip2(\WEIGHT_2/mem_w2[8][8] ), .op(n4083) );
  nand2_1 U4322 ( .ip1(w2SramWeOffChip), .ip2(q_w2[8]), .op(n4082) );
  nand2_1 U4323 ( .ip1(n4267), .ip2(\WEIGHT_2/mem_w2[9][8] ), .op(n4081) );
  nand2_1 U4324 ( .ip1(n8541), .ip2(\WEIGHT_2/mem_w2[2][8] ), .op(n4078) );
  and2_1 U4325 ( .ip1(n8560), .ip2(\WEIGHT_2/mem_w2[0][8] ), .op(n4075) );
  nand2_1 U4326 ( .ip1(n8556), .ip2(\WEIGHT_2/mem_w2[7][8] ), .op(n4073) );
  nand2_1 U4327 ( .ip1(n8544), .ip2(\WEIGHT_2/mem_w2[3][8] ), .op(n4072) );
  nand2_1 U4328 ( .ip1(n8547), .ip2(\WEIGHT_2/mem_w2[4][8] ), .op(n4071) );
  nand2_1 U4329 ( .ip1(n8562), .ip2(\WEIGHT_2/mem_w2[1][8] ), .op(n4070) );
  nand4_1 U4330 ( .ip1(n4073), .ip2(n4072), .ip3(n4071), .ip4(n4070), .op(
        n4074) );
  not_ab_or_c_or_d U4331 ( .ip1(\WEIGHT_2/mem_w2[5][8] ), .ip2(n8550), .ip3(
        n4075), .ip4(n4074), .op(n4077) );
  nand2_1 U4332 ( .ip1(n8553), .ip2(\WEIGHT_2/mem_w2[6][8] ), .op(n4076) );
  nand3_1 U4333 ( .ip1(n4078), .ip2(n4077), .ip3(n4076), .op(n4079) );
  nand2_1 U4334 ( .ip1(n4278), .ip2(n4079), .op(n4080) );
  nand4_1 U4335 ( .ip1(n4083), .ip2(n4082), .ip3(n4081), .ip4(n4080), .op(
        n2136) );
  nand2_1 U4336 ( .ip1(q_w2[3]), .ip2(w2SramWeOffChip), .op(n4097) );
  nand2_1 U4337 ( .ip1(n4266), .ip2(\WEIGHT_2/mem_w2[8][3] ), .op(n4096) );
  nand2_1 U4338 ( .ip1(n4267), .ip2(\WEIGHT_2/mem_w2[9][3] ), .op(n4095) );
  nand2_1 U4339 ( .ip1(n8544), .ip2(\WEIGHT_2/mem_w2[3][3] ), .op(n4092) );
  and2_1 U4340 ( .ip1(n8560), .ip2(\WEIGHT_2/mem_w2[0][3] ), .op(n4089) );
  nand2_1 U4341 ( .ip1(n8556), .ip2(\WEIGHT_2/mem_w2[7][3] ), .op(n4087) );
  nand2_1 U4342 ( .ip1(n8547), .ip2(\WEIGHT_2/mem_w2[4][3] ), .op(n4086) );
  nand2_1 U4343 ( .ip1(n8562), .ip2(\WEIGHT_2/mem_w2[1][3] ), .op(n4085) );
  nand2_1 U4344 ( .ip1(n8550), .ip2(\WEIGHT_2/mem_w2[5][3] ), .op(n4084) );
  nand4_1 U4345 ( .ip1(n4087), .ip2(n4086), .ip3(n4085), .ip4(n4084), .op(
        n4088) );
  not_ab_or_c_or_d U4346 ( .ip1(\WEIGHT_2/mem_w2[2][3] ), .ip2(n8541), .ip3(
        n4089), .ip4(n4088), .op(n4091) );
  nand2_1 U4347 ( .ip1(n8553), .ip2(\WEIGHT_2/mem_w2[6][3] ), .op(n4090) );
  nand3_1 U4348 ( .ip1(n4092), .ip2(n4091), .ip3(n4090), .op(n4093) );
  nand2_1 U4349 ( .ip1(n4278), .ip2(n4093), .op(n4094) );
  nand4_1 U4350 ( .ip1(n4097), .ip2(n4096), .ip3(n4095), .ip4(n4094), .op(
        n2141) );
  nand2_1 U4351 ( .ip1(n4266), .ip2(\WEIGHT_2/mem_w2[8][12] ), .op(n4111) );
  nand2_1 U4352 ( .ip1(w2SramWeOffChip), .ip2(q_w2[12]), .op(n4110) );
  nand2_1 U4353 ( .ip1(n4267), .ip2(\WEIGHT_2/mem_w2[9][12] ), .op(n4109) );
  nand2_1 U4354 ( .ip1(n8544), .ip2(\WEIGHT_2/mem_w2[3][12] ), .op(n4106) );
  and2_1 U4355 ( .ip1(n8560), .ip2(\WEIGHT_2/mem_w2[0][12] ), .op(n4103) );
  nand2_1 U4356 ( .ip1(n8556), .ip2(\WEIGHT_2/mem_w2[7][12] ), .op(n4101) );
  nand2_1 U4357 ( .ip1(n8553), .ip2(\WEIGHT_2/mem_w2[6][12] ), .op(n4100) );
  nand2_1 U4358 ( .ip1(n8562), .ip2(\WEIGHT_2/mem_w2[1][12] ), .op(n4099) );
  nand2_1 U4359 ( .ip1(n8550), .ip2(\WEIGHT_2/mem_w2[5][12] ), .op(n4098) );
  nand4_1 U4360 ( .ip1(n4101), .ip2(n4100), .ip3(n4099), .ip4(n4098), .op(
        n4102) );
  not_ab_or_c_or_d U4361 ( .ip1(\WEIGHT_2/mem_w2[2][12] ), .ip2(n8541), .ip3(
        n4103), .ip4(n4102), .op(n4105) );
  nand2_1 U4362 ( .ip1(n8547), .ip2(\WEIGHT_2/mem_w2[4][12] ), .op(n4104) );
  nand3_1 U4363 ( .ip1(n4106), .ip2(n4105), .ip3(n4104), .op(n4107) );
  nand2_1 U4364 ( .ip1(n4278), .ip2(n4107), .op(n4108) );
  nand4_1 U4365 ( .ip1(n4111), .ip2(n4110), .ip3(n4109), .ip4(n4108), .op(
        n2132) );
  nand2_1 U4366 ( .ip1(w2SramWeOffChip), .ip2(q_w2[7]), .op(n4125) );
  nand2_1 U4367 ( .ip1(n4266), .ip2(\WEIGHT_2/mem_w2[8][7] ), .op(n4124) );
  nand2_1 U4368 ( .ip1(n4267), .ip2(\WEIGHT_2/mem_w2[9][7] ), .op(n4123) );
  nand2_1 U4369 ( .ip1(n8544), .ip2(\WEIGHT_2/mem_w2[3][7] ), .op(n4120) );
  and2_1 U4370 ( .ip1(n8560), .ip2(\WEIGHT_2/mem_w2[0][7] ), .op(n4117) );
  nand2_1 U4371 ( .ip1(n8556), .ip2(\WEIGHT_2/mem_w2[7][7] ), .op(n4115) );
  nand2_1 U4372 ( .ip1(n8550), .ip2(\WEIGHT_2/mem_w2[5][7] ), .op(n4114) );
  nand2_1 U4373 ( .ip1(n8553), .ip2(\WEIGHT_2/mem_w2[6][7] ), .op(n4113) );
  nand2_1 U4374 ( .ip1(n8547), .ip2(\WEIGHT_2/mem_w2[4][7] ), .op(n4112) );
  nand4_1 U4375 ( .ip1(n4115), .ip2(n4114), .ip3(n4113), .ip4(n4112), .op(
        n4116) );
  not_ab_or_c_or_d U4376 ( .ip1(\WEIGHT_2/mem_w2[1][7] ), .ip2(n8562), .ip3(
        n4117), .ip4(n4116), .op(n4119) );
  nand2_1 U4377 ( .ip1(n8541), .ip2(\WEIGHT_2/mem_w2[2][7] ), .op(n4118) );
  nand3_1 U4378 ( .ip1(n4120), .ip2(n4119), .ip3(n4118), .op(n4121) );
  nand2_1 U4379 ( .ip1(n4278), .ip2(n4121), .op(n4122) );
  nand4_1 U4380 ( .ip1(n4125), .ip2(n4124), .ip3(n4123), .ip4(n4122), .op(
        n2137) );
  nand2_1 U4381 ( .ip1(w2SramWeOffChip), .ip2(q_w2[11]), .op(n4139) );
  nand2_1 U4382 ( .ip1(n4266), .ip2(\WEIGHT_2/mem_w2[8][11] ), .op(n4138) );
  nand2_1 U4383 ( .ip1(n4267), .ip2(\WEIGHT_2/mem_w2[9][11] ), .op(n4137) );
  nand2_1 U4384 ( .ip1(\WEIGHT_2/mem_w2[2][11] ), .ip2(n8541), .op(n4134) );
  and2_1 U4385 ( .ip1(n8560), .ip2(\WEIGHT_2/mem_w2[0][11] ), .op(n4131) );
  nand2_1 U4386 ( .ip1(n8544), .ip2(\WEIGHT_2/mem_w2[3][11] ), .op(n4129) );
  nand2_1 U4387 ( .ip1(n8556), .ip2(\WEIGHT_2/mem_w2[7][11] ), .op(n4128) );
  nand2_1 U4388 ( .ip1(n8553), .ip2(\WEIGHT_2/mem_w2[6][11] ), .op(n4127) );
  nand2_1 U4389 ( .ip1(n8562), .ip2(\WEIGHT_2/mem_w2[1][11] ), .op(n4126) );
  nand4_1 U4390 ( .ip1(n4129), .ip2(n4128), .ip3(n4127), .ip4(n4126), .op(
        n4130) );
  not_ab_or_c_or_d U4391 ( .ip1(\WEIGHT_2/mem_w2[4][11] ), .ip2(n8547), .ip3(
        n4131), .ip4(n4130), .op(n4133) );
  nand2_1 U4392 ( .ip1(n8550), .ip2(\WEIGHT_2/mem_w2[5][11] ), .op(n4132) );
  nand3_1 U4393 ( .ip1(n4134), .ip2(n4133), .ip3(n4132), .op(n4135) );
  nand2_1 U4394 ( .ip1(n4278), .ip2(n4135), .op(n4136) );
  nand4_1 U4395 ( .ip1(n4139), .ip2(n4138), .ip3(n4137), .ip4(n4136), .op(
        n2133) );
  nand2_1 U4396 ( .ip1(w2SramWeOffChip), .ip2(q_w2[5]), .op(n4153) );
  nand2_1 U4397 ( .ip1(n4266), .ip2(\WEIGHT_2/mem_w2[8][5] ), .op(n4152) );
  nand2_1 U4398 ( .ip1(n4267), .ip2(\WEIGHT_2/mem_w2[9][5] ), .op(n4151) );
  nand2_1 U4399 ( .ip1(\WEIGHT_2/mem_w2[7][5] ), .ip2(n8556), .op(n4148) );
  and2_1 U4400 ( .ip1(n8560), .ip2(\WEIGHT_2/mem_w2[0][5] ), .op(n4145) );
  nand2_1 U4401 ( .ip1(n8541), .ip2(\WEIGHT_2/mem_w2[2][5] ), .op(n4143) );
  nand2_1 U4402 ( .ip1(n8544), .ip2(\WEIGHT_2/mem_w2[3][5] ), .op(n4142) );
  nand2_1 U4403 ( .ip1(n8562), .ip2(\WEIGHT_2/mem_w2[1][5] ), .op(n4141) );
  nand2_1 U4404 ( .ip1(n8550), .ip2(\WEIGHT_2/mem_w2[5][5] ), .op(n4140) );
  nand4_1 U4405 ( .ip1(n4143), .ip2(n4142), .ip3(n4141), .ip4(n4140), .op(
        n4144) );
  not_ab_or_c_or_d U4406 ( .ip1(n8547), .ip2(\WEIGHT_2/mem_w2[4][5] ), .ip3(
        n4145), .ip4(n4144), .op(n4147) );
  nand2_1 U4407 ( .ip1(n8553), .ip2(\WEIGHT_2/mem_w2[6][5] ), .op(n4146) );
  nand3_1 U4408 ( .ip1(n4148), .ip2(n4147), .ip3(n4146), .op(n4149) );
  nand2_1 U4409 ( .ip1(n4278), .ip2(n4149), .op(n4150) );
  nand4_1 U4410 ( .ip1(n4153), .ip2(n4152), .ip3(n4151), .ip4(n4150), .op(
        n2139) );
  nand2_1 U4411 ( .ip1(n4266), .ip2(\WEIGHT_2/mem_w2[8][0] ), .op(n4167) );
  nand2_1 U4412 ( .ip1(q_w2[0]), .ip2(w2SramWeOffChip), .op(n4166) );
  nand2_1 U4413 ( .ip1(n4267), .ip2(\WEIGHT_2/mem_w2[9][0] ), .op(n4165) );
  nand2_1 U4414 ( .ip1(n8541), .ip2(\WEIGHT_2/mem_w2[2][0] ), .op(n4162) );
  and2_1 U4415 ( .ip1(n8560), .ip2(\WEIGHT_2/mem_w2[0][0] ), .op(n4159) );
  nand2_1 U4416 ( .ip1(n8556), .ip2(\WEIGHT_2/mem_w2[7][0] ), .op(n4157) );
  nand2_1 U4417 ( .ip1(n8544), .ip2(\WEIGHT_2/mem_w2[3][0] ), .op(n4156) );
  nand2_1 U4418 ( .ip1(n8550), .ip2(\WEIGHT_2/mem_w2[5][0] ), .op(n4155) );
  nand2_1 U4419 ( .ip1(n8553), .ip2(\WEIGHT_2/mem_w2[6][0] ), .op(n4154) );
  nand4_1 U4420 ( .ip1(n4157), .ip2(n4156), .ip3(n4155), .ip4(n4154), .op(
        n4158) );
  not_ab_or_c_or_d U4421 ( .ip1(n8562), .ip2(\WEIGHT_2/mem_w2[1][0] ), .ip3(
        n4159), .ip4(n4158), .op(n4161) );
  nand2_1 U4422 ( .ip1(n8547), .ip2(\WEIGHT_2/mem_w2[4][0] ), .op(n4160) );
  nand3_1 U4423 ( .ip1(n4162), .ip2(n4161), .ip3(n4160), .op(n4163) );
  nand2_1 U4424 ( .ip1(n4278), .ip2(n4163), .op(n4164) );
  nand4_1 U4425 ( .ip1(n4167), .ip2(n4166), .ip3(n4165), .ip4(n4164), .op(
        n2144) );
  nand2_1 U4426 ( .ip1(n4266), .ip2(\WEIGHT_2/mem_w2[8][10] ), .op(n4181) );
  nand2_1 U4427 ( .ip1(w2SramWeOffChip), .ip2(q_w2[10]), .op(n4180) );
  nand2_1 U4428 ( .ip1(n4267), .ip2(\WEIGHT_2/mem_w2[9][10] ), .op(n4179) );
  nand2_1 U4429 ( .ip1(n8556), .ip2(\WEIGHT_2/mem_w2[7][10] ), .op(n4176) );
  and2_1 U4430 ( .ip1(n8560), .ip2(\WEIGHT_2/mem_w2[0][10] ), .op(n4173) );
  nand2_1 U4431 ( .ip1(n8547), .ip2(\WEIGHT_2/mem_w2[4][10] ), .op(n4171) );
  nand2_1 U4432 ( .ip1(n8562), .ip2(\WEIGHT_2/mem_w2[1][10] ), .op(n4170) );
  nand2_1 U4433 ( .ip1(n8553), .ip2(\WEIGHT_2/mem_w2[6][10] ), .op(n4169) );
  nand2_1 U4434 ( .ip1(n8544), .ip2(\WEIGHT_2/mem_w2[3][10] ), .op(n4168) );
  nand4_1 U4435 ( .ip1(n4171), .ip2(n4170), .ip3(n4169), .ip4(n4168), .op(
        n4172) );
  not_ab_or_c_or_d U4436 ( .ip1(n8550), .ip2(\WEIGHT_2/mem_w2[5][10] ), .ip3(
        n4173), .ip4(n4172), .op(n4175) );
  nand2_1 U4437 ( .ip1(n8541), .ip2(\WEIGHT_2/mem_w2[2][10] ), .op(n4174) );
  nand3_1 U4438 ( .ip1(n4176), .ip2(n4175), .ip3(n4174), .op(n4177) );
  nand2_1 U4439 ( .ip1(n4278), .ip2(n4177), .op(n4178) );
  nand4_1 U4440 ( .ip1(n4181), .ip2(n4180), .ip3(n4179), .ip4(n4178), .op(
        n2134) );
  nand2_1 U4441 ( .ip1(n4266), .ip2(\WEIGHT_2/mem_w2[8][13] ), .op(n4195) );
  nand2_1 U4442 ( .ip1(w2SramWeOffChip), .ip2(q_w2[13]), .op(n4194) );
  nand2_1 U4443 ( .ip1(n4267), .ip2(\WEIGHT_2/mem_w2[9][13] ), .op(n4193) );
  nand2_1 U4444 ( .ip1(\WEIGHT_2/mem_w2[3][13] ), .ip2(n8544), .op(n4190) );
  and2_1 U4445 ( .ip1(n8560), .ip2(\WEIGHT_2/mem_w2[0][13] ), .op(n4187) );
  nand2_1 U4446 ( .ip1(n8541), .ip2(\WEIGHT_2/mem_w2[2][13] ), .op(n4185) );
  nand2_1 U4447 ( .ip1(n8547), .ip2(\WEIGHT_2/mem_w2[4][13] ), .op(n4184) );
  nand2_1 U4448 ( .ip1(n8562), .ip2(\WEIGHT_2/mem_w2[1][13] ), .op(n4183) );
  nand2_1 U4449 ( .ip1(n8556), .ip2(\WEIGHT_2/mem_w2[7][13] ), .op(n4182) );
  nand4_1 U4450 ( .ip1(n4185), .ip2(n4184), .ip3(n4183), .ip4(n4182), .op(
        n4186) );
  not_ab_or_c_or_d U4451 ( .ip1(n8550), .ip2(\WEIGHT_2/mem_w2[5][13] ), .ip3(
        n4187), .ip4(n4186), .op(n4189) );
  nand2_1 U4452 ( .ip1(n8553), .ip2(\WEIGHT_2/mem_w2[6][13] ), .op(n4188) );
  nand3_1 U4453 ( .ip1(n4190), .ip2(n4189), .ip3(n4188), .op(n4191) );
  nand2_1 U4454 ( .ip1(n4278), .ip2(n4191), .op(n4192) );
  nand4_1 U4455 ( .ip1(n4195), .ip2(n4194), .ip3(n4193), .ip4(n4192), .op(
        n2131) );
  nand2_1 U4456 ( .ip1(w2SramWeOffChip), .ip2(q_w2[4]), .op(n4209) );
  nand2_1 U4457 ( .ip1(n4266), .ip2(\WEIGHT_2/mem_w2[8][4] ), .op(n4208) );
  nand2_1 U4458 ( .ip1(n4267), .ip2(\WEIGHT_2/mem_w2[9][4] ), .op(n4207) );
  nand2_1 U4459 ( .ip1(\WEIGHT_2/mem_w2[7][4] ), .ip2(n8556), .op(n4204) );
  and2_1 U4460 ( .ip1(n8560), .ip2(\WEIGHT_2/mem_w2[0][4] ), .op(n4201) );
  nand2_1 U4461 ( .ip1(n8562), .ip2(\WEIGHT_2/mem_w2[1][4] ), .op(n4199) );
  nand2_1 U4462 ( .ip1(n8547), .ip2(\WEIGHT_2/mem_w2[4][4] ), .op(n4198) );
  nand2_1 U4463 ( .ip1(n8541), .ip2(\WEIGHT_2/mem_w2[2][4] ), .op(n4197) );
  nand2_1 U4464 ( .ip1(n8553), .ip2(\WEIGHT_2/mem_w2[6][4] ), .op(n4196) );
  nand4_1 U4465 ( .ip1(n4199), .ip2(n4198), .ip3(n4197), .ip4(n4196), .op(
        n4200) );
  not_ab_or_c_or_d U4466 ( .ip1(n8550), .ip2(\WEIGHT_2/mem_w2[5][4] ), .ip3(
        n4201), .ip4(n4200), .op(n4203) );
  nand2_1 U4467 ( .ip1(n8544), .ip2(\WEIGHT_2/mem_w2[3][4] ), .op(n4202) );
  nand3_1 U4468 ( .ip1(n4204), .ip2(n4203), .ip3(n4202), .op(n4205) );
  nand2_1 U4469 ( .ip1(n4278), .ip2(n4205), .op(n4206) );
  nand4_1 U4470 ( .ip1(n4209), .ip2(n4208), .ip3(n4207), .ip4(n4206), .op(
        n2140) );
  nand2_1 U4471 ( .ip1(n4266), .ip2(\WEIGHT_2/mem_w2[8][1] ), .op(n4223) );
  nand2_1 U4472 ( .ip1(q_w2[1]), .ip2(w2SramWeOffChip), .op(n4222) );
  nand2_1 U4473 ( .ip1(n4267), .ip2(\WEIGHT_2/mem_w2[9][1] ), .op(n4221) );
  nand2_1 U4474 ( .ip1(\WEIGHT_2/mem_w2[7][1] ), .ip2(n8556), .op(n4218) );
  and2_1 U4475 ( .ip1(n8560), .ip2(\WEIGHT_2/mem_w2[0][1] ), .op(n4215) );
  nand2_1 U4476 ( .ip1(n8541), .ip2(\WEIGHT_2/mem_w2[2][1] ), .op(n4213) );
  nand2_1 U4477 ( .ip1(n8553), .ip2(\WEIGHT_2/mem_w2[6][1] ), .op(n4212) );
  nand2_1 U4478 ( .ip1(n8562), .ip2(\WEIGHT_2/mem_w2[1][1] ), .op(n4211) );
  nand2_1 U4479 ( .ip1(n8550), .ip2(\WEIGHT_2/mem_w2[5][1] ), .op(n4210) );
  nand4_1 U4480 ( .ip1(n4213), .ip2(n4212), .ip3(n4211), .ip4(n4210), .op(
        n4214) );
  not_ab_or_c_or_d U4481 ( .ip1(n8547), .ip2(\WEIGHT_2/mem_w2[4][1] ), .ip3(
        n4215), .ip4(n4214), .op(n4217) );
  nand2_1 U4482 ( .ip1(n8544), .ip2(\WEIGHT_2/mem_w2[3][1] ), .op(n4216) );
  nand3_1 U4483 ( .ip1(n4218), .ip2(n4217), .ip3(n4216), .op(n4219) );
  nand2_1 U4484 ( .ip1(n4278), .ip2(n4219), .op(n4220) );
  nand4_1 U4485 ( .ip1(n4223), .ip2(n4222), .ip3(n4221), .ip4(n4220), .op(
        n2143) );
  nand2_1 U4486 ( .ip1(w2SramWeOffChip), .ip2(q_w2[9]), .op(n4237) );
  nand2_1 U4487 ( .ip1(n4266), .ip2(\WEIGHT_2/mem_w2[8][9] ), .op(n4236) );
  nand2_1 U4488 ( .ip1(n4267), .ip2(\WEIGHT_2/mem_w2[9][9] ), .op(n4235) );
  nand2_1 U4489 ( .ip1(\WEIGHT_2/mem_w2[7][9] ), .ip2(n8556), .op(n4232) );
  and2_1 U4490 ( .ip1(n8560), .ip2(\WEIGHT_2/mem_w2[0][9] ), .op(n4229) );
  nand2_1 U4491 ( .ip1(n8562), .ip2(\WEIGHT_2/mem_w2[1][9] ), .op(n4227) );
  nand2_1 U4492 ( .ip1(n8544), .ip2(\WEIGHT_2/mem_w2[3][9] ), .op(n4226) );
  nand2_1 U4493 ( .ip1(n8541), .ip2(\WEIGHT_2/mem_w2[2][9] ), .op(n4225) );
  nand2_1 U4494 ( .ip1(n8553), .ip2(\WEIGHT_2/mem_w2[6][9] ), .op(n4224) );
  nand4_1 U4495 ( .ip1(n4227), .ip2(n4226), .ip3(n4225), .ip4(n4224), .op(
        n4228) );
  not_ab_or_c_or_d U4496 ( .ip1(n8550), .ip2(\WEIGHT_2/mem_w2[5][9] ), .ip3(
        n4229), .ip4(n4228), .op(n4231) );
  nand2_1 U4497 ( .ip1(n8547), .ip2(\WEIGHT_2/mem_w2[4][9] ), .op(n4230) );
  nand3_1 U4498 ( .ip1(n4232), .ip2(n4231), .ip3(n4230), .op(n4233) );
  nand2_1 U4499 ( .ip1(n4278), .ip2(n4233), .op(n4234) );
  nand4_1 U4500 ( .ip1(n4237), .ip2(n4236), .ip3(n4235), .ip4(n4234), .op(
        n2135) );
  nand2_1 U4501 ( .ip1(w2SramWeOffChip), .ip2(q_w2[6]), .op(n4251) );
  nand2_1 U4502 ( .ip1(n4266), .ip2(\WEIGHT_2/mem_w2[8][6] ), .op(n4250) );
  nand2_1 U4503 ( .ip1(n4267), .ip2(\WEIGHT_2/mem_w2[9][6] ), .op(n4249) );
  nand2_1 U4504 ( .ip1(n8550), .ip2(\WEIGHT_2/mem_w2[5][6] ), .op(n4246) );
  and2_1 U4505 ( .ip1(n8560), .ip2(\WEIGHT_2/mem_w2[0][6] ), .op(n4243) );
  nand2_1 U4506 ( .ip1(n8553), .ip2(\WEIGHT_2/mem_w2[6][6] ), .op(n4241) );
  nand2_1 U4507 ( .ip1(n8541), .ip2(\WEIGHT_2/mem_w2[2][6] ), .op(n4240) );
  nand2_1 U4508 ( .ip1(n8544), .ip2(\WEIGHT_2/mem_w2[3][6] ), .op(n4239) );
  nand2_1 U4509 ( .ip1(n8547), .ip2(\WEIGHT_2/mem_w2[4][6] ), .op(n4238) );
  nand4_1 U4510 ( .ip1(n4241), .ip2(n4240), .ip3(n4239), .ip4(n4238), .op(
        n4242) );
  not_ab_or_c_or_d U4511 ( .ip1(n8556), .ip2(\WEIGHT_2/mem_w2[7][6] ), .ip3(
        n4243), .ip4(n4242), .op(n4245) );
  nand2_1 U4512 ( .ip1(n8562), .ip2(\WEIGHT_2/mem_w2[1][6] ), .op(n4244) );
  nand3_1 U4513 ( .ip1(n4246), .ip2(n4245), .ip3(n4244), .op(n4247) );
  nand2_1 U4514 ( .ip1(n4278), .ip2(n4247), .op(n4248) );
  nand4_1 U4515 ( .ip1(n4251), .ip2(n4250), .ip3(n4249), .ip4(n4248), .op(
        n2138) );
  nand2_1 U4516 ( .ip1(w2SramWeOffChip), .ip2(q_w2[15]), .op(n4265) );
  nand2_1 U4517 ( .ip1(n4266), .ip2(\WEIGHT_2/mem_w2[8][15] ), .op(n4264) );
  nand2_1 U4518 ( .ip1(n4267), .ip2(\WEIGHT_2/mem_w2[9][15] ), .op(n4263) );
  nand2_1 U4519 ( .ip1(\WEIGHT_2/mem_w2[3][15] ), .ip2(n8544), .op(n4260) );
  and2_1 U4520 ( .ip1(n8560), .ip2(\WEIGHT_2/mem_w2[0][15] ), .op(n4257) );
  nand2_1 U4521 ( .ip1(n8550), .ip2(\WEIGHT_2/mem_w2[5][15] ), .op(n4255) );
  nand2_1 U4522 ( .ip1(n8541), .ip2(\WEIGHT_2/mem_w2[2][15] ), .op(n4254) );
  nand2_1 U4523 ( .ip1(n8547), .ip2(\WEIGHT_2/mem_w2[4][15] ), .op(n4253) );
  nand2_1 U4524 ( .ip1(n8562), .ip2(\WEIGHT_2/mem_w2[1][15] ), .op(n4252) );
  nand4_1 U4525 ( .ip1(n4255), .ip2(n4254), .ip3(n4253), .ip4(n4252), .op(
        n4256) );
  not_ab_or_c_or_d U4526 ( .ip1(n8556), .ip2(\WEIGHT_2/mem_w2[7][15] ), .ip3(
        n4257), .ip4(n4256), .op(n4259) );
  nand2_1 U4527 ( .ip1(n8553), .ip2(\WEIGHT_2/mem_w2[6][15] ), .op(n4258) );
  nand3_1 U4528 ( .ip1(n4260), .ip2(n4259), .ip3(n4258), .op(n4261) );
  nand2_1 U4529 ( .ip1(n4278), .ip2(n4261), .op(n4262) );
  nand4_1 U4530 ( .ip1(n4265), .ip2(n4264), .ip3(n4263), .ip4(n4262), .op(
        n2129) );
  nand2_1 U4531 ( .ip1(n4266), .ip2(\WEIGHT_2/mem_w2[8][14] ), .op(n4282) );
  nand2_1 U4532 ( .ip1(w2SramWeOffChip), .ip2(q_w2[14]), .op(n4281) );
  nand2_1 U4533 ( .ip1(n4267), .ip2(\WEIGHT_2/mem_w2[9][14] ), .op(n4280) );
  nand2_1 U4534 ( .ip1(\WEIGHT_2/mem_w2[7][14] ), .ip2(n8556), .op(n4276) );
  and2_1 U4535 ( .ip1(n8560), .ip2(\WEIGHT_2/mem_w2[0][14] ), .op(n4273) );
  nand2_1 U4536 ( .ip1(n8562), .ip2(\WEIGHT_2/mem_w2[1][14] ), .op(n4271) );
  nand2_1 U4537 ( .ip1(n8553), .ip2(\WEIGHT_2/mem_w2[6][14] ), .op(n4270) );
  nand2_1 U4538 ( .ip1(n8550), .ip2(\WEIGHT_2/mem_w2[5][14] ), .op(n4269) );
  nand2_1 U4539 ( .ip1(n8541), .ip2(\WEIGHT_2/mem_w2[2][14] ), .op(n4268) );
  nand4_1 U4540 ( .ip1(n4271), .ip2(n4270), .ip3(n4269), .ip4(n4268), .op(
        n4272) );
  not_ab_or_c_or_d U4541 ( .ip1(n8547), .ip2(\WEIGHT_2/mem_w2[4][14] ), .ip3(
        n4273), .ip4(n4272), .op(n4275) );
  nand2_1 U4542 ( .ip1(n8544), .ip2(\WEIGHT_2/mem_w2[3][14] ), .op(n4274) );
  nand3_1 U4543 ( .ip1(n4276), .ip2(n4275), .ip3(n4274), .op(n4277) );
  nand2_1 U4544 ( .ip1(n4278), .ip2(n4277), .op(n4279) );
  nand4_1 U4545 ( .ip1(n4282), .ip2(n4281), .ip3(n4280), .ip4(n4279), .op(
        n2130) );
  inv_1 U4546 ( .ip(rdata[8]), .op(n9486) );
  inv_1 U4547 ( .ip(m2DataIn[8]), .op(n9817) );
  nand3_1 U4548 ( .ip1(\CNTRL/currentState [2]), .ip2(\CNTRL/currentState [1]), 
        .ip3(n8195), .op(n4293) );
  mux2_1 U4549 ( .ip1(n9486), .ip2(n9817), .s(n4293), .op(n4285) );
  mux2_1 U4550 ( .ip1(rdata[15]), .ip2(m2DataIn[15]), .s(n4293), .op(
        \sig_in[15] ) );
  inv_1 U4551 ( .ip(\sig_in[15] ), .op(n4328) );
  inv_1 U4552 ( .ip(rdata[6]), .op(n9216) );
  inv_1 U4553 ( .ip(m2DataIn[6]), .op(n9467) );
  mux2_1 U4554 ( .ip1(n9216), .ip2(n9467), .s(n4293), .op(n4330) );
  mux2_1 U4555 ( .ip1(rdata[5]), .ip2(m2DataIn[5]), .s(n4293), .op(n4325) );
  mux2_1 U4556 ( .ip1(rdata[4]), .ip2(m2DataIn[4]), .s(n4293), .op(n4322) );
  inv_1 U4557 ( .ip(rdata[3]), .op(n8999) );
  inv_1 U4558 ( .ip(m2DataIn[3]), .op(n9530) );
  mux2_1 U4559 ( .ip1(n8999), .ip2(n9530), .s(n4293), .op(n4318) );
  mux2_1 U4560 ( .ip1(rdata[2]), .ip2(m2DataIn[2]), .s(n4293), .op(n4315) );
  inv_1 U4561 ( .ip(rdata[1]), .op(n8873) );
  inv_1 U4562 ( .ip(m2DataIn[1]), .op(n9417) );
  mux2_1 U4563 ( .ip1(n8873), .ip2(n9417), .s(n4293), .op(n4313) );
  inv_1 U4564 ( .ip(rdata[0]), .op(n8756) );
  inv_1 U4565 ( .ip(m2DataIn[0]), .op(n9335) );
  mux2_1 U4566 ( .ip1(n8756), .ip2(n9335), .s(n4293), .op(n4311) );
  nand2_1 U4567 ( .ip1(n4313), .ip2(n4311), .op(n4332) );
  nor2_1 U4568 ( .ip1(n4315), .ip2(n4332), .op(n4316) );
  nand2_1 U4569 ( .ip1(n4318), .ip2(n4316), .op(n4320) );
  or2_1 U4570 ( .ip1(n4322), .ip2(n4320), .op(n4323) );
  nor2_1 U4571 ( .ip1(n4325), .ip2(n4323), .op(n4327) );
  nand2_1 U4572 ( .ip1(n4330), .ip2(n4327), .op(n4308) );
  mux2_1 U4573 ( .ip1(rdata[7]), .ip2(m2DataIn[7]), .s(n4293), .op(n4310) );
  nor2_1 U4574 ( .ip1(n4308), .ip2(n4310), .op(n4284) );
  nor2_1 U4575 ( .ip1(n4328), .ip2(n4284), .op(n4283) );
  xor2_1 U4576 ( .ip1(n4285), .ip2(n4283), .op(n4358) );
  mux2_1 U4577 ( .ip1(rdata[9]), .ip2(m2DataIn[9]), .s(n4293), .op(n4295) );
  nand2_1 U4578 ( .ip1(n4285), .ip2(n4284), .op(n4294) );
  inv_1 U4579 ( .ip(n4294), .op(n8593) );
  nor2_1 U4580 ( .ip1(n4328), .ip2(n8593), .op(n4286) );
  xor2_1 U4581 ( .ip1(n4295), .ip2(n4286), .op(n4353) );
  inv_1 U4582 ( .ip(n4353), .op(n8592) );
  nand2_1 U4583 ( .ip1(n4358), .ip2(n8592), .op(n4363) );
  inv_1 U4584 ( .ip(n4363), .op(n4355) );
  inv_1 U4585 ( .ip(rdata[13]), .op(n9742) );
  inv_1 U4586 ( .ip(m2DataIn[13]), .op(n9799) );
  mux2_1 U4587 ( .ip1(n9742), .ip2(n9799), .s(n4293), .op(n4291) );
  inv_1 U4588 ( .ip(rdata[12]), .op(n9754) );
  inv_1 U4589 ( .ip(m2DataIn[12]), .op(n9815) );
  mux2_1 U4590 ( .ip1(n9754), .ip2(n9815), .s(n4293), .op(n4288) );
  nor2_1 U4591 ( .ip1(n4291), .ip2(n4288), .op(n4287) );
  nor2_1 U4592 ( .ip1(n4328), .ip2(n4287), .op(n4290) );
  mux2_1 U4593 ( .ip1(rdata[11]), .ip2(m2DataIn[11]), .s(n4293), .op(n4292) );
  nor2_1 U4594 ( .ip1(n4288), .ip2(n4292), .op(n4289) );
  nor2_1 U4595 ( .ip1(n4290), .ip2(n4289), .op(n4304) );
  inv_1 U4596 ( .ip(rdata[14]), .op(n9895) );
  inv_1 U4597 ( .ip(m2DataIn[14]), .op(n9863) );
  mux2_1 U4598 ( .ip1(n9895), .ip2(n9863), .s(n4293), .op(n4302) );
  inv_1 U4599 ( .ip(n4291), .op(n4301) );
  and2_1 U4600 ( .ip1(n4292), .ip2(n4328), .op(n4300) );
  inv_1 U4601 ( .ip(rdata[10]), .op(n9557) );
  inv_1 U4602 ( .ip(m2DataIn[10]), .op(n9792) );
  mux2_1 U4603 ( .ip1(n9557), .ip2(n9792), .s(n4293), .op(n4307) );
  or2_1 U4604 ( .ip1(n4307), .ip2(n4328), .op(n4297) );
  nor2_1 U4605 ( .ip1(n4295), .ip2(n4294), .op(n4305) );
  or2_1 U4606 ( .ip1(n4305), .ip2(n4328), .op(n4296) );
  nand2_1 U4607 ( .ip1(n4297), .ip2(n4296), .op(n4298) );
  nor2_1 U4608 ( .ip1(n4298), .ip2(n4302), .op(n4299) );
  not_ab_or_c_or_d U4609 ( .ip1(n4302), .ip2(n4301), .ip3(n4300), .ip4(n4299), 
        .op(n4303) );
  nand2_1 U4610 ( .ip1(n4304), .ip2(n4303), .op(n8594) );
  nor2_1 U4611 ( .ip1(n4328), .ip2(n4305), .op(n4306) );
  xor2_1 U4612 ( .ip1(n4307), .ip2(n4306), .op(n8591) );
  inv_1 U4613 ( .ip(n8591), .op(n4359) );
  nor2_1 U4614 ( .ip1(n8594), .ip2(n4359), .op(n4366) );
  nand2_1 U4615 ( .ip1(n4355), .ip2(n4366), .op(n4348) );
  nand2_1 U4616 ( .ip1(n4308), .ip2(\sig_in[15] ), .op(n4309) );
  xor2_1 U4617 ( .ip1(n4310), .ip2(n4309), .op(n8599) );
  inv_1 U4618 ( .ip(n8599), .op(n4391) );
  inv_1 U4619 ( .ip(n4311), .op(n4319) );
  nand2_1 U4620 ( .ip1(\sig_in[15] ), .ip2(n4319), .op(n4312) );
  xor2_1 U4621 ( .ip1(n4313), .ip2(n4312), .op(n4339) );
  and2_1 U4622 ( .ip1(\sig_in[15] ), .ip2(n4332), .op(n4314) );
  xor2_1 U4623 ( .ip1(n4315), .ip2(n4314), .op(n4338) );
  nor2_1 U4624 ( .ip1(n4328), .ip2(n4316), .op(n4317) );
  xor2_1 U4625 ( .ip1(n4318), .ip2(n4317), .op(n4340) );
  inv_1 U4626 ( .ip(n4340), .op(n4335) );
  not_ab_or_c_or_d U4627 ( .ip1(n4319), .ip2(n4339), .ip3(n4338), .ip4(n4335), 
        .op(n4326) );
  nand2_1 U4628 ( .ip1(n4320), .ip2(\sig_in[15] ), .op(n4321) );
  xor2_1 U4629 ( .ip1(n4322), .ip2(n4321), .op(n4341) );
  nand2_1 U4630 ( .ip1(n4323), .ip2(\sig_in[15] ), .op(n4324) );
  xor2_1 U4631 ( .ip1(n4325), .ip2(n4324), .op(n4344) );
  nor3_1 U4632 ( .ip1(n4326), .ip2(n4341), .ip3(n4344), .op(n4331) );
  nor2_1 U4633 ( .ip1(n4328), .ip2(n4327), .op(n4329) );
  xor2_1 U4634 ( .ip1(n4330), .ip2(n4329), .op(n4347) );
  inv_1 U4635 ( .ip(n4347), .op(n4350) );
  or2_1 U4636 ( .ip1(n4331), .ip2(n4350), .op(n4399) );
  nand2_1 U4637 ( .ip1(n4391), .ip2(n4399), .op(n8565) );
  inv_1 U4638 ( .ip(n8565), .op(n4367) );
  nand3_1 U4639 ( .ip1(n4332), .ip2(n4338), .ip3(n4335), .op(n4333) );
  nand3_1 U4640 ( .ip1(n4341), .ip2(n4344), .ip3(n4333), .op(n4334) );
  nand2_1 U4641 ( .ip1(n4350), .ip2(n4334), .op(n4400) );
  nand2_1 U4642 ( .ip1(n4367), .ip2(n4400), .op(n8617) );
  nor2_1 U4643 ( .ip1(n4348), .ip2(n8617), .op(n8633) );
  inv_1 U4644 ( .ip(n4341), .op(n4336) );
  not_ab_or_c_or_d U4645 ( .ip1(n4338), .ip2(n4339), .ip3(n4336), .ip4(n4335), 
        .op(n4337) );
  nor2_1 U4646 ( .ip1(n4344), .ip2(n4337), .op(n4351) );
  nor2_1 U4647 ( .ip1(n4351), .ip2(n4400), .op(n4349) );
  nand2_1 U4648 ( .ip1(n4349), .ip2(n4391), .op(n4373) );
  nor2_1 U4649 ( .ip1(n4348), .ip2(n4373), .op(n4384) );
  inv_1 U4650 ( .ip(n4366), .op(n8569) );
  nor3_1 U4651 ( .ip1(n4353), .ip2(n8569), .ip3(n4358), .op(n8635) );
  inv_1 U4652 ( .ip(n8635), .op(n8572) );
  inv_1 U4653 ( .ip(n4338), .op(n4343) );
  inv_1 U4654 ( .ip(n4339), .op(n4342) );
  not_ab_or_c_or_d U4655 ( .ip1(n4343), .ip2(n4342), .ip3(n4341), .ip4(n4340), 
        .op(n4346) );
  inv_1 U4656 ( .ip(n4344), .op(n4345) );
  nor2_1 U4657 ( .ip1(n4346), .ip2(n4345), .op(n4352) );
  nand2_1 U4658 ( .ip1(n4347), .ip2(n4352), .op(n8601) );
  inv_1 U4659 ( .ip(n8601), .op(n8582) );
  nand2_1 U4660 ( .ip1(n8599), .ip2(n8582), .op(n4386) );
  nor2_1 U4661 ( .ip1(n8572), .ip2(n4386), .op(n8632) );
  inv_1 U4662 ( .ip(n4348), .op(n8585) );
  nand2_1 U4663 ( .ip1(n8599), .ip2(n4349), .op(n4371) );
  inv_1 U4664 ( .ip(n4371), .op(n8581) );
  nand2_1 U4665 ( .ip1(n8585), .ip2(n8581), .op(n4402) );
  nand2_1 U4666 ( .ip1(n4351), .ip2(n4350), .op(n8564) );
  nor2_1 U4667 ( .ip1(n4391), .ip2(n8564), .op(n8571) );
  nand2_1 U4668 ( .ip1(n8585), .ip2(n8571), .op(n8598) );
  nand2_1 U4669 ( .ip1(n4402), .ip2(n8598), .op(n8628) );
  nor4_1 U4670 ( .ip1(n8633), .ip2(n4384), .ip3(n8632), .ip4(n8628), .op(n8597) );
  nor2_1 U4671 ( .ip1(n4352), .ip2(n4399), .op(n4398) );
  inv_1 U4672 ( .ip(n4398), .op(n8600) );
  nand3_1 U4673 ( .ip1(n4353), .ip2(n4358), .ip3(n4366), .op(n8616) );
  nor3_1 U4674 ( .ip1(n4391), .ip2(n8600), .ip3(n8616), .op(n4389) );
  nor2_1 U4675 ( .ip1(n4386), .ip2(n8616), .op(n4354) );
  not_ab_or_c_or_d U4676 ( .ip1(n8635), .ip2(n8581), .ip3(n4389), .ip4(n4354), 
        .op(n4380) );
  nor2_1 U4677 ( .ip1(n4373), .ip2(n8572), .op(n4378) );
  or2_1 U4678 ( .ip1(n4355), .ip2(n8591), .op(n4357) );
  inv_1 U4679 ( .ip(n4386), .op(n4392) );
  or2_1 U4680 ( .ip1(n4392), .ip2(n8591), .op(n4356) );
  nand2_1 U4681 ( .ip1(n4357), .ip2(n4356), .op(n4364) );
  nor2_1 U4682 ( .ip1(n8599), .ip2(n8564), .op(n4385) );
  or2_1 U4683 ( .ip1(n4385), .ip2(n4359), .op(n4361) );
  nor2_1 U4684 ( .ip1(n4358), .ip2(n8592), .op(n4365) );
  or2_1 U4685 ( .ip1(n4365), .ip2(n4359), .op(n4360) );
  nand2_1 U4686 ( .ip1(n4361), .ip2(n4360), .op(n4362) );
  or2_1 U4687 ( .ip1(n4364), .ip2(n4362), .op(n8586) );
  nor2_1 U4688 ( .ip1(n8586), .ip2(n8594), .op(n4370) );
  and2_1 U4689 ( .ip1(n4400), .ip2(n8599), .op(n8567) );
  nor2_1 U4690 ( .ip1(n8594), .ip2(n4363), .op(n8566) );
  and3_1 U4691 ( .ip1(n8567), .ip2(n8566), .ip3(n4364), .op(n4369) );
  nand2_1 U4692 ( .ip1(n4366), .ip2(n4365), .op(n4394) );
  inv_1 U4693 ( .ip(n4394), .op(n8576) );
  nand3_1 U4694 ( .ip1(n8564), .ip2(n8576), .ip3(n4367), .op(n4368) );
  nor2_1 U4695 ( .ip1(n8599), .ip2(n8600), .op(n4383) );
  nand2_1 U4696 ( .ip1(n4383), .ip2(n8576), .op(n8578) );
  nand2_1 U4697 ( .ip1(n4368), .ip2(n8578), .op(n8607) );
  nor3_1 U4698 ( .ip1(n4370), .ip2(n4369), .ip3(n8607), .op(n8640) );
  inv_1 U4699 ( .ip(n8640), .op(n4377) );
  inv_1 U4700 ( .ip(n8616), .op(n8583) );
  nor2_1 U4701 ( .ip1(n4371), .ip2(n8616), .op(n8614) );
  or2_1 U4702 ( .ip1(n8571), .ip2(n8614), .op(n4372) );
  nand2_1 U4703 ( .ip1(n8583), .ip2(n4372), .op(n8620) );
  inv_1 U4704 ( .ip(n8620), .op(n4376) );
  nor2_1 U4705 ( .ip1(n4373), .ip2(n8616), .op(n8604) );
  or2_1 U4706 ( .ip1(n4385), .ip2(n8604), .op(n4374) );
  nand2_1 U4707 ( .ip1(n4374), .ip2(n8583), .op(n8570) );
  nand2_1 U4708 ( .ip1(n4392), .ip2(n8576), .op(n4375) );
  nand2_1 U4709 ( .ip1(n8570), .ip2(n4375), .op(n4397) );
  nor4_1 U4710 ( .ip1(n4378), .ip2(n4377), .ip3(n4376), .ip4(n4397), .op(n4379) );
  nor2_1 U4711 ( .ip1(n8599), .ip2(n8601), .op(n8575) );
  nand2_1 U4712 ( .ip1(n8635), .ip2(n8575), .op(n4382) );
  nand4_1 U4713 ( .ip1(n8597), .ip2(n4380), .ip3(n4379), .ip4(n4382), .op(
        n3840) );
  nor2_1 U4714 ( .ip1(n8599), .ip2(n8572), .op(n8631) );
  nand2_1 U4715 ( .ip1(n4398), .ip2(n8631), .op(n4381) );
  nand2_1 U4716 ( .ip1(n4382), .ip2(n4381), .op(n8574) );
  inv_1 U4717 ( .ip(n8574), .op(n4404) );
  nand2_1 U4718 ( .ip1(n8585), .ip2(n4383), .op(n8579) );
  inv_1 U4719 ( .ip(n8579), .op(n8622) );
  not_ab_or_c_or_d U4720 ( .ip1(n8585), .ip2(n4385), .ip3(n4384), .ip4(n8622), 
        .op(n8637) );
  or2_1 U4721 ( .ip1(n4386), .ip2(n8616), .op(n4388) );
  nand2_1 U4722 ( .ip1(n4399), .ip2(n8567), .op(n4390) );
  or2_1 U4723 ( .ip1(n4390), .ip2(n8616), .op(n4387) );
  nand2_1 U4724 ( .ip1(n4388), .ip2(n4387), .op(n8608) );
  nor2_1 U4725 ( .ip1(n4389), .ip2(n8608), .op(n8621) );
  inv_1 U4726 ( .ip(n4390), .op(n8584) );
  nor3_1 U4727 ( .ip1(n4392), .ip2(n4399), .ip3(n4391), .op(n8634) );
  nor2_1 U4728 ( .ip1(n8584), .ip2(n8634), .op(n4393) );
  nor2_1 U4729 ( .ip1(n4394), .ip2(n4393), .op(n8613) );
  nor3_1 U4730 ( .ip1(n8575), .ip2(n8581), .ip3(n8571), .op(n4395) );
  nor2_1 U4731 ( .ip1(n4395), .ip2(n4394), .op(n4396) );
  nor3_1 U4732 ( .ip1(n4397), .ip2(n8613), .ip3(n4396), .op(n8639) );
  nand3_1 U4733 ( .ip1(n8585), .ip2(n8599), .ip3(n4398), .op(n8623) );
  nand3_1 U4734 ( .ip1(n8635), .ip2(n4400), .ip3(n4399), .op(n4401) );
  and4_1 U4735 ( .ip1(n8639), .ip2(n4402), .ip3(n8623), .ip4(n4401), .op(n4403) );
  nand4_1 U4736 ( .ip1(n4404), .ip2(n8637), .ip3(n8621), .ip4(n4403), .op(
        n3839) );
  nor2_1 U4737 ( .ip1(\CNTRL/currentState [2]), .ip2(n8195), .op(n8223) );
  nand2_1 U4738 ( .ip1(n8223), .ip2(n4405), .op(n10017) );
  nand3_1 U4739 ( .ip1(\CNTRL/currentState [1]), .ip2(n8223), .ip3(
        \CNTRL/count_20Q [0]), .op(n10018) );
  nand2_1 U4740 ( .ip1(n10017), .ip2(n10018), .op(n10053) );
  inv_1 U4741 ( .ip(\CNTRL/count_20Q [1]), .op(n8801) );
  inv_1 U4742 ( .ip(\CNTRL/currentState [2]), .op(n8807) );
  nor2_1 U4743 ( .ip1(n8810), .ip2(n8807), .op(n8804) );
  or2_1 U4744 ( .ip1(n4405), .ip2(n8804), .op(n4406) );
  nand2_1 U4745 ( .ip1(n8802), .ip2(n4406), .op(n8328) );
  nor2_1 U4746 ( .ip1(\CNTRL/count_20Q [2]), .ip2(\CNTRL/count_20Q [3]), .op(
        n8336) );
  nand3_1 U4747 ( .ip1(\CNTRL/count_20Q [4]), .ip2(n8328), .ip3(n8336), .op(
        n8314) );
  nor2_1 U4748 ( .ip1(n8801), .ip2(n8314), .op(n8523) );
  and2_1 U4749 ( .ip1(n10053), .ip2(n8523), .op(weight2_loadNextRow) );
  nand3_1 U4750 ( .ip1(\CNTRL/currentState [2]), .ip2(\CNTRL/currentState [0]), 
        .ip3(\CNTRL/currentState [1]), .op(n9445) );
  inv_1 U4751 ( .ip(n9445), .op(n9907) );
  nor4_1 U4752 ( .ip1(n8810), .ip2(reset), .ip3(n9907), .ip4(
        weight2_loadNextRow), .op(n4040) );
  inv_1 U4753 ( .ip(\STAGE_1/weightReg [1]), .op(n5535) );
  inv_1 U4754 ( .ip(n5535), .op(n6248) );
  inv_1 U4755 ( .ip(\STAGE_1/weightReg [3]), .op(n5500) );
  inv_1 U4756 ( .ip(n5500), .op(n8001) );
  nand2_1 U4757 ( .ip1(m1Inputs[146]), .ip2(\STAGE_1/weightReg [3]), .op(n4408) );
  inv_1 U4758 ( .ip(\STAGE_1/weightReg [0]), .op(n5552) );
  nand2_1 U4759 ( .ip1(m1Inputs[149]), .ip2(\STAGE_1/weightReg [0]), .op(n4407) );
  xor2_1 U4760 ( .ip1(n4408), .ip2(n4407), .op(n4466) );
  inv_1 U4761 ( .ip(\STAGE_1/weightReg [5]), .op(n7624) );
  nand3_1 U4762 ( .ip1(m1Inputs[144]), .ip2(n4466), .ip3(
        \STAGE_1/weightReg [5]), .op(n4410) );
  nand4_1 U4763 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n8001), .ip3(
        m1Inputs[146]), .ip4(m1Inputs[149]), .op(n4409) );
  nand2_1 U4764 ( .ip1(n4410), .ip2(n4409), .op(n4462) );
  buf_1 U4765 ( .ip(\STAGE_1/weightReg [2]), .op(n6280) );
  nand2_1 U4766 ( .ip1(n6280), .ip2(m1Inputs[148]), .op(n6282) );
  buf_1 U4767 ( .ip(n5535), .op(n5414) );
  inv_1 U4768 ( .ip(m1Inputs[149]), .op(n8060) );
  nor3_1 U4769 ( .ip1(n5414), .ip2(n6282), .ip3(n8060), .op(n4453) );
  or2_1 U4770 ( .ip1(n6282), .ip2(n4453), .op(n4413) );
  nand2_1 U4771 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[149]), .op(n4411) );
  or2_1 U4772 ( .ip1(n4411), .ip2(n4453), .op(n4412) );
  nand2_1 U4773 ( .ip1(n4413), .ip2(n4412), .op(n4461) );
  inv_1 U4774 ( .ip(m1Inputs[145]), .op(n4482) );
  inv_1 U4775 ( .ip(\STAGE_1/weightReg [5]), .op(n7813) );
  nor2_1 U4776 ( .ip1(n4482), .ip2(n7813), .op(n4436) );
  inv_1 U4777 ( .ip(\STAGE_1/weightReg [0]), .op(n5475) );
  inv_1 U4778 ( .ip(m1Inputs[150]), .op(n8046) );
  nor2_1 U4779 ( .ip1(n5475), .ip2(n8046), .op(n4435) );
  inv_1 U4780 ( .ip(m1Inputs[144]), .op(n4493) );
  inv_1 U4781 ( .ip(\STAGE_1/weightReg [6]), .op(n5669) );
  nor2_1 U4782 ( .ip1(n4493), .ip2(n5669), .op(n4434) );
  and3_1 U4783 ( .ip1(n6248), .ip2(m1Inputs[150]), .ip3(n4450), .op(n6275) );
  inv_1 U4784 ( .ip(m1Inputs[148]), .op(n8077) );
  nand2_1 U4785 ( .ip1(n8001), .ip2(m1Inputs[151]), .op(n8004) );
  nor3_1 U4786 ( .ip1(n5552), .ip2(n8077), .ip3(n8004), .op(n4430) );
  inv_1 U4787 ( .ip(\STAGE_1/weightReg [3]), .op(n6246) );
  nor2_1 U4788 ( .ip1(n6246), .ip2(n8077), .op(n4414) );
  or2_1 U4789 ( .ip1(m1Inputs[151]), .ip2(n4414), .op(n4416) );
  or2_1 U4790 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n4414), .op(n4415) );
  nand2_1 U4791 ( .ip1(n4416), .ip2(n4415), .op(n4429) );
  nand2_1 U4792 ( .ip1(n6280), .ip2(m1Inputs[149]), .op(n4431) );
  nor2_1 U4793 ( .ip1(n4429), .ip2(n4431), .op(n4417) );
  nor2_1 U4794 ( .ip1(n4430), .ip2(n4417), .op(n6265) );
  nand2_1 U4795 ( .ip1(\STAGE_1/weightReg [5]), .ip2(m1Inputs[146]), .op(n4419) );
  buf_1 U4796 ( .ip(\STAGE_1/weightReg [4]), .op(n8078) );
  nand2_1 U4797 ( .ip1(n8078), .ip2(m1Inputs[147]), .op(n4418) );
  xor2_1 U4798 ( .ip1(n4419), .ip2(n4418), .op(n4425) );
  inv_1 U4799 ( .ip(m1Inputs[147]), .op(n8000) );
  nand2_1 U4800 ( .ip1(m1Inputs[146]), .ip2(\STAGE_1/weightReg [4]), .op(n4464) );
  nor3_1 U4801 ( .ip1(n8000), .ip2(n7813), .ip3(n4464), .op(n4420) );
  or2_1 U4802 ( .ip1(n4425), .ip2(n4420), .op(n4422) );
  inv_1 U4803 ( .ip(\STAGE_1/weightReg [7]), .op(n7685) );
  nor2_1 U4804 ( .ip1(n4493), .ip2(n7685), .op(n4424) );
  or2_1 U4805 ( .ip1(n4424), .ip2(n4420), .op(n4421) );
  nand2_1 U4806 ( .ip1(n4422), .ip2(n4421), .op(n6264) );
  nand2_1 U4807 ( .ip1(m1Inputs[146]), .ip2(\STAGE_1/weightReg [6]), .op(n6263) );
  inv_1 U4808 ( .ip(n4423), .op(n6272) );
  xnor2_1 U4809 ( .ip1(n4425), .ip2(n4424), .op(n4447) );
  nand2_1 U4810 ( .ip1(n6248), .ip2(m1Inputs[147]), .op(n6294) );
  nor2_1 U4811 ( .ip1(n6282), .ip2(n6294), .op(n4459) );
  and2_1 U4812 ( .ip1(n8001), .ip2(n4459), .op(n4428) );
  nand2_1 U4813 ( .ip1(n8001), .ip2(m1Inputs[147]), .op(n4426) );
  mux2_1 U4814 ( .ip1(n4426), .ip2(n8001), .s(n4459), .op(n4463) );
  nor2_1 U4815 ( .ip1(n4464), .ip2(n4463), .op(n4427) );
  nor2_1 U4816 ( .ip1(n4428), .ip2(n4427), .op(n4446) );
  nor2_1 U4817 ( .ip1(n4430), .ip2(n4429), .op(n4432) );
  xor2_1 U4818 ( .ip1(n4432), .ip2(n4431), .op(n4445) );
  inv_1 U4819 ( .ip(n4433), .op(n6271) );
  nor2_1 U4820 ( .ip1(n4482), .ip2(n5669), .op(n4454) );
  fulladder U4821 ( .a(n4436), .b(n4435), .ci(n4434), .co(n4452), .s(n4460) );
  nor2_1 U4822 ( .ip1(n5060), .ip2(n8060), .op(n6298) );
  and3_1 U4823 ( .ip1(n8001), .ip2(m1Inputs[148]), .ip3(n6298), .op(n6242) );
  nor2_1 U4824 ( .ip1(n6246), .ip2(n8060), .op(n4437) );
  or2_1 U4825 ( .ip1(m1Inputs[148]), .ip2(n4437), .op(n4439) );
  or2_1 U4826 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n4437), .op(n4438) );
  nand2_1 U4827 ( .ip1(n4439), .ip2(n4438), .op(n4440) );
  nor2_1 U4828 ( .ip1(n6242), .ip2(n4440), .op(n6241) );
  nor2_1 U4829 ( .ip1(n4482), .ip2(n7685), .op(n6243) );
  xor2_1 U4830 ( .ip1(n6241), .ip2(n6243), .op(n6262) );
  nor2_1 U4831 ( .ip1(n8000), .ip2(n7813), .op(n6257) );
  inv_1 U4832 ( .ip(m1Inputs[152]), .op(n8030) );
  nor2_1 U4833 ( .ip1(n5552), .ip2(n8030), .op(n6256) );
  nand2_1 U4834 ( .ip1(m1Inputs[144]), .ip2(\STAGE_1/weightReg [15]), .op(
        n6255) );
  inv_1 U4835 ( .ip(m1Inputs[151]), .op(n8031) );
  nor2_1 U4836 ( .ip1(n5535), .ip2(n8031), .op(n6259) );
  nor2_1 U4837 ( .ip1(\CNTRL/count_layer1_784Q [0]), .ip2(
        \CNTRL/count_layer1_784Q [1]), .op(n8198) );
  nor4_1 U4838 ( .ip1(\CNTRL/count_layer1_784Q [2]), .ip2(
        \CNTRL/count_layer1_784Q [3]), .ip3(\CNTRL/count_layer1_784Q [8]), 
        .ip4(\CNTRL/count_layer1_784Q [9]), .op(n4443) );
  or4_1 U4839 ( .ip1(\CNTRL/currentState [2]), .ip2(
        \CNTRL/count_layer1_784Q [6]), .ip3(\CNTRL/count_layer1_784Q [7]), 
        .ip4(\CNTRL/count_layer1_784Q [5]), .op(n4441) );
  nor3_1 U4840 ( .ip1(\CNTRL/count_layer1_784Q [4]), .ip2(n4442), .ip3(n4441), 
        .op(n8187) );
  nand3_1 U4841 ( .ip1(n8198), .ip2(n4443), .ip3(n8187), .op(n4444) );
  nand2_1 U4842 ( .ip1(n4444), .ip2(n10017), .op(n8180) );
  inv_1 U4843 ( .ip(n8180), .op(n8175) );
  nand2_1 U4844 ( .ip1(n8175), .ip2(column[144]), .op(n6267) );
  inv_1 U4845 ( .ip(\STAGE_1/weightReg [2]), .op(n5593) );
  nor2_1 U4846 ( .ip1(n5593), .ip2(n8046), .op(n6258) );
  fulladder U4847 ( .a(n4447), .b(n4446), .ci(n4445), .co(n4433), .s(n4448) );
  inv_1 U4848 ( .ip(n4448), .op(n4529) );
  nor2_1 U4849 ( .ip1(n5535), .ip2(n8046), .op(n4449) );
  nor2_1 U4850 ( .ip1(n4450), .ip2(n4449), .op(n4451) );
  nor2_1 U4851 ( .ip1(n6275), .ip2(n4451), .op(n4528) );
  fulladder U4852 ( .a(n4454), .b(n4453), .ci(n4452), .co(n6270), .s(n4527) );
  nand2_1 U4853 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[146]), .op(n4492) );
  nor3_1 U4854 ( .ip1(n5593), .ip2(n8000), .ip3(n4492), .op(n4473) );
  nor2_1 U4855 ( .ip1(n5593), .ip2(n8000), .op(n4455) );
  or2_1 U4856 ( .ip1(m1Inputs[148]), .ip2(n4455), .op(n4457) );
  or2_1 U4857 ( .ip1(\STAGE_1/weightReg [1]), .ip2(n4455), .op(n4456) );
  nand2_1 U4858 ( .ip1(n4457), .ip2(n4456), .op(n4458) );
  nor2_1 U4859 ( .ip1(n4459), .ip2(n4458), .op(n4468) );
  nor2_1 U4860 ( .ip1(n4482), .ip2(n5060), .op(n4467) );
  fulladder U4861 ( .a(n4462), .b(n4461), .ci(n4460), .co(n4450), .s(n4471) );
  xor2_1 U4862 ( .ip1(n4464), .ip2(n4463), .op(n4470) );
  nand2_1 U4863 ( .ip1(n4518), .ip2(n4517), .op(n4526) );
  nor2_1 U4864 ( .ip1(n4493), .ip2(n7813), .op(n4465) );
  xor2_1 U4865 ( .ip1(n4466), .ip2(n4465), .op(n4510) );
  fulladder U4866 ( .a(n4473), .b(n4468), .ci(n4467), .co(n4472), .s(n4509) );
  nor2_1 U4867 ( .ip1(n5552), .ip2(n8077), .op(n4479) );
  nor2_1 U4868 ( .ip1(n6246), .ip2(n4482), .op(n4478) );
  nor2_1 U4869 ( .ip1(n4493), .ip2(n5060), .op(n4477) );
  inv_1 U4870 ( .ip(n4469), .op(n4524) );
  fulladder U4871 ( .a(n4472), .b(n4471), .ci(n4470), .co(n4517), .s(n4520) );
  nor3_1 U4872 ( .ip1(n6246), .ip2(n4493), .ip3(n4492), .op(n4497) );
  or2_1 U4873 ( .ip1(n6294), .ip2(n4473), .op(n4476) );
  nand2_1 U4874 ( .ip1(n6280), .ip2(m1Inputs[146]), .op(n4474) );
  or2_1 U4875 ( .ip1(n4474), .ip2(n4473), .op(n4475) );
  nand2_1 U4876 ( .ip1(n4476), .ip2(n4475), .op(n4481) );
  fulladder U4877 ( .a(n4479), .b(n4478), .ci(n4477), .co(n4508), .s(n4480) );
  fulladder U4878 ( .a(n4497), .b(n4481), .ci(n4480), .co(n4511), .s(n4502) );
  nand4_1 U4879 ( .ip1(\STAGE_1/weightReg [1]), .ip2(\STAGE_1/weightReg [2]), 
        .ip3(m1Inputs[145]), .ip4(m1Inputs[144]), .op(n4484) );
  not_ab_or_c_or_d U4880 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[144]), 
        .ip3(n5593), .ip4(n4482), .op(n4491) );
  nand3_1 U4881 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n4491), .ip3(
        m1Inputs[147]), .op(n4483) );
  nand2_1 U4882 ( .ip1(n4484), .ip2(n4483), .op(n4504) );
  nand2_1 U4883 ( .ip1(n4502), .ip2(n4504), .op(n4507) );
  inv_1 U4884 ( .ip(\STAGE_1/weightReg [2]), .op(n5175) );
  nand2_1 U4885 ( .ip1(m1Inputs[144]), .ip2(n5175), .op(n4485) );
  inv_1 U4886 ( .ip(m1Inputs[146]), .op(n6279) );
  nand2_1 U4887 ( .ip1(n4485), .ip2(n6279), .op(n4489) );
  nand2_1 U4888 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[145]), .op(n4487) );
  nand2_1 U4889 ( .ip1(n6280), .ip2(m1Inputs[144]), .op(n4486) );
  nand2_1 U4890 ( .ip1(n4487), .ip2(n4486), .op(n4488) );
  nand3_1 U4891 ( .ip1(n4489), .ip2(\STAGE_1/weightReg [0]), .ip3(n4488), .op(
        n4498) );
  nand2_1 U4892 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[147]), .op(n4490) );
  xor2_1 U4893 ( .ip1(n4491), .ip2(n4490), .op(n4499) );
  nor2_1 U4894 ( .ip1(n4498), .ip2(n4499), .op(n4501) );
  inv_1 U4895 ( .ip(n4492), .op(n4495) );
  nor2_1 U4896 ( .ip1(n6246), .ip2(n4493), .op(n4494) );
  nor2_1 U4897 ( .ip1(n4495), .ip2(n4494), .op(n4496) );
  not_ab_or_c_or_d U4898 ( .ip1(n4499), .ip2(n4498), .ip3(n4497), .ip4(n4496), 
        .op(n4500) );
  or2_1 U4899 ( .ip1(n4501), .ip2(n4500), .op(n4503) );
  nand2_1 U4900 ( .ip1(n4502), .ip2(n4503), .op(n4506) );
  nand2_1 U4901 ( .ip1(n4504), .ip2(n4503), .op(n4505) );
  nand3_1 U4902 ( .ip1(n4507), .ip2(n4506), .ip3(n4505), .op(n4513) );
  nand2_1 U4903 ( .ip1(n4511), .ip2(n4513), .op(n4516) );
  fulladder U4904 ( .a(n4510), .b(n4509), .ci(n4508), .co(n4469), .s(n4512) );
  nand2_1 U4905 ( .ip1(n4511), .ip2(n4512), .op(n4515) );
  nand2_1 U4906 ( .ip1(n4513), .ip2(n4512), .op(n4514) );
  nand3_1 U4907 ( .ip1(n4516), .ip2(n4515), .ip3(n4514), .op(n4519) );
  nand2_1 U4908 ( .ip1(n4520), .ip2(n4519), .op(n4523) );
  nor2_1 U4909 ( .ip1(n4518), .ip2(n4517), .op(n4522) );
  nor2_1 U4910 ( .ip1(n4520), .ip2(n4519), .op(n4521) );
  ab_or_c_or_d U4911 ( .ip1(n4524), .ip2(n4523), .ip3(n4522), .ip4(n4521), 
        .op(n4525) );
  nand2_1 U4912 ( .ip1(n4526), .ip2(n4525), .op(n6277) );
  fulladder U4913 ( .a(n4529), .b(n4528), .ci(n4527), .co(n6276), .s(n4518) );
  inv_1 U4914 ( .ip(m1Inputs[133]), .op(n7865) );
  nor2_1 U4915 ( .ip1(n5475), .ip2(n7865), .op(n4580) );
  inv_1 U4916 ( .ip(m1Inputs[130]), .op(n6221) );
  nor2_1 U4917 ( .ip1(n6246), .ip2(n6221), .op(n4579) );
  inv_1 U4918 ( .ip(m1Inputs[128]), .op(n4611) );
  nor2_1 U4919 ( .ip1(n4611), .ip2(n7813), .op(n4578) );
  nand2_1 U4920 ( .ip1(n6280), .ip2(m1Inputs[132]), .op(n6223) );
  nor3_1 U4921 ( .ip1(n5414), .ip2(n6223), .ip3(n7865), .op(n4566) );
  or2_1 U4922 ( .ip1(n6223), .ip2(n4566), .op(n4532) );
  nand2_1 U4923 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[133]), .op(n4530) );
  or2_1 U4924 ( .ip1(n4530), .ip2(n4566), .op(n4531) );
  nand2_1 U4925 ( .ip1(n4532), .ip2(n4531), .op(n4574) );
  inv_1 U4926 ( .ip(m1Inputs[129]), .op(n4610) );
  nor2_1 U4927 ( .ip1(n4610), .ip2(n7813), .op(n4555) );
  inv_1 U4928 ( .ip(m1Inputs[134]), .op(n7849) );
  nor2_1 U4929 ( .ip1(n5475), .ip2(n7849), .op(n4554) );
  nor2_1 U4930 ( .ip1(n4611), .ip2(n5669), .op(n4553) );
  and3_1 U4931 ( .ip1(n6248), .ip2(m1Inputs[134]), .ip3(n4563), .op(n6202) );
  inv_1 U4932 ( .ip(m1Inputs[132]), .op(n7881) );
  nand2_1 U4933 ( .ip1(n8001), .ip2(m1Inputs[135]), .op(n7819) );
  nor3_1 U4934 ( .ip1(n5475), .ip2(n7881), .ip3(n7819), .op(n4549) );
  nor2_1 U4935 ( .ip1(n6246), .ip2(n7881), .op(n4533) );
  or2_1 U4936 ( .ip1(m1Inputs[135]), .ip2(n4533), .op(n4535) );
  or2_1 U4937 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n4533), .op(n4534) );
  nand2_1 U4938 ( .ip1(n4535), .ip2(n4534), .op(n4548) );
  nand2_1 U4939 ( .ip1(n6280), .ip2(m1Inputs[133]), .op(n4550) );
  nor2_1 U4940 ( .ip1(n4548), .ip2(n4550), .op(n4536) );
  nor2_1 U4941 ( .ip1(n4549), .ip2(n4536), .op(n6192) );
  nand2_1 U4942 ( .ip1(n8078), .ip2(m1Inputs[131]), .op(n4538) );
  nand2_1 U4943 ( .ip1(\STAGE_1/weightReg [5]), .ip2(m1Inputs[130]), .op(n4537) );
  xor2_1 U4944 ( .ip1(n4538), .ip2(n4537), .op(n4544) );
  inv_1 U4945 ( .ip(m1Inputs[131]), .op(n7820) );
  nand2_1 U4946 ( .ip1(m1Inputs[130]), .ip2(\STAGE_1/weightReg [4]), .op(n4577) );
  nor3_1 U4947 ( .ip1(n7820), .ip2(n7624), .ip3(n4577), .op(n4539) );
  or2_1 U4948 ( .ip1(n4544), .ip2(n4539), .op(n4541) );
  nor2_1 U4949 ( .ip1(n4611), .ip2(n7685), .op(n4543) );
  or2_1 U4950 ( .ip1(n4543), .ip2(n4539), .op(n4540) );
  nand2_1 U4951 ( .ip1(n4541), .ip2(n4540), .op(n6191) );
  nand2_1 U4952 ( .ip1(m1Inputs[130]), .ip2(\STAGE_1/weightReg [6]), .op(n6190) );
  inv_1 U4953 ( .ip(n4542), .op(n6199) );
  xnor2_1 U4954 ( .ip1(n4544), .ip2(n4543), .op(n4560) );
  nor3_1 U4955 ( .ip1(n5414), .ip2(n7820), .ip3(n6223), .op(n4572) );
  and2_1 U4956 ( .ip1(n8001), .ip2(n4572), .op(n4547) );
  nand2_1 U4957 ( .ip1(n8001), .ip2(m1Inputs[131]), .op(n4545) );
  mux2_1 U4958 ( .ip1(n4545), .ip2(n8001), .s(n4572), .op(n4576) );
  nor2_1 U4959 ( .ip1(n4577), .ip2(n4576), .op(n4546) );
  nor2_1 U4960 ( .ip1(n4547), .ip2(n4546), .op(n4559) );
  nor2_1 U4961 ( .ip1(n4549), .ip2(n4548), .op(n4551) );
  xor2_1 U4962 ( .ip1(n4551), .ip2(n4550), .op(n4558) );
  inv_1 U4963 ( .ip(n4552), .op(n6198) );
  nor2_1 U4964 ( .ip1(n4610), .ip2(n5669), .op(n4567) );
  fulladder U4965 ( .a(n4555), .b(n4554), .ci(n4553), .co(n4565), .s(n4573) );
  nand2_1 U4966 ( .ip1(m1Inputs[132]), .ip2(\STAGE_1/weightReg [4]), .op(n4557) );
  nand2_1 U4967 ( .ip1(m1Inputs[133]), .ip2(\STAGE_1/weightReg [3]), .op(n4556) );
  xor2_1 U4968 ( .ip1(n4557), .ip2(n4556), .op(n6170) );
  nor2_1 U4969 ( .ip1(n4610), .ip2(n7685), .op(n6172) );
  xor2_1 U4970 ( .ip1(n6170), .ip2(n6172), .op(n6189) );
  nor2_1 U4971 ( .ip1(n7820), .ip2(n7624), .op(n6184) );
  inv_1 U4972 ( .ip(m1Inputs[136]), .op(n7840) );
  nor2_1 U4973 ( .ip1(n5475), .ip2(n7840), .op(n6183) );
  nand2_1 U4974 ( .ip1(m1Inputs[128]), .ip2(\STAGE_1/weightReg [15]), .op(
        n6182) );
  inv_1 U4975 ( .ip(m1Inputs[135]), .op(n7841) );
  nor2_1 U4976 ( .ip1(n5414), .ip2(n7841), .op(n6186) );
  nand2_1 U4977 ( .ip1(n8175), .ip2(column[128]), .op(n6194) );
  nor2_1 U4978 ( .ip1(n5593), .ip2(n7849), .op(n6185) );
  fulladder U4979 ( .a(n4560), .b(n4559), .ci(n4558), .co(n4552), .s(n4561) );
  inv_1 U4980 ( .ip(n4561), .op(n4643) );
  nor2_1 U4981 ( .ip1(n5535), .ip2(n7849), .op(n4562) );
  nor2_1 U4982 ( .ip1(n4563), .ip2(n4562), .op(n4564) );
  nor2_1 U4983 ( .ip1(n6202), .ip2(n4564), .op(n4642) );
  fulladder U4984 ( .a(n4567), .b(n4566), .ci(n4565), .co(n6197), .s(n4641) );
  nand2_1 U4985 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[130]), .op(n4599) );
  nor3_1 U4986 ( .ip1(n5593), .ip2(n4599), .ip3(n7820), .op(n4587) );
  nor2_1 U4987 ( .ip1(n5593), .ip2(n7820), .op(n4568) );
  or2_1 U4988 ( .ip1(m1Inputs[132]), .ip2(n4568), .op(n4570) );
  or2_1 U4989 ( .ip1(\STAGE_1/weightReg [1]), .ip2(n4568), .op(n4569) );
  nand2_1 U4990 ( .ip1(n4570), .ip2(n4569), .op(n4571) );
  nor2_1 U4991 ( .ip1(n4572), .ip2(n4571), .op(n4582) );
  nor2_1 U4992 ( .ip1(n4610), .ip2(n5060), .op(n4581) );
  fulladder U4993 ( .a(n4575), .b(n4574), .ci(n4573), .co(n4563), .s(n4629) );
  xor2_1 U4994 ( .ip1(n4577), .ip2(n4576), .op(n4628) );
  and2_1 U4995 ( .ip1(n4638), .ip2(n4637), .op(n4632) );
  fulladder U4996 ( .a(n4580), .b(n4579), .ci(n4578), .co(n4575), .s(n4621) );
  fulladder U4997 ( .a(n4587), .b(n4582), .ci(n4581), .co(n4630), .s(n4620) );
  nor2_1 U4998 ( .ip1(n5475), .ip2(n7881), .op(n4590) );
  nor2_1 U4999 ( .ip1(n4611), .ip2(n5060), .op(n4589) );
  nor2_1 U5000 ( .ip1(n6246), .ip2(n4610), .op(n4588) );
  nor3_1 U5001 ( .ip1(n6246), .ip2(n4611), .ip3(n4599), .op(n4600) );
  nor2_1 U5002 ( .ip1(n5414), .ip2(n7820), .op(n4583) );
  or2_1 U5003 ( .ip1(m1Inputs[130]), .ip2(n4583), .op(n4585) );
  or2_1 U5004 ( .ip1(\STAGE_1/weightReg [2]), .ip2(n4583), .op(n4584) );
  nand2_1 U5005 ( .ip1(n4585), .ip2(n4584), .op(n4586) );
  nor2_1 U5006 ( .ip1(n4587), .ip2(n4586), .op(n4592) );
  fulladder U5007 ( .a(n4590), .b(n4589), .ci(n4588), .co(n4619), .s(n4591) );
  fulladder U5008 ( .a(n4600), .b(n4592), .ci(n4591), .co(n4622), .s(n4615) );
  nand2_1 U5009 ( .ip1(n6280), .ip2(m1Inputs[128]), .op(n4597) );
  nand2_1 U5010 ( .ip1(n6248), .ip2(m1Inputs[129]), .op(n4596) );
  or2_1 U5011 ( .ip1(m1Inputs[128]), .ip2(m1Inputs[130]), .op(n4594) );
  or2_1 U5012 ( .ip1(n5593), .ip2(m1Inputs[130]), .op(n4593) );
  nand2_1 U5013 ( .ip1(n4594), .ip2(n4593), .op(n4595) );
  not_ab_or_c_or_d U5014 ( .ip1(n4597), .ip2(n4596), .ip3(n4595), .ip4(n5552), 
        .op(n4604) );
  not_ab_or_c_or_d U5015 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[128]), 
        .ip3(n5593), .ip4(n4610), .op(n4612) );
  nor2_1 U5016 ( .ip1(n5552), .ip2(n7820), .op(n4598) );
  xor2_1 U5017 ( .ip1(n4612), .ip2(n4598), .op(n4606) );
  nand2_1 U5018 ( .ip1(n4604), .ip2(n4606), .op(n4609) );
  or2_1 U5019 ( .ip1(n4599), .ip2(n4600), .op(n4603) );
  nand2_1 U5020 ( .ip1(n8001), .ip2(m1Inputs[128]), .op(n4601) );
  or2_1 U5021 ( .ip1(n4601), .ip2(n4600), .op(n4602) );
  nand2_1 U5022 ( .ip1(n4603), .ip2(n4602), .op(n4605) );
  nand2_1 U5023 ( .ip1(n4604), .ip2(n4605), .op(n4608) );
  nand2_1 U5024 ( .ip1(n4606), .ip2(n4605), .op(n4607) );
  nand3_1 U5025 ( .ip1(n4609), .ip2(n4608), .ip3(n4607), .op(n4616) );
  nor2_1 U5026 ( .ip1(n4615), .ip2(n4616), .op(n4618) );
  nor4_1 U5027 ( .ip1(n5414), .ip2(n5175), .ip3(n4611), .ip4(n4610), .op(n4614) );
  and3_1 U5028 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n4612), .ip3(m1Inputs[131]), .op(n4613) );
  not_ab_or_c_or_d U5029 ( .ip1(n4616), .ip2(n4615), .ip3(n4614), .ip4(n4613), 
        .op(n4617) );
  nor2_1 U5030 ( .ip1(n4618), .ip2(n4617), .op(n4624) );
  nand2_1 U5031 ( .ip1(n4622), .ip2(n4624), .op(n4627) );
  fulladder U5032 ( .a(n4621), .b(n4620), .ci(n4619), .co(n4633), .s(n4623) );
  nand2_1 U5033 ( .ip1(n4622), .ip2(n4623), .op(n4626) );
  nand2_1 U5034 ( .ip1(n4624), .ip2(n4623), .op(n4625) );
  nand3_1 U5035 ( .ip1(n4627), .ip2(n4626), .ip3(n4625), .op(n4634) );
  nor3_1 U5036 ( .ip1(n4632), .ip2(n4633), .ip3(n4634), .op(n4636) );
  fulladder U5037 ( .a(n4630), .b(n4629), .ci(n4628), .co(n4637), .s(n4631) );
  not_ab_or_c_or_d U5038 ( .ip1(n4634), .ip2(n4633), .ip3(n4632), .ip4(n4631), 
        .op(n4635) );
  or2_1 U5039 ( .ip1(n4636), .ip2(n4635), .op(n4640) );
  nor2_1 U5040 ( .ip1(n4638), .ip2(n4637), .op(n4639) );
  nor2_1 U5041 ( .ip1(n4640), .ip2(n4639), .op(n6204) );
  fulladder U5042 ( .a(n4643), .b(n4642), .ci(n4641), .co(n6203), .s(n4638) );
  nand2_1 U5043 ( .ip1(m1Inputs[114]), .ip2(\STAGE_1/weightReg [3]), .op(n4645) );
  nand2_1 U5044 ( .ip1(m1Inputs[117]), .ip2(\STAGE_1/weightReg [0]), .op(n4644) );
  xor2_1 U5045 ( .ip1(n4645), .ip2(n4644), .op(n4700) );
  nand3_1 U5046 ( .ip1(m1Inputs[112]), .ip2(n4700), .ip3(n8064), .op(n4647) );
  nand4_1 U5047 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n8001), .ip3(
        m1Inputs[114]), .ip4(m1Inputs[117]), .op(n4646) );
  nand2_1 U5048 ( .ip1(n4647), .ip2(n4646), .op(n4696) );
  nand2_1 U5049 ( .ip1(n6280), .ip2(m1Inputs[116]), .op(n6152) );
  inv_1 U5050 ( .ip(m1Inputs[117]), .op(n7684) );
  nor3_1 U5051 ( .ip1(n5414), .ip2(n6152), .ip3(n7684), .op(n4687) );
  or2_1 U5052 ( .ip1(n6152), .ip2(n4687), .op(n4650) );
  nand2_1 U5053 ( .ip1(n6248), .ip2(m1Inputs[117]), .op(n4648) );
  or2_1 U5054 ( .ip1(n4648), .ip2(n4687), .op(n4649) );
  nand2_1 U5055 ( .ip1(n4650), .ip2(n4649), .op(n4695) );
  inv_1 U5056 ( .ip(m1Inputs[113]), .op(n4719) );
  nor2_1 U5057 ( .ip1(n4719), .ip2(n7624), .op(n4674) );
  inv_1 U5058 ( .ip(m1Inputs[118]), .op(n7663) );
  nor2_1 U5059 ( .ip1(n5475), .ip2(n7663), .op(n4673) );
  inv_1 U5060 ( .ip(m1Inputs[112]), .op(n4718) );
  nor2_1 U5061 ( .ip1(n4718), .ip2(n5669), .op(n4672) );
  and3_1 U5062 ( .ip1(n6248), .ip2(m1Inputs[118]), .ip3(n4684), .op(n6130) );
  inv_1 U5063 ( .ip(m1Inputs[116]), .op(n6107) );
  nand2_1 U5064 ( .ip1(n8001), .ip2(m1Inputs[119]), .op(n7631) );
  nor3_1 U5065 ( .ip1(n5552), .ip2(n6107), .ip3(n7631), .op(n4668) );
  nor2_1 U5066 ( .ip1(n6246), .ip2(n6107), .op(n4651) );
  or2_1 U5067 ( .ip1(m1Inputs[119]), .ip2(n4651), .op(n4653) );
  or2_1 U5068 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n4651), .op(n4652) );
  nand2_1 U5069 ( .ip1(n4653), .ip2(n4652), .op(n4667) );
  nand2_1 U5070 ( .ip1(n6280), .ip2(m1Inputs[117]), .op(n4669) );
  nor2_1 U5071 ( .ip1(n4667), .ip2(n4669), .op(n4654) );
  nor2_1 U5072 ( .ip1(n4668), .ip2(n4654), .op(n6120) );
  inv_1 U5073 ( .ip(n7813), .op(n8064) );
  nand2_1 U5074 ( .ip1(n8064), .ip2(m1Inputs[114]), .op(n4656) );
  nand2_1 U5075 ( .ip1(n8078), .ip2(m1Inputs[115]), .op(n4655) );
  xor2_1 U5076 ( .ip1(n4656), .ip2(n4655), .op(n4662) );
  inv_1 U5077 ( .ip(m1Inputs[114]), .op(n6150) );
  inv_1 U5078 ( .ip(\STAGE_1/weightReg [4]), .op(n5060) );
  nor2_1 U5079 ( .ip1(n6150), .ip2(n5060), .op(n4698) );
  inv_1 U5080 ( .ip(m1Inputs[115]), .op(n7629) );
  nor2_1 U5081 ( .ip1(n7629), .ip2(n7624), .op(n6112) );
  and2_1 U5082 ( .ip1(n4698), .ip2(n6112), .op(n4657) );
  or2_1 U5083 ( .ip1(n4662), .ip2(n4657), .op(n4659) );
  nor2_1 U5084 ( .ip1(n4718), .ip2(n7685), .op(n4661) );
  or2_1 U5085 ( .ip1(n4661), .ip2(n4657), .op(n4658) );
  nand2_1 U5086 ( .ip1(n4659), .ip2(n4658), .op(n6119) );
  nand2_1 U5087 ( .ip1(m1Inputs[114]), .ip2(\STAGE_1/weightReg [6]), .op(n6118) );
  inv_1 U5088 ( .ip(n4660), .op(n6127) );
  xnor2_1 U5089 ( .ip1(n4662), .ip2(n4661), .op(n4681) );
  nor3_1 U5090 ( .ip1(n5414), .ip2(n7629), .ip3(n6152), .op(n4693) );
  and2_1 U5091 ( .ip1(\STAGE_1/weightReg [3]), .ip2(n4693), .op(n4664) );
  or2_1 U5092 ( .ip1(n4698), .ip2(n4664), .op(n4666) );
  nor2_1 U5093 ( .ip1(n4693), .ip2(n7629), .op(n4663) );
  mux2_1 U5094 ( .ip1(n4663), .ip2(n4693), .s(n5500), .op(n4697) );
  or2_1 U5095 ( .ip1(n4697), .ip2(n4664), .op(n4665) );
  nand2_1 U5096 ( .ip1(n4666), .ip2(n4665), .op(n4680) );
  nor2_1 U5097 ( .ip1(n4668), .ip2(n4667), .op(n4670) );
  xor2_1 U5098 ( .ip1(n4670), .ip2(n4669), .op(n4679) );
  inv_1 U5099 ( .ip(n4671), .op(n6126) );
  nor2_1 U5100 ( .ip1(n4719), .ip2(n5669), .op(n4688) );
  fulladder U5101 ( .a(n4674), .b(n4673), .ci(n4672), .co(n4686), .s(n4694) );
  inv_1 U5102 ( .ip(m1Inputs[120]), .op(n7683) );
  nor2_1 U5103 ( .ip1(n5552), .ip2(n7683), .op(n6111) );
  nand2_1 U5104 ( .ip1(m1Inputs[112]), .ip2(\STAGE_1/weightReg [15]), .op(
        n6110) );
  nor2_1 U5105 ( .ip1(n5060), .ip2(n7684), .op(n6142) );
  and3_1 U5106 ( .ip1(n8001), .ip2(m1Inputs[116]), .ip3(n6142), .op(n6098) );
  nor2_1 U5107 ( .ip1(n6246), .ip2(n7684), .op(n4675) );
  or2_1 U5108 ( .ip1(m1Inputs[116]), .ip2(n4675), .op(n4677) );
  or2_1 U5109 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n4675), .op(n4676) );
  nand2_1 U5110 ( .ip1(n4677), .ip2(n4676), .op(n4678) );
  nor2_1 U5111 ( .ip1(n6098), .ip2(n4678), .op(n6097) );
  nor2_1 U5112 ( .ip1(n4719), .ip2(n7685), .op(n6099) );
  xor2_1 U5113 ( .ip1(n6097), .ip2(n6099), .op(n6116) );
  inv_1 U5114 ( .ip(m1Inputs[119]), .op(n7652) );
  nor2_1 U5115 ( .ip1(n5414), .ip2(n7652), .op(n6114) );
  buf_1 U5116 ( .ip(n8175), .op(n8009) );
  nand2_1 U5117 ( .ip1(n8009), .ip2(column[112]), .op(n6122) );
  nor2_1 U5118 ( .ip1(n5593), .ip2(n7663), .op(n6113) );
  fulladder U5119 ( .a(n4681), .b(n4680), .ci(n4679), .co(n4671), .s(n4682) );
  inv_1 U5120 ( .ip(n4682), .op(n4767) );
  nor2_1 U5121 ( .ip1(n5414), .ip2(n7663), .op(n4683) );
  nor2_1 U5122 ( .ip1(n4684), .ip2(n4683), .op(n4685) );
  nor2_1 U5123 ( .ip1(n6130), .ip2(n4685), .op(n4766) );
  fulladder U5124 ( .a(n4688), .b(n4687), .ci(n4686), .co(n6125), .s(n4765) );
  nand2_1 U5125 ( .ip1(n6248), .ip2(m1Inputs[114]), .op(n4721) );
  nor3_1 U5126 ( .ip1(n5593), .ip2(n7629), .ip3(n4721), .op(n4705) );
  nor2_1 U5127 ( .ip1(n5593), .ip2(n7629), .op(n4689) );
  or2_1 U5128 ( .ip1(m1Inputs[116]), .ip2(n4689), .op(n4691) );
  or2_1 U5129 ( .ip1(\STAGE_1/weightReg [1]), .ip2(n4689), .op(n4690) );
  nand2_1 U5130 ( .ip1(n4691), .ip2(n4690), .op(n4692) );
  nor2_1 U5131 ( .ip1(n4693), .ip2(n4692), .op(n4702) );
  nor2_1 U5132 ( .ip1(n4719), .ip2(n5060), .op(n4701) );
  fulladder U5133 ( .a(n4696), .b(n4695), .ci(n4694), .co(n4684), .s(n4753) );
  xor2_1 U5134 ( .ip1(n4698), .ip2(n4697), .op(n4752) );
  nand2_1 U5135 ( .ip1(n4756), .ip2(n4755), .op(n4764) );
  nor2_1 U5136 ( .ip1(n4718), .ip2(n7813), .op(n4699) );
  xor2_1 U5137 ( .ip1(n4700), .ip2(n4699), .op(n4742) );
  fulladder U5138 ( .a(n4705), .b(n4702), .ci(n4701), .co(n4754), .s(n4741) );
  nor2_1 U5139 ( .ip1(n5475), .ip2(n6107), .op(n4711) );
  nor2_1 U5140 ( .ip1(n4718), .ip2(n5060), .op(n4710) );
  nor2_1 U5141 ( .ip1(n6246), .ip2(n4719), .op(n4709) );
  inv_1 U5142 ( .ip(n4703), .op(n4762) );
  nor3_1 U5143 ( .ip1(n6246), .ip2(n4718), .ip3(n4721), .op(n4745) );
  nand2_1 U5144 ( .ip1(n6280), .ip2(m1Inputs[114]), .op(n4704) );
  or2_1 U5145 ( .ip1(n4704), .ip2(n4705), .op(n4708) );
  nand2_1 U5146 ( .ip1(n6248), .ip2(m1Inputs[115]), .op(n4706) );
  or2_1 U5147 ( .ip1(n4706), .ip2(n4705), .op(n4707) );
  nand2_1 U5148 ( .ip1(n4708), .ip2(n4707), .op(n4744) );
  fulladder U5149 ( .a(n4711), .b(n4710), .ci(n4709), .co(n4740), .s(n4743) );
  nor2_1 U5150 ( .ip1(n5414), .ip2(n4719), .op(n4712) );
  nor3_1 U5151 ( .ip1(n6150), .ip2(n5175), .ip3(n4718), .op(n4713) );
  or2_1 U5152 ( .ip1(n4712), .ip2(n4713), .op(n4716) );
  nand2_1 U5153 ( .ip1(n6280), .ip2(m1Inputs[112]), .op(n4714) );
  or2_1 U5154 ( .ip1(n4714), .ip2(n4713), .op(n4715) );
  nand2_1 U5155 ( .ip1(n4716), .ip2(n4715), .op(n4717) );
  not_ab_or_c_or_d U5156 ( .ip1(n4718), .ip2(n6150), .ip3(n4717), .ip4(n5475), 
        .op(n4725) );
  not_ab_or_c_or_d U5157 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[112]), 
        .ip3(n5593), .ip4(n4719), .op(n4731) );
  nor2_1 U5158 ( .ip1(n5552), .ip2(n7629), .op(n4720) );
  xor2_1 U5159 ( .ip1(n4731), .ip2(n4720), .op(n4727) );
  nand2_1 U5160 ( .ip1(n4725), .ip2(n4727), .op(n4730) );
  or2_1 U5161 ( .ip1(n4721), .ip2(n4745), .op(n4724) );
  nand2_1 U5162 ( .ip1(n8001), .ip2(m1Inputs[112]), .op(n4722) );
  or2_1 U5163 ( .ip1(n4722), .ip2(n4745), .op(n4723) );
  nand2_1 U5164 ( .ip1(n4724), .ip2(n4723), .op(n4726) );
  nand2_1 U5165 ( .ip1(n4725), .ip2(n4726), .op(n4729) );
  nand2_1 U5166 ( .ip1(n4727), .ip2(n4726), .op(n4728) );
  nand3_1 U5167 ( .ip1(n4730), .ip2(n4729), .ip3(n4728), .op(n4736) );
  nand2_1 U5168 ( .ip1(n4734), .ip2(n4736), .op(n4739) );
  nand4_1 U5169 ( .ip1(n6248), .ip2(\STAGE_1/weightReg [2]), .ip3(
        m1Inputs[112]), .ip4(m1Inputs[113]), .op(n4733) );
  nand3_1 U5170 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n4731), .ip3(
        m1Inputs[115]), .op(n4732) );
  nand2_1 U5171 ( .ip1(n4733), .ip2(n4732), .op(n4735) );
  nand2_1 U5172 ( .ip1(n4734), .ip2(n4735), .op(n4738) );
  nand2_1 U5173 ( .ip1(n4736), .ip2(n4735), .op(n4737) );
  nand3_1 U5174 ( .ip1(n4739), .ip2(n4738), .ip3(n4737), .op(n4746) );
  fulladder U5175 ( .a(n4742), .b(n4741), .ci(n4740), .co(n4703), .s(n4748) );
  nand2_1 U5176 ( .ip1(n4746), .ip2(n4748), .op(n4751) );
  fulladder U5177 ( .a(n4745), .b(n4744), .ci(n4743), .co(n4747), .s(n4734) );
  nand2_1 U5178 ( .ip1(n4746), .ip2(n4747), .op(n4750) );
  nand2_1 U5179 ( .ip1(n4748), .ip2(n4747), .op(n4749) );
  nand3_1 U5180 ( .ip1(n4751), .ip2(n4750), .ip3(n4749), .op(n4758) );
  fulladder U5181 ( .a(n4754), .b(n4753), .ci(n4752), .co(n4755), .s(n4757) );
  nand2_1 U5182 ( .ip1(n4758), .ip2(n4757), .op(n4761) );
  nor2_1 U5183 ( .ip1(n4756), .ip2(n4755), .op(n4760) );
  nor2_1 U5184 ( .ip1(n4758), .ip2(n4757), .op(n4759) );
  ab_or_c_or_d U5185 ( .ip1(n4762), .ip2(n4761), .ip3(n4760), .ip4(n4759), 
        .op(n4763) );
  nand2_1 U5186 ( .ip1(n4764), .ip2(n4763), .op(n6132) );
  fulladder U5187 ( .a(n4767), .b(n4766), .ci(n4765), .co(n6131), .s(n4756) );
  inv_1 U5188 ( .ip(m1Inputs[101]), .op(n7496) );
  nor2_1 U5189 ( .ip1(n5552), .ip2(n7496), .op(n4820) );
  inv_1 U5190 ( .ip(m1Inputs[98]), .op(n6062) );
  nor2_1 U5191 ( .ip1(n6246), .ip2(n6062), .op(n4819) );
  inv_1 U5192 ( .ip(m1Inputs[96]), .op(n4823) );
  nor2_1 U5193 ( .ip1(n4823), .ip2(n7813), .op(n4818) );
  nand2_1 U5194 ( .ip1(n6280), .ip2(m1Inputs[100]), .op(n6064) );
  nor3_1 U5195 ( .ip1(n5535), .ip2(n6064), .ip3(n7496), .op(n4803) );
  or2_1 U5196 ( .ip1(n6064), .ip2(n4803), .op(n4770) );
  nand2_1 U5197 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[101]), .op(n4768) );
  or2_1 U5198 ( .ip1(n4768), .ip2(n4803), .op(n4769) );
  nand2_1 U5199 ( .ip1(n4770), .ip2(n4769), .op(n4811) );
  inv_1 U5200 ( .ip(m1Inputs[97]), .op(n4832) );
  nor2_1 U5201 ( .ip1(n4832), .ip2(n7813), .op(n4792) );
  inv_1 U5202 ( .ip(m1Inputs[102]), .op(n7475) );
  nor2_1 U5203 ( .ip1(n5552), .ip2(n7475), .op(n4791) );
  nor2_1 U5204 ( .ip1(n4823), .ip2(n5669), .op(n4790) );
  and3_1 U5205 ( .ip1(n6248), .ip2(m1Inputs[102]), .ip3(n4800), .op(n6058) );
  inv_1 U5206 ( .ip(m1Inputs[100]), .op(n6024) );
  nand2_1 U5207 ( .ip1(n8001), .ip2(m1Inputs[103]), .op(n7443) );
  nor3_1 U5208 ( .ip1(n5552), .ip2(n6024), .ip3(n7443), .op(n4786) );
  nor2_1 U5209 ( .ip1(n6246), .ip2(n6024), .op(n6032) );
  or2_1 U5210 ( .ip1(m1Inputs[103]), .ip2(n6032), .op(n4772) );
  or2_1 U5211 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n6032), .op(n4771) );
  nand2_1 U5212 ( .ip1(n4772), .ip2(n4771), .op(n4785) );
  nand2_1 U5213 ( .ip1(n6280), .ip2(m1Inputs[101]), .op(n4787) );
  nor2_1 U5214 ( .ip1(n4785), .ip2(n4787), .op(n4773) );
  nor2_1 U5215 ( .ip1(n4786), .ip2(n4773), .op(n6048) );
  nand2_1 U5216 ( .ip1(\STAGE_1/weightReg [5]), .ip2(m1Inputs[98]), .op(n4775)
         );
  nand2_1 U5217 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[99]), .op(n4774)
         );
  xor2_1 U5218 ( .ip1(n4775), .ip2(n4774), .op(n4781) );
  inv_1 U5219 ( .ip(m1Inputs[99]), .op(n7444) );
  nand2_1 U5220 ( .ip1(m1Inputs[98]), .ip2(n8078), .op(n4814) );
  nor3_1 U5221 ( .ip1(n7444), .ip2(n7813), .ip3(n4814), .op(n4776) );
  or2_1 U5222 ( .ip1(n4781), .ip2(n4776), .op(n4778) );
  nor2_1 U5223 ( .ip1(n4823), .ip2(n7685), .op(n4780) );
  or2_1 U5224 ( .ip1(n4780), .ip2(n4776), .op(n4777) );
  nand2_1 U5225 ( .ip1(n4778), .ip2(n4777), .op(n6047) );
  nand2_1 U5226 ( .ip1(m1Inputs[98]), .ip2(\STAGE_1/weightReg [6]), .op(n6046)
         );
  inv_1 U5227 ( .ip(n4779), .op(n6055) );
  xnor2_1 U5228 ( .ip1(n4781), .ip2(n4780), .op(n4797) );
  nor3_1 U5229 ( .ip1(n5414), .ip2(n7444), .ip3(n6064), .op(n4809) );
  and2_1 U5230 ( .ip1(\STAGE_1/weightReg [3]), .ip2(n4809), .op(n4784) );
  nand2_1 U5231 ( .ip1(n8001), .ip2(m1Inputs[99]), .op(n4782) );
  mux2_1 U5232 ( .ip1(n4782), .ip2(n8001), .s(n4809), .op(n4813) );
  nor2_1 U5233 ( .ip1(n4814), .ip2(n4813), .op(n4783) );
  nor2_1 U5234 ( .ip1(n4784), .ip2(n4783), .op(n4796) );
  nor2_1 U5235 ( .ip1(n4786), .ip2(n4785), .op(n4788) );
  xor2_1 U5236 ( .ip1(n4788), .ip2(n4787), .op(n4795) );
  inv_1 U5237 ( .ip(n4789), .op(n6054) );
  nor2_1 U5238 ( .ip1(n4832), .ip2(n5669), .op(n4804) );
  fulladder U5239 ( .a(n4792), .b(n4791), .ci(n4790), .co(n4802), .s(n4810) );
  nand2_1 U5240 ( .ip1(m1Inputs[100]), .ip2(n8078), .op(n4794) );
  nand2_1 U5241 ( .ip1(m1Inputs[101]), .ip2(\STAGE_1/weightReg [3]), .op(n4793) );
  xor2_1 U5242 ( .ip1(n4794), .ip2(n4793), .op(n6033) );
  nor2_1 U5243 ( .ip1(n4832), .ip2(n7685), .op(n6035) );
  xor2_1 U5244 ( .ip1(n6033), .ip2(n6035), .op(n6045) );
  nor2_1 U5245 ( .ip1(n7444), .ip2(n7813), .op(n6029) );
  inv_1 U5246 ( .ip(m1Inputs[104]), .op(n7495) );
  nor2_1 U5247 ( .ip1(n5552), .ip2(n7495), .op(n6028) );
  nand2_1 U5248 ( .ip1(m1Inputs[96]), .ip2(\STAGE_1/weightReg [15]), .op(n6027) );
  inv_1 U5249 ( .ip(m1Inputs[103]), .op(n7464) );
  nor2_1 U5250 ( .ip1(n5414), .ip2(n7464), .op(n6031) );
  nand2_1 U5251 ( .ip1(n8175), .ip2(column[96]), .op(n6050) );
  nor2_1 U5252 ( .ip1(n5593), .ip2(n7475), .op(n6030) );
  fulladder U5253 ( .a(n4797), .b(n4796), .ci(n4795), .co(n4789), .s(n4798) );
  inv_1 U5254 ( .ip(n4798), .op(n4882) );
  nor2_1 U5255 ( .ip1(n5414), .ip2(n7475), .op(n4799) );
  nor2_1 U5256 ( .ip1(n4800), .ip2(n4799), .op(n4801) );
  nor2_1 U5257 ( .ip1(n6058), .ip2(n4801), .op(n4881) );
  fulladder U5258 ( .a(n4804), .b(n4803), .ci(n4802), .co(n6053), .s(n4880) );
  nand2_1 U5259 ( .ip1(n6248), .ip2(m1Inputs[98]), .op(n4842) );
  nor3_1 U5260 ( .ip1(n5593), .ip2(n7444), .ip3(n4842), .op(n4828) );
  nor2_1 U5261 ( .ip1(n5593), .ip2(n7444), .op(n4805) );
  or2_1 U5262 ( .ip1(m1Inputs[100]), .ip2(n4805), .op(n4807) );
  or2_1 U5263 ( .ip1(\STAGE_1/weightReg [1]), .ip2(n4805), .op(n4806) );
  nand2_1 U5264 ( .ip1(n4807), .ip2(n4806), .op(n4808) );
  nor2_1 U5265 ( .ip1(n4809), .ip2(n4808), .op(n4822) );
  nor2_1 U5266 ( .ip1(n4832), .ip2(n5060), .op(n4821) );
  fulladder U5267 ( .a(n4812), .b(n4811), .ci(n4810), .co(n4800), .s(n4816) );
  xor2_1 U5268 ( .ip1(n4814), .ip2(n4813), .op(n4815) );
  and2_1 U5269 ( .ip1(n4877), .ip2(n4876), .op(n4871) );
  fulladder U5270 ( .a(n4817), .b(n4816), .ci(n4815), .co(n4876), .s(n4872) );
  fulladder U5271 ( .a(n4820), .b(n4819), .ci(n4818), .co(n4812), .s(n4860) );
  fulladder U5272 ( .a(n4828), .b(n4822), .ci(n4821), .co(n4817), .s(n4859) );
  nor2_1 U5273 ( .ip1(n5552), .ip2(n6024), .op(n4831) );
  nor2_1 U5274 ( .ip1(n4823), .ip2(n5060), .op(n4830) );
  nor2_1 U5275 ( .ip1(n6246), .ip2(n4832), .op(n4829) );
  nor3_1 U5276 ( .ip1(n4871), .ip2(n4872), .ip3(n4873), .op(n4875) );
  nor3_1 U5277 ( .ip1(n6246), .ip2(n4823), .ip3(n4842), .op(n4863) );
  nor2_1 U5278 ( .ip1(n5414), .ip2(n7444), .op(n4824) );
  or2_1 U5279 ( .ip1(m1Inputs[98]), .ip2(n4824), .op(n4826) );
  or2_1 U5280 ( .ip1(\STAGE_1/weightReg [2]), .ip2(n4824), .op(n4825) );
  nand2_1 U5281 ( .ip1(n4826), .ip2(n4825), .op(n4827) );
  nor2_1 U5282 ( .ip1(n4828), .ip2(n4827), .op(n4862) );
  fulladder U5283 ( .a(n4831), .b(n4830), .ci(n4829), .co(n4858), .s(n4861) );
  nand4_1 U5284 ( .ip1(\STAGE_1/weightReg [1]), .ip2(\STAGE_1/weightReg [2]), 
        .ip3(m1Inputs[97]), .ip4(m1Inputs[96]), .op(n4834) );
  not_ab_or_c_or_d U5285 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[96]), 
        .ip3(n5593), .ip4(n4832), .op(n4841) );
  nand3_1 U5286 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n4841), .ip3(m1Inputs[99]), .op(n4833) );
  nand2_1 U5287 ( .ip1(n4834), .ip2(n4833), .op(n4854) );
  nand2_1 U5288 ( .ip1(n4852), .ip2(n4854), .op(n4857) );
  nand2_1 U5289 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[97]), .op(n4839)
         );
  nand2_1 U5290 ( .ip1(n6280), .ip2(m1Inputs[96]), .op(n4838) );
  or2_1 U5291 ( .ip1(m1Inputs[96]), .ip2(m1Inputs[98]), .op(n4836) );
  or2_1 U5292 ( .ip1(n5593), .ip2(m1Inputs[98]), .op(n4835) );
  nand2_1 U5293 ( .ip1(n4836), .ip2(n4835), .op(n4837) );
  not_ab_or_c_or_d U5294 ( .ip1(n4839), .ip2(n4838), .ip3(n4837), .ip4(n5475), 
        .op(n4846) );
  nor2_1 U5295 ( .ip1(n5475), .ip2(n7444), .op(n4840) );
  xor2_1 U5296 ( .ip1(n4841), .ip2(n4840), .op(n4848) );
  nand2_1 U5297 ( .ip1(n4846), .ip2(n4848), .op(n4851) );
  or2_1 U5298 ( .ip1(n4842), .ip2(n4863), .op(n4845) );
  nand2_1 U5299 ( .ip1(n8001), .ip2(m1Inputs[96]), .op(n4843) );
  or2_1 U5300 ( .ip1(n4843), .ip2(n4863), .op(n4844) );
  nand2_1 U5301 ( .ip1(n4845), .ip2(n4844), .op(n4847) );
  nand2_1 U5302 ( .ip1(n4846), .ip2(n4847), .op(n4850) );
  nand2_1 U5303 ( .ip1(n4848), .ip2(n4847), .op(n4849) );
  nand3_1 U5304 ( .ip1(n4851), .ip2(n4850), .ip3(n4849), .op(n4853) );
  nand2_1 U5305 ( .ip1(n4852), .ip2(n4853), .op(n4856) );
  nand2_1 U5306 ( .ip1(n4854), .ip2(n4853), .op(n4855) );
  nand3_1 U5307 ( .ip1(n4857), .ip2(n4856), .ip3(n4855), .op(n4864) );
  fulladder U5308 ( .a(n4860), .b(n4859), .ci(n4858), .co(n4873), .s(n4866) );
  nand2_1 U5309 ( .ip1(n4864), .ip2(n4866), .op(n4869) );
  fulladder U5310 ( .a(n4863), .b(n4862), .ci(n4861), .co(n4865), .s(n4852) );
  nand2_1 U5311 ( .ip1(n4864), .ip2(n4865), .op(n4868) );
  nand2_1 U5312 ( .ip1(n4866), .ip2(n4865), .op(n4867) );
  nand3_1 U5313 ( .ip1(n4869), .ip2(n4868), .ip3(n4867), .op(n4870) );
  not_ab_or_c_or_d U5314 ( .ip1(n4873), .ip2(n4872), .ip3(n4871), .ip4(n4870), 
        .op(n4874) );
  or2_1 U5315 ( .ip1(n4875), .ip2(n4874), .op(n4879) );
  nor2_1 U5316 ( .ip1(n4877), .ip2(n4876), .op(n4878) );
  nor2_1 U5317 ( .ip1(n4879), .ip2(n4878), .op(n6060) );
  fulladder U5318 ( .a(n4882), .b(n4881), .ci(n4880), .co(n6059), .s(n4877) );
  nand2_1 U5319 ( .ip1(m1Inputs[82]), .ip2(\STAGE_1/weightReg [3]), .op(n4884)
         );
  nand2_1 U5320 ( .ip1(m1Inputs[85]), .ip2(\STAGE_1/weightReg [0]), .op(n4883)
         );
  xor2_1 U5321 ( .ip1(n4884), .ip2(n4883), .op(n4976) );
  nand3_1 U5322 ( .ip1(m1Inputs[80]), .ip2(n4976), .ip3(\STAGE_1/weightReg [5]), .op(n4886) );
  nand4_1 U5323 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n8001), .ip3(m1Inputs[82]), .ip4(m1Inputs[85]), .op(n4885) );
  nand2_1 U5324 ( .ip1(n4886), .ip2(n4885), .op(n4936) );
  nand2_1 U5325 ( .ip1(n6280), .ip2(m1Inputs[84]), .op(n5990) );
  inv_1 U5326 ( .ip(m1Inputs[85]), .op(n7306) );
  nor3_1 U5327 ( .ip1(n5414), .ip2(n5990), .ip3(n7306), .op(n4927) );
  or2_1 U5328 ( .ip1(n5990), .ip2(n4927), .op(n4889) );
  nand2_1 U5329 ( .ip1(n6248), .ip2(m1Inputs[85]), .op(n4887) );
  or2_1 U5330 ( .ip1(n4887), .ip2(n4927), .op(n4888) );
  nand2_1 U5331 ( .ip1(n4889), .ip2(n4888), .op(n4935) );
  inv_1 U5332 ( .ip(m1Inputs[81]), .op(n4967) );
  nor2_1 U5333 ( .ip1(n4967), .ip2(n7624), .op(n4912) );
  inv_1 U5334 ( .ip(m1Inputs[86]), .op(n7293) );
  nor2_1 U5335 ( .ip1(n5552), .ip2(n7293), .op(n4911) );
  inv_1 U5336 ( .ip(m1Inputs[80]), .op(n4974) );
  nor2_1 U5337 ( .ip1(n4974), .ip2(n5669), .op(n4910) );
  and3_1 U5338 ( .ip1(n6248), .ip2(m1Inputs[86]), .ip3(n4924), .op(n5985) );
  inv_1 U5339 ( .ip(m1Inputs[84]), .op(n7322) );
  nand2_1 U5340 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[87]), .op(n7256)
         );
  nor3_1 U5341 ( .ip1(n5552), .ip2(n7322), .ip3(n7256), .op(n4906) );
  nor2_1 U5342 ( .ip1(n6246), .ip2(n7322), .op(n4914) );
  or2_1 U5343 ( .ip1(m1Inputs[87]), .ip2(n4914), .op(n4891) );
  or2_1 U5344 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n4914), .op(n4890) );
  nand2_1 U5345 ( .ip1(n4891), .ip2(n4890), .op(n4905) );
  nand2_1 U5346 ( .ip1(n6280), .ip2(m1Inputs[85]), .op(n4907) );
  nor2_1 U5347 ( .ip1(n4905), .ip2(n4907), .op(n4892) );
  nor2_1 U5348 ( .ip1(n4906), .ip2(n4892), .op(n5975) );
  nand2_1 U5349 ( .ip1(n8064), .ip2(m1Inputs[82]), .op(n4894) );
  nand2_1 U5350 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[83]), .op(n4893)
         );
  xor2_1 U5351 ( .ip1(n4894), .ip2(n4893), .op(n4900) );
  inv_1 U5352 ( .ip(m1Inputs[82]), .op(n5989) );
  nand2_1 U5353 ( .ip1(m1Inputs[83]), .ip2(\STAGE_1/weightReg [5]), .op(n5956)
         );
  nor3_1 U5354 ( .ip1(n5989), .ip2(n5060), .ip3(n5956), .op(n4895) );
  or2_1 U5355 ( .ip1(n4900), .ip2(n4895), .op(n4897) );
  nor2_1 U5356 ( .ip1(n4974), .ip2(n7685), .op(n4899) );
  or2_1 U5357 ( .ip1(n4899), .ip2(n4895), .op(n4896) );
  nand2_1 U5358 ( .ip1(n4897), .ip2(n4896), .op(n5974) );
  inv_1 U5359 ( .ip(n5669), .op(n8037) );
  nand2_1 U5360 ( .ip1(m1Inputs[82]), .ip2(n8037), .op(n5973) );
  inv_1 U5361 ( .ip(n4898), .op(n5982) );
  xnor2_1 U5362 ( .ip1(n4900), .ip2(n4899), .op(n4921) );
  nor2_1 U5363 ( .ip1(n5989), .ip2(n5060), .op(n4938) );
  inv_1 U5364 ( .ip(m1Inputs[83]), .op(n7253) );
  nor3_1 U5365 ( .ip1(n5414), .ip2(n7253), .ip3(n5990), .op(n4933) );
  and2_1 U5366 ( .ip1(\STAGE_1/weightReg [3]), .ip2(n4933), .op(n4902) );
  or2_1 U5367 ( .ip1(n4938), .ip2(n4902), .op(n4904) );
  nor2_1 U5368 ( .ip1(n4933), .ip2(n7253), .op(n4901) );
  mux2_1 U5369 ( .ip1(n4901), .ip2(n4933), .s(n5500), .op(n4937) );
  or2_1 U5370 ( .ip1(n4937), .ip2(n4902), .op(n4903) );
  nand2_1 U5371 ( .ip1(n4904), .ip2(n4903), .op(n4920) );
  nor2_1 U5372 ( .ip1(n4906), .ip2(n4905), .op(n4908) );
  xor2_1 U5373 ( .ip1(n4908), .ip2(n4907), .op(n4919) );
  inv_1 U5374 ( .ip(n4909), .op(n5981) );
  nor2_1 U5375 ( .ip1(n4967), .ip2(n5669), .op(n4928) );
  fulladder U5376 ( .a(n4912), .b(n4911), .ci(n4910), .co(n4926), .s(n4934) );
  inv_1 U5377 ( .ip(\STAGE_1/weightReg [15]), .op(n7628) );
  nor2_1 U5378 ( .ip1(n4974), .ip2(n7628), .op(n5958) );
  nand2_1 U5379 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[88]), .op(n5957)
         );
  inv_1 U5380 ( .ip(n4913), .op(n5972) );
  nor2_1 U5381 ( .ip1(n5060), .ip2(n7306), .op(n6011) );
  and2_1 U5382 ( .ip1(n6011), .ip2(n4914), .op(n5962) );
  nor2_1 U5383 ( .ip1(n6246), .ip2(n7306), .op(n4915) );
  or2_1 U5384 ( .ip1(m1Inputs[84]), .ip2(n4915), .op(n4917) );
  or2_1 U5385 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n4915), .op(n4916) );
  nand2_1 U5386 ( .ip1(n4917), .ip2(n4916), .op(n4918) );
  nor2_1 U5387 ( .ip1(n5962), .ip2(n4918), .op(n5961) );
  nor2_1 U5388 ( .ip1(n4967), .ip2(n7685), .op(n5963) );
  xor2_1 U5389 ( .ip1(n5961), .ip2(n5963), .op(n5971) );
  inv_1 U5390 ( .ip(m1Inputs[87]), .op(n7279) );
  nor2_1 U5391 ( .ip1(n5414), .ip2(n7279), .op(n5954) );
  nor2_1 U5392 ( .ip1(n5593), .ip2(n7293), .op(n5953) );
  nand2_1 U5393 ( .ip1(n8009), .ip2(column[80]), .op(n5977) );
  fulladder U5394 ( .a(n4921), .b(n4920), .ci(n4919), .co(n4909), .s(n4922) );
  inv_1 U5395 ( .ip(n4922), .op(n5007) );
  nor2_1 U5396 ( .ip1(n5414), .ip2(n7293), .op(n4923) );
  nor2_1 U5397 ( .ip1(n4924), .ip2(n4923), .op(n4925) );
  nor2_1 U5398 ( .ip1(n5985), .ip2(n4925), .op(n5006) );
  fulladder U5399 ( .a(n4928), .b(n4927), .ci(n4926), .co(n5980), .s(n5005) );
  nand2_1 U5400 ( .ip1(n6248), .ip2(m1Inputs[82]), .op(n4943) );
  nor3_1 U5401 ( .ip1(n5593), .ip2(n7253), .ip3(n4943), .op(n4979) );
  nor2_1 U5402 ( .ip1(n5593), .ip2(n7253), .op(n4929) );
  or2_1 U5403 ( .ip1(m1Inputs[84]), .ip2(n4929), .op(n4931) );
  or2_1 U5404 ( .ip1(\STAGE_1/weightReg [1]), .ip2(n4929), .op(n4930) );
  nand2_1 U5405 ( .ip1(n4931), .ip2(n4930), .op(n4932) );
  nor2_1 U5406 ( .ip1(n4933), .ip2(n4932), .op(n4978) );
  nor2_1 U5407 ( .ip1(n4967), .ip2(n5060), .op(n4977) );
  fulladder U5408 ( .a(n4936), .b(n4935), .ci(n4934), .co(n4924), .s(n4940) );
  xor2_1 U5409 ( .ip1(n4938), .ip2(n4937), .op(n4939) );
  nand2_1 U5410 ( .ip1(n4996), .ip2(n4995), .op(n5004) );
  fulladder U5411 ( .a(n4941), .b(n4940), .ci(n4939), .co(n4995), .s(n4942) );
  inv_1 U5412 ( .ip(n4942), .op(n5002) );
  nor3_1 U5413 ( .ip1(n6246), .ip2(n4974), .ip3(n4943), .op(n4985) );
  or2_1 U5414 ( .ip1(n4943), .ip2(n4985), .op(n4946) );
  nand2_1 U5415 ( .ip1(n8001), .ip2(m1Inputs[80]), .op(n4944) );
  or2_1 U5416 ( .ip1(n4944), .ip2(n4985), .op(n4945) );
  nand2_1 U5417 ( .ip1(n4946), .ip2(n4945), .op(n4954) );
  not_ab_or_c_or_d U5418 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[80]), 
        .ip3(n5593), .ip4(n4967), .op(n4960) );
  nor2_1 U5419 ( .ip1(n5552), .ip2(n7253), .op(n4947) );
  xor2_1 U5420 ( .ip1(n4960), .ip2(n4947), .op(n4956) );
  nand2_1 U5421 ( .ip1(n4954), .ip2(n4956), .op(n4959) );
  nor2_1 U5422 ( .ip1(n5414), .ip2(n4967), .op(n4948) );
  nor3_1 U5423 ( .ip1(n5989), .ip2(n5175), .ip3(n4974), .op(n4949) );
  or2_1 U5424 ( .ip1(n4948), .ip2(n4949), .op(n4952) );
  nand2_1 U5425 ( .ip1(n6280), .ip2(m1Inputs[80]), .op(n4950) );
  or2_1 U5426 ( .ip1(n4950), .ip2(n4949), .op(n4951) );
  nand2_1 U5427 ( .ip1(n4952), .ip2(n4951), .op(n4953) );
  not_ab_or_c_or_d U5428 ( .ip1(n4974), .ip2(n5989), .ip3(n4953), .ip4(n5552), 
        .op(n4955) );
  nand2_1 U5429 ( .ip1(n4954), .ip2(n4955), .op(n4958) );
  nand2_1 U5430 ( .ip1(n4956), .ip2(n4955), .op(n4957) );
  nand3_1 U5431 ( .ip1(n4959), .ip2(n4958), .ip3(n4957), .op(n4968) );
  nand4_1 U5432 ( .ip1(n6248), .ip2(\STAGE_1/weightReg [2]), .ip3(m1Inputs[81]), .ip4(m1Inputs[80]), .op(n4962) );
  nand3_1 U5433 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n4960), .ip3(m1Inputs[83]), .op(n4961) );
  nand2_1 U5434 ( .ip1(n4962), .ip2(n4961), .op(n4970) );
  nand2_1 U5435 ( .ip1(n4968), .ip2(n4970), .op(n4973) );
  nand2_1 U5436 ( .ip1(n6280), .ip2(m1Inputs[82]), .op(n4963) );
  or2_1 U5437 ( .ip1(n4963), .ip2(n4979), .op(n4966) );
  nand2_1 U5438 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[83]), .op(n4964)
         );
  or2_1 U5439 ( .ip1(n4964), .ip2(n4979), .op(n4965) );
  nand2_1 U5440 ( .ip1(n4966), .ip2(n4965), .op(n4984) );
  nor2_1 U5441 ( .ip1(n5552), .ip2(n7322), .op(n4982) );
  nor2_1 U5442 ( .ip1(n4974), .ip2(n5060), .op(n4981) );
  nor2_1 U5443 ( .ip1(n6246), .ip2(n4967), .op(n4980) );
  nand2_1 U5444 ( .ip1(n4968), .ip2(n4969), .op(n4972) );
  nand2_1 U5445 ( .ip1(n4970), .ip2(n4969), .op(n4971) );
  nand3_1 U5446 ( .ip1(n4973), .ip2(n4972), .ip3(n4971), .op(n4986) );
  nor2_1 U5447 ( .ip1(n4974), .ip2(n7813), .op(n4975) );
  xor2_1 U5448 ( .ip1(n4976), .ip2(n4975), .op(n4994) );
  fulladder U5449 ( .a(n4979), .b(n4978), .ci(n4977), .co(n4941), .s(n4993) );
  fulladder U5450 ( .a(n4982), .b(n4981), .ci(n4980), .co(n4992), .s(n4983) );
  nand2_1 U5451 ( .ip1(n4986), .ip2(n4988), .op(n4991) );
  fulladder U5452 ( .a(n4985), .b(n4984), .ci(n4983), .co(n4987), .s(n4969) );
  nand2_1 U5453 ( .ip1(n4986), .ip2(n4987), .op(n4990) );
  nand2_1 U5454 ( .ip1(n4988), .ip2(n4987), .op(n4989) );
  nand3_1 U5455 ( .ip1(n4991), .ip2(n4990), .ip3(n4989), .op(n4998) );
  fulladder U5456 ( .a(n4994), .b(n4993), .ci(n4992), .co(n4997), .s(n4988) );
  nand2_1 U5457 ( .ip1(n4998), .ip2(n4997), .op(n5001) );
  nor2_1 U5458 ( .ip1(n4996), .ip2(n4995), .op(n5000) );
  nor2_1 U5459 ( .ip1(n4998), .ip2(n4997), .op(n4999) );
  ab_or_c_or_d U5460 ( .ip1(n5002), .ip2(n5001), .ip3(n5000), .ip4(n4999), 
        .op(n5003) );
  nand2_1 U5461 ( .ip1(n5004), .ip2(n5003), .op(n5987) );
  fulladder U5462 ( .a(n5007), .b(n5006), .ci(n5005), .co(n5986), .s(n4996) );
  inv_1 U5463 ( .ip(m1Inputs[69]), .op(n7122) );
  nor2_1 U5464 ( .ip1(n5552), .ip2(n7122), .op(n5065) );
  inv_1 U5465 ( .ip(m1Inputs[66]), .op(n5931) );
  nor2_1 U5466 ( .ip1(n6246), .ip2(n5931), .op(n5064) );
  inv_1 U5467 ( .ip(m1Inputs[64]), .op(n5089) );
  nor2_1 U5468 ( .ip1(n5089), .ip2(n7624), .op(n5063) );
  nand2_1 U5469 ( .ip1(n6280), .ip2(m1Inputs[68]), .op(n5933) );
  nor3_1 U5470 ( .ip1(n5414), .ip2(n5933), .ip3(n7122), .op(n5054) );
  or2_1 U5471 ( .ip1(n5933), .ip2(n5054), .op(n5010) );
  nand2_1 U5472 ( .ip1(n6248), .ip2(m1Inputs[69]), .op(n5008) );
  or2_1 U5473 ( .ip1(n5008), .ip2(n5054), .op(n5009) );
  nand2_1 U5474 ( .ip1(n5010), .ip2(n5009), .op(n5042) );
  inv_1 U5475 ( .ip(m1Inputs[65]), .op(n5078) );
  nor2_1 U5476 ( .ip1(n5078), .ip2(n7624), .op(n5033) );
  inv_1 U5477 ( .ip(m1Inputs[70]), .op(n7101) );
  nor2_1 U5478 ( .ip1(n5552), .ip2(n7101), .op(n5032) );
  nor2_1 U5479 ( .ip1(n5089), .ip2(n5669), .op(n5031) );
  and3_1 U5480 ( .ip1(n6248), .ip2(m1Inputs[70]), .ip3(n5051), .op(n5911) );
  inv_1 U5481 ( .ip(m1Inputs[68]), .op(n5879) );
  nand2_1 U5482 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[71]), .op(n7069)
         );
  nor3_1 U5483 ( .ip1(n5475), .ip2(n5879), .ip3(n7069), .op(n5027) );
  nor2_1 U5484 ( .ip1(n6246), .ip2(n5879), .op(n5011) );
  or2_1 U5485 ( .ip1(m1Inputs[71]), .ip2(n5011), .op(n5013) );
  or2_1 U5486 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n5011), .op(n5012) );
  nand2_1 U5487 ( .ip1(n5013), .ip2(n5012), .op(n5026) );
  nand2_1 U5488 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[69]), .op(n5028)
         );
  nor2_1 U5489 ( .ip1(n5026), .ip2(n5028), .op(n5014) );
  nor2_1 U5490 ( .ip1(n5027), .ip2(n5014), .op(n5901) );
  nand2_1 U5491 ( .ip1(n8064), .ip2(m1Inputs[66]), .op(n5016) );
  nand2_1 U5492 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[67]), .op(n5015)
         );
  xor2_1 U5493 ( .ip1(n5016), .ip2(n5015), .op(n5022) );
  inv_1 U5494 ( .ip(m1Inputs[67]), .op(n7070) );
  nand2_1 U5495 ( .ip1(m1Inputs[66]), .ip2(n8078), .op(n5045) );
  nor3_1 U5496 ( .ip1(n7070), .ip2(n7624), .ip3(n5045), .op(n5017) );
  or2_1 U5497 ( .ip1(n5022), .ip2(n5017), .op(n5019) );
  nor2_1 U5498 ( .ip1(n5089), .ip2(n7685), .op(n5021) );
  or2_1 U5499 ( .ip1(n5021), .ip2(n5017), .op(n5018) );
  nand2_1 U5500 ( .ip1(n5019), .ip2(n5018), .op(n5900) );
  nand2_1 U5501 ( .ip1(m1Inputs[66]), .ip2(n8037), .op(n5899) );
  inv_1 U5502 ( .ip(n5020), .op(n5908) );
  xnor2_1 U5503 ( .ip1(n5022), .ip2(n5021), .op(n5048) );
  nand2_1 U5504 ( .ip1(n6248), .ip2(m1Inputs[67]), .op(n5919) );
  nor2_1 U5505 ( .ip1(n5933), .ip2(n5919), .op(n5040) );
  and2_1 U5506 ( .ip1(\STAGE_1/weightReg [3]), .ip2(n5040), .op(n5025) );
  nand2_1 U5507 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[67]), .op(n5023)
         );
  mux2_1 U5508 ( .ip1(n5023), .ip2(n8001), .s(n5040), .op(n5044) );
  nor2_1 U5509 ( .ip1(n5045), .ip2(n5044), .op(n5024) );
  nor2_1 U5510 ( .ip1(n5025), .ip2(n5024), .op(n5047) );
  nor2_1 U5511 ( .ip1(n5027), .ip2(n5026), .op(n5029) );
  xor2_1 U5512 ( .ip1(n5029), .ip2(n5028), .op(n5046) );
  inv_1 U5513 ( .ip(n5030), .op(n5907) );
  nor2_1 U5514 ( .ip1(n5078), .ip2(n5669), .op(n5055) );
  fulladder U5515 ( .a(n5033), .b(n5032), .ci(n5031), .co(n5053), .s(n5041) );
  nand2_1 U5516 ( .ip1(m1Inputs[69]), .ip2(\STAGE_1/weightReg [3]), .op(n5035)
         );
  nor2_1 U5517 ( .ip1(n5879), .ip2(n5060), .op(n5034) );
  xor2_1 U5518 ( .ip1(n5035), .ip2(n5034), .op(n5888) );
  nand2_1 U5519 ( .ip1(m1Inputs[65]), .ip2(n7882), .op(n5887) );
  xor2_1 U5520 ( .ip1(n5888), .ip2(n5887), .op(n5898) );
  nor2_1 U5521 ( .ip1(n7070), .ip2(n7624), .op(n5884) );
  inv_1 U5522 ( .ip(m1Inputs[72]), .op(n7121) );
  nor2_1 U5523 ( .ip1(n5552), .ip2(n7121), .op(n5883) );
  nand2_1 U5524 ( .ip1(m1Inputs[64]), .ip2(\STAGE_1/weightReg [15]), .op(n5882) );
  inv_1 U5525 ( .ip(m1Inputs[71]), .op(n7090) );
  nor2_1 U5526 ( .ip1(n5414), .ip2(n7090), .op(n5886) );
  nand2_1 U5527 ( .ip1(n8009), .ip2(column[64]), .op(n5903) );
  nor2_1 U5528 ( .ip1(n5593), .ip2(n7101), .op(n5885) );
  nand2_1 U5529 ( .ip1(n6248), .ip2(m1Inputs[66]), .op(n5088) );
  nor3_1 U5530 ( .ip1(n5593), .ip2(n7070), .ip3(n5088), .op(n5069) );
  nor2_1 U5531 ( .ip1(n5593), .ip2(n7070), .op(n5036) );
  or2_1 U5532 ( .ip1(m1Inputs[68]), .ip2(n5036), .op(n5038) );
  or2_1 U5533 ( .ip1(\STAGE_1/weightReg [1]), .ip2(n5036), .op(n5037) );
  nand2_1 U5534 ( .ip1(n5038), .ip2(n5037), .op(n5039) );
  nor2_1 U5535 ( .ip1(n5040), .ip2(n5039), .op(n5062) );
  nor2_1 U5536 ( .ip1(n5078), .ip2(n5060), .op(n5061) );
  fulladder U5537 ( .a(n5043), .b(n5042), .ci(n5041), .co(n5051), .s(n5057) );
  xor2_1 U5538 ( .ip1(n5045), .ip2(n5044), .op(n5056) );
  fulladder U5539 ( .a(n5048), .b(n5047), .ci(n5046), .co(n5030), .s(n5049) );
  inv_1 U5540 ( .ip(n5049), .op(n5122) );
  nor2_1 U5541 ( .ip1(n5414), .ip2(n7101), .op(n5050) );
  nor2_1 U5542 ( .ip1(n5051), .ip2(n5050), .op(n5052) );
  nor2_1 U5543 ( .ip1(n5911), .ip2(n5052), .op(n5121) );
  fulladder U5544 ( .a(n5055), .b(n5054), .ci(n5053), .co(n5906), .s(n5120) );
  nand2_1 U5545 ( .ip1(n5111), .ip2(n5110), .op(n5119) );
  fulladder U5546 ( .a(n5058), .b(n5057), .ci(n5056), .co(n5111), .s(n5059) );
  inv_1 U5547 ( .ip(n5059), .op(n5117) );
  nor2_1 U5548 ( .ip1(n5552), .ip2(n5879), .op(n5068) );
  nor2_1 U5549 ( .ip1(n5089), .ip2(n5060), .op(n5067) );
  nor2_1 U5550 ( .ip1(n6246), .ip2(n5078), .op(n5066) );
  fulladder U5551 ( .a(n5069), .b(n5062), .ci(n5061), .co(n5058), .s(n5074) );
  fulladder U5552 ( .a(n5065), .b(n5064), .ci(n5063), .co(n5043), .s(n5073) );
  fulladder U5553 ( .a(n5068), .b(n5067), .ci(n5066), .co(n5075), .s(n5077) );
  nor3_1 U5554 ( .ip1(n6246), .ip2(n5089), .ip3(n5088), .op(n5093) );
  or2_1 U5555 ( .ip1(n5919), .ip2(n5069), .op(n5072) );
  nand2_1 U5556 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[66]), .op(n5070)
         );
  or2_1 U5557 ( .ip1(n5070), .ip2(n5069), .op(n5071) );
  nand2_1 U5558 ( .ip1(n5072), .ip2(n5071), .op(n5076) );
  fulladder U5559 ( .a(n5075), .b(n5074), .ci(n5073), .co(n5113), .s(n5106) );
  nand2_1 U5560 ( .ip1(n5104), .ip2(n5106), .op(n5109) );
  fulladder U5561 ( .a(n5077), .b(n5093), .ci(n5076), .co(n5104), .s(n5098) );
  nand4_1 U5562 ( .ip1(n6248), .ip2(\STAGE_1/weightReg [2]), .ip3(m1Inputs[65]), .ip4(m1Inputs[64]), .op(n5080) );
  not_ab_or_c_or_d U5563 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[64]), 
        .ip3(n5593), .ip4(n5078), .op(n5087) );
  nand3_1 U5564 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n5087), .ip3(m1Inputs[67]), .op(n5079) );
  nand2_1 U5565 ( .ip1(n5080), .ip2(n5079), .op(n5100) );
  nand2_1 U5566 ( .ip1(n5098), .ip2(n5100), .op(n5103) );
  nand2_1 U5567 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[65]), .op(n5085)
         );
  nand2_1 U5568 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[64]), .op(n5084)
         );
  or2_1 U5569 ( .ip1(m1Inputs[64]), .ip2(m1Inputs[66]), .op(n5082) );
  or2_1 U5570 ( .ip1(n5593), .ip2(m1Inputs[66]), .op(n5081) );
  nand2_1 U5571 ( .ip1(n5082), .ip2(n5081), .op(n5083) );
  ab_or_c_or_d U5572 ( .ip1(n5085), .ip2(n5084), .ip3(n5083), .ip4(n5475), 
        .op(n5094) );
  nand2_1 U5573 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[67]), .op(n5086)
         );
  xor2_1 U5574 ( .ip1(n5087), .ip2(n5086), .op(n5095) );
  nor2_1 U5575 ( .ip1(n5094), .ip2(n5095), .op(n5097) );
  inv_1 U5576 ( .ip(n5088), .op(n5091) );
  nor2_1 U5577 ( .ip1(n6246), .ip2(n5089), .op(n5090) );
  nor2_1 U5578 ( .ip1(n5091), .ip2(n5090), .op(n5092) );
  not_ab_or_c_or_d U5579 ( .ip1(n5095), .ip2(n5094), .ip3(n5093), .ip4(n5092), 
        .op(n5096) );
  or2_1 U5580 ( .ip1(n5097), .ip2(n5096), .op(n5099) );
  nand2_1 U5581 ( .ip1(n5098), .ip2(n5099), .op(n5102) );
  nand2_1 U5582 ( .ip1(n5100), .ip2(n5099), .op(n5101) );
  nand3_1 U5583 ( .ip1(n5103), .ip2(n5102), .ip3(n5101), .op(n5105) );
  nand2_1 U5584 ( .ip1(n5104), .ip2(n5105), .op(n5108) );
  nand2_1 U5585 ( .ip1(n5106), .ip2(n5105), .op(n5107) );
  nand3_1 U5586 ( .ip1(n5109), .ip2(n5108), .ip3(n5107), .op(n5112) );
  nand2_1 U5587 ( .ip1(n5113), .ip2(n5112), .op(n5116) );
  nor2_1 U5588 ( .ip1(n5111), .ip2(n5110), .op(n5115) );
  nor2_1 U5589 ( .ip1(n5113), .ip2(n5112), .op(n5114) );
  ab_or_c_or_d U5590 ( .ip1(n5117), .ip2(n5116), .ip3(n5115), .ip4(n5114), 
        .op(n5118) );
  nand2_1 U5591 ( .ip1(n5119), .ip2(n5118), .op(n5913) );
  fulladder U5592 ( .a(n5122), .b(n5121), .ci(n5120), .co(n5912), .s(n5110) );
  inv_1 U5593 ( .ip(m1Inputs[53]), .op(n6931) );
  nor2_1 U5594 ( .ip1(n5552), .ip2(n6931), .op(n5172) );
  inv_1 U5595 ( .ip(m1Inputs[50]), .op(n5844) );
  nor2_1 U5596 ( .ip1(n5844), .ip2(n5500), .op(n5171) );
  inv_1 U5597 ( .ip(m1Inputs[48]), .op(n5187) );
  nor2_1 U5598 ( .ip1(n5187), .ip2(n7624), .op(n5170) );
  nand2_1 U5599 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[52]), .op(n5846)
         );
  nor3_1 U5600 ( .ip1(n5414), .ip2(n5846), .ip3(n6931), .op(n5158) );
  or2_1 U5601 ( .ip1(n5846), .ip2(n5158), .op(n5125) );
  nand2_1 U5602 ( .ip1(n6248), .ip2(m1Inputs[53]), .op(n5123) );
  or2_1 U5603 ( .ip1(n5123), .ip2(n5158), .op(n5124) );
  nand2_1 U5604 ( .ip1(n5125), .ip2(n5124), .op(n5166) );
  inv_1 U5605 ( .ip(m1Inputs[49]), .op(n5176) );
  nor2_1 U5606 ( .ip1(n5176), .ip2(n7624), .op(n5147) );
  inv_1 U5607 ( .ip(m1Inputs[54]), .op(n6918) );
  nor2_1 U5608 ( .ip1(n5552), .ip2(n6918), .op(n5146) );
  nor2_1 U5609 ( .ip1(n5187), .ip2(n5669), .op(n5145) );
  and3_1 U5610 ( .ip1(n6248), .ip2(m1Inputs[54]), .ip3(n5155), .op(n5840) );
  inv_1 U5611 ( .ip(m1Inputs[52]), .op(n6947) );
  nand2_1 U5612 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[55]), .op(n6885)
         );
  nor3_1 U5613 ( .ip1(n5475), .ip2(n6947), .ip3(n6885), .op(n5141) );
  nor2_1 U5614 ( .ip1(n6246), .ip2(n6947), .op(n5815) );
  or2_1 U5615 ( .ip1(m1Inputs[55]), .ip2(n5815), .op(n5127) );
  or2_1 U5616 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n5815), .op(n5126) );
  nand2_1 U5617 ( .ip1(n5127), .ip2(n5126), .op(n5140) );
  nand2_1 U5618 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[53]), .op(n5142)
         );
  nor2_1 U5619 ( .ip1(n5140), .ip2(n5142), .op(n5128) );
  nor2_1 U5620 ( .ip1(n5141), .ip2(n5128), .op(n5830) );
  nand2_1 U5621 ( .ip1(n8064), .ip2(m1Inputs[50]), .op(n5130) );
  nand2_1 U5622 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[51]), .op(n5129)
         );
  xor2_1 U5623 ( .ip1(n5130), .ip2(n5129), .op(n5136) );
  inv_1 U5624 ( .ip(m1Inputs[51]), .op(n6886) );
  nand2_1 U5625 ( .ip1(m1Inputs[50]), .ip2(\STAGE_1/weightReg [4]), .op(n5169)
         );
  nor3_1 U5626 ( .ip1(n6886), .ip2(n7813), .ip3(n5169), .op(n5131) );
  or2_1 U5627 ( .ip1(n5136), .ip2(n5131), .op(n5133) );
  nor2_1 U5628 ( .ip1(n5187), .ip2(n7685), .op(n5135) );
  or2_1 U5629 ( .ip1(n5135), .ip2(n5131), .op(n5132) );
  nand2_1 U5630 ( .ip1(n5133), .ip2(n5132), .op(n5829) );
  nand2_1 U5631 ( .ip1(m1Inputs[50]), .ip2(\STAGE_1/weightReg [6]), .op(n5828)
         );
  inv_1 U5632 ( .ip(n5134), .op(n5837) );
  xnor2_1 U5633 ( .ip1(n5136), .ip2(n5135), .op(n5152) );
  nor3_1 U5634 ( .ip1(n6886), .ip2(n5414), .ip3(n5846), .op(n5164) );
  and2_1 U5635 ( .ip1(\STAGE_1/weightReg [3]), .ip2(n5164), .op(n5139) );
  nand2_1 U5636 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[51]), .op(n5137)
         );
  mux2_1 U5637 ( .ip1(n5137), .ip2(n8001), .s(n5164), .op(n5168) );
  nor2_1 U5638 ( .ip1(n5169), .ip2(n5168), .op(n5138) );
  nor2_1 U5639 ( .ip1(n5139), .ip2(n5138), .op(n5151) );
  nor2_1 U5640 ( .ip1(n5141), .ip2(n5140), .op(n5143) );
  xor2_1 U5641 ( .ip1(n5143), .ip2(n5142), .op(n5150) );
  inv_1 U5642 ( .ip(n5144), .op(n5836) );
  nor2_1 U5643 ( .ip1(n5176), .ip2(n5669), .op(n5159) );
  fulladder U5644 ( .a(n5147), .b(n5146), .ci(n5145), .co(n5157), .s(n5165) );
  nand2_1 U5645 ( .ip1(m1Inputs[53]), .ip2(\STAGE_1/weightReg [3]), .op(n5149)
         );
  nor2_1 U5646 ( .ip1(n6947), .ip2(n5060), .op(n5148) );
  xor2_1 U5647 ( .ip1(n5149), .ip2(n5148), .op(n5817) );
  nand2_1 U5648 ( .ip1(m1Inputs[49]), .ip2(\STAGE_1/weightReg [7]), .op(n5816)
         );
  xor2_1 U5649 ( .ip1(n5817), .ip2(n5816), .op(n5827) );
  nor2_1 U5650 ( .ip1(n6886), .ip2(n7813), .op(n5812) );
  inv_1 U5651 ( .ip(m1Inputs[56]), .op(n6906) );
  nor2_1 U5652 ( .ip1(n5552), .ip2(n6906), .op(n5811) );
  nand2_1 U5653 ( .ip1(m1Inputs[48]), .ip2(\STAGE_1/weightReg [15]), .op(n5810) );
  inv_1 U5654 ( .ip(m1Inputs[55]), .op(n6907) );
  nor2_1 U5655 ( .ip1(n5414), .ip2(n6907), .op(n5814) );
  nand2_1 U5656 ( .ip1(n8009), .ip2(column[48]), .op(n5832) );
  nor2_1 U5657 ( .ip1(n5593), .ip2(n6918), .op(n5813) );
  fulladder U5658 ( .a(n5152), .b(n5151), .ci(n5150), .co(n5144), .s(n5153) );
  inv_1 U5659 ( .ip(n5153), .op(n5239) );
  nor2_1 U5660 ( .ip1(n5535), .ip2(n6918), .op(n5154) );
  nor2_1 U5661 ( .ip1(n5155), .ip2(n5154), .op(n5156) );
  nor2_1 U5662 ( .ip1(n5840), .ip2(n5156), .op(n5238) );
  fulladder U5663 ( .a(n5159), .b(n5158), .ci(n5157), .co(n5835), .s(n5237) );
  nand2_1 U5664 ( .ip1(n6248), .ip2(m1Inputs[50]), .op(n5188) );
  nor3_1 U5665 ( .ip1(n6886), .ip2(n5593), .ip3(n5188), .op(n5202) );
  nor2_1 U5666 ( .ip1(n6886), .ip2(n5593), .op(n5160) );
  or2_1 U5667 ( .ip1(m1Inputs[52]), .ip2(n5160), .op(n5162) );
  or2_1 U5668 ( .ip1(\STAGE_1/weightReg [1]), .ip2(n5160), .op(n5161) );
  nand2_1 U5669 ( .ip1(n5162), .ip2(n5161), .op(n5163) );
  nor2_1 U5670 ( .ip1(n5164), .ip2(n5163), .op(n5174) );
  nor2_1 U5671 ( .ip1(n5176), .ip2(n5060), .op(n5173) );
  fulladder U5672 ( .a(n5167), .b(n5166), .ci(n5165), .co(n5155), .s(n5225) );
  xor2_1 U5673 ( .ip1(n5169), .ip2(n5168), .op(n5224) );
  and2_1 U5674 ( .ip1(n5234), .ip2(n5233), .op(n5228) );
  fulladder U5675 ( .a(n5172), .b(n5171), .ci(n5170), .co(n5167), .s(n5214) );
  fulladder U5676 ( .a(n5202), .b(n5174), .ci(n5173), .co(n5226), .s(n5213) );
  nor2_1 U5677 ( .ip1(n5552), .ip2(n6947), .op(n5205) );
  nor2_1 U5678 ( .ip1(n5187), .ip2(n5060), .op(n5204) );
  nor2_1 U5679 ( .ip1(n5176), .ip2(n5500), .op(n5203) );
  nor2_1 U5680 ( .ip1(n5552), .ip2(n6886), .op(n5184) );
  nor4_1 U5681 ( .ip1(n5414), .ip2(n5176), .ip3(n5175), .ip4(n5187), .op(n5183) );
  nor2_1 U5682 ( .ip1(n5184), .ip2(n5183), .op(n5177) );
  nand2_1 U5683 ( .ip1(m1Inputs[49]), .ip2(\STAGE_1/weightReg [2]), .op(n5186)
         );
  nor2_1 U5684 ( .ip1(n5177), .ip2(n5186), .op(n5206) );
  nand2_1 U5685 ( .ip1(n6248), .ip2(m1Inputs[49]), .op(n5182) );
  nand2_1 U5686 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[48]), .op(n5181)
         );
  or2_1 U5687 ( .ip1(m1Inputs[48]), .ip2(m1Inputs[50]), .op(n5179) );
  or2_1 U5688 ( .ip1(n5593), .ip2(m1Inputs[50]), .op(n5178) );
  nand2_1 U5689 ( .ip1(n5179), .ip2(n5178), .op(n5180) );
  not_ab_or_c_or_d U5690 ( .ip1(n5182), .ip2(n5181), .ip3(n5180), .ip4(n5475), 
        .op(n5192) );
  xnor2_1 U5691 ( .ip1(n5184), .ip2(n5183), .op(n5185) );
  xor2_1 U5692 ( .ip1(n5186), .ip2(n5185), .op(n5194) );
  nand2_1 U5693 ( .ip1(n5192), .ip2(n5194), .op(n5197) );
  nor3_1 U5694 ( .ip1(n5187), .ip2(n5188), .ip3(n5500), .op(n5217) );
  or2_1 U5695 ( .ip1(n5188), .ip2(n5217), .op(n5191) );
  nand2_1 U5696 ( .ip1(m1Inputs[48]), .ip2(\STAGE_1/weightReg [3]), .op(n5189)
         );
  or2_1 U5697 ( .ip1(n5189), .ip2(n5217), .op(n5190) );
  nand2_1 U5698 ( .ip1(n5191), .ip2(n5190), .op(n5193) );
  nand2_1 U5699 ( .ip1(n5192), .ip2(n5193), .op(n5196) );
  nand2_1 U5700 ( .ip1(n5194), .ip2(n5193), .op(n5195) );
  nand3_1 U5701 ( .ip1(n5197), .ip2(n5196), .ip3(n5195), .op(n5208) );
  nand2_1 U5702 ( .ip1(n5206), .ip2(n5208), .op(n5211) );
  nor2_1 U5703 ( .ip1(n6886), .ip2(n5414), .op(n5198) );
  or2_1 U5704 ( .ip1(m1Inputs[50]), .ip2(n5198), .op(n5200) );
  or2_1 U5705 ( .ip1(\STAGE_1/weightReg [2]), .ip2(n5198), .op(n5199) );
  nand2_1 U5706 ( .ip1(n5200), .ip2(n5199), .op(n5201) );
  nor2_1 U5707 ( .ip1(n5202), .ip2(n5201), .op(n5216) );
  fulladder U5708 ( .a(n5205), .b(n5204), .ci(n5203), .co(n5212), .s(n5215) );
  nand2_1 U5709 ( .ip1(n5206), .ip2(n5207), .op(n5210) );
  nand2_1 U5710 ( .ip1(n5208), .ip2(n5207), .op(n5209) );
  nand3_1 U5711 ( .ip1(n5211), .ip2(n5210), .ip3(n5209), .op(n5218) );
  fulladder U5712 ( .a(n5214), .b(n5213), .ci(n5212), .co(n5229), .s(n5220) );
  nand2_1 U5713 ( .ip1(n5218), .ip2(n5220), .op(n5223) );
  fulladder U5714 ( .a(n5217), .b(n5216), .ci(n5215), .co(n5219), .s(n5207) );
  nand2_1 U5715 ( .ip1(n5218), .ip2(n5219), .op(n5222) );
  nand2_1 U5716 ( .ip1(n5220), .ip2(n5219), .op(n5221) );
  nand3_1 U5717 ( .ip1(n5223), .ip2(n5222), .ip3(n5221), .op(n5230) );
  nor3_1 U5718 ( .ip1(n5228), .ip2(n5229), .ip3(n5230), .op(n5232) );
  fulladder U5719 ( .a(n5226), .b(n5225), .ci(n5224), .co(n5233), .s(n5227) );
  not_ab_or_c_or_d U5720 ( .ip1(n5230), .ip2(n5229), .ip3(n5228), .ip4(n5227), 
        .op(n5231) );
  or2_1 U5721 ( .ip1(n5232), .ip2(n5231), .op(n5236) );
  nor2_1 U5722 ( .ip1(n5234), .ip2(n5233), .op(n5235) );
  nor2_1 U5723 ( .ip1(n5236), .ip2(n5235), .op(n5842) );
  fulladder U5724 ( .a(n5239), .b(n5238), .ci(n5237), .co(n5841), .s(n5234) );
  inv_1 U5725 ( .ip(m1Inputs[37]), .op(n6749) );
  nor2_1 U5726 ( .ip1(n5552), .ip2(n6749), .op(n5269) );
  inv_1 U5727 ( .ip(m1Inputs[34]), .op(n5772) );
  nor2_1 U5728 ( .ip1(n6246), .ip2(n5772), .op(n5268) );
  inv_1 U5729 ( .ip(m1Inputs[32]), .op(n5295) );
  nor2_1 U5730 ( .ip1(n5295), .ip2(n7813), .op(n5267) );
  nand2_1 U5731 ( .ip1(n6280), .ip2(m1Inputs[36]), .op(n5774) );
  nor3_1 U5732 ( .ip1(n5414), .ip2(n5774), .ip3(n6749), .op(n5290) );
  or2_1 U5733 ( .ip1(n5774), .ip2(n5290), .op(n5242) );
  nand2_1 U5734 ( .ip1(n6248), .ip2(m1Inputs[37]), .op(n5240) );
  or2_1 U5735 ( .ip1(n5240), .ip2(n5290), .op(n5241) );
  nand2_1 U5736 ( .ip1(n5242), .ip2(n5241), .op(n5278) );
  inv_1 U5737 ( .ip(m1Inputs[33]), .op(n5309) );
  nor2_1 U5738 ( .ip1(n5309), .ip2(n7813), .op(n5264) );
  inv_1 U5739 ( .ip(m1Inputs[38]), .op(n6728) );
  nor2_1 U5740 ( .ip1(n5552), .ip2(n6728), .op(n5263) );
  nor2_1 U5741 ( .ip1(n5295), .ip2(n5669), .op(n5262) );
  and3_1 U5742 ( .ip1(n6248), .ip2(m1Inputs[38]), .ip3(n5287), .op(n5768) );
  inv_1 U5743 ( .ip(m1Inputs[36]), .op(n5735) );
  nand2_1 U5744 ( .ip1(n8001), .ip2(m1Inputs[39]), .op(n6694) );
  nor3_1 U5745 ( .ip1(n5552), .ip2(n5735), .ip3(n6694), .op(n5258) );
  nor2_1 U5746 ( .ip1(n6246), .ip2(n5735), .op(n5743) );
  or2_1 U5747 ( .ip1(m1Inputs[39]), .ip2(n5743), .op(n5244) );
  or2_1 U5748 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n5743), .op(n5243) );
  nand2_1 U5749 ( .ip1(n5244), .ip2(n5243), .op(n5257) );
  nand2_1 U5750 ( .ip1(n6280), .ip2(m1Inputs[37]), .op(n5259) );
  nor2_1 U5751 ( .ip1(n5257), .ip2(n5259), .op(n5245) );
  nor2_1 U5752 ( .ip1(n5258), .ip2(n5245), .op(n5758) );
  nand2_1 U5753 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[35]), .op(n5247)
         );
  nand2_1 U5754 ( .ip1(n8064), .ip2(m1Inputs[34]), .op(n5246) );
  xor2_1 U5755 ( .ip1(n5247), .ip2(n5246), .op(n5253) );
  inv_1 U5756 ( .ip(m1Inputs[35]), .op(n6691) );
  nand2_1 U5757 ( .ip1(m1Inputs[34]), .ip2(\STAGE_1/weightReg [4]), .op(n5281)
         );
  nor3_1 U5758 ( .ip1(n6691), .ip2(n7624), .ip3(n5281), .op(n5248) );
  or2_1 U5759 ( .ip1(n5253), .ip2(n5248), .op(n5250) );
  nor2_1 U5760 ( .ip1(n5295), .ip2(n7685), .op(n5252) );
  or2_1 U5761 ( .ip1(n5252), .ip2(n5248), .op(n5249) );
  nand2_1 U5762 ( .ip1(n5250), .ip2(n5249), .op(n5757) );
  nand2_1 U5763 ( .ip1(m1Inputs[34]), .ip2(\STAGE_1/weightReg [6]), .op(n5756)
         );
  inv_1 U5764 ( .ip(n5251), .op(n5765) );
  xnor2_1 U5765 ( .ip1(n5253), .ip2(n5252), .op(n5284) );
  nor3_1 U5766 ( .ip1(n5414), .ip2(n6691), .ip3(n5774), .op(n5274) );
  and2_1 U5767 ( .ip1(\STAGE_1/weightReg [3]), .ip2(n5274), .op(n5256) );
  nand2_1 U5768 ( .ip1(n8001), .ip2(m1Inputs[35]), .op(n5254) );
  mux2_1 U5769 ( .ip1(n5254), .ip2(n8001), .s(n5274), .op(n5280) );
  nor2_1 U5770 ( .ip1(n5281), .ip2(n5280), .op(n5255) );
  nor2_1 U5771 ( .ip1(n5256), .ip2(n5255), .op(n5283) );
  nor2_1 U5772 ( .ip1(n5258), .ip2(n5257), .op(n5260) );
  xor2_1 U5773 ( .ip1(n5260), .ip2(n5259), .op(n5282) );
  inv_1 U5774 ( .ip(n5261), .op(n5764) );
  nor2_1 U5775 ( .ip1(n5309), .ip2(n5669), .op(n5291) );
  fulladder U5776 ( .a(n5264), .b(n5263), .ci(n5262), .co(n5289), .s(n5277) );
  nand2_1 U5777 ( .ip1(m1Inputs[37]), .ip2(n8001), .op(n5266) );
  nor2_1 U5778 ( .ip1(n5735), .ip2(n5060), .op(n5265) );
  xor2_1 U5779 ( .ip1(n5266), .ip2(n5265), .op(n5745) );
  nand2_1 U5780 ( .ip1(m1Inputs[33]), .ip2(n7882), .op(n5744) );
  xor2_1 U5781 ( .ip1(n5745), .ip2(n5744), .op(n5755) );
  nor2_1 U5782 ( .ip1(n6691), .ip2(n7624), .op(n5740) );
  inv_1 U5783 ( .ip(m1Inputs[40]), .op(n6748) );
  nor2_1 U5784 ( .ip1(n5552), .ip2(n6748), .op(n5739) );
  nand2_1 U5785 ( .ip1(m1Inputs[32]), .ip2(\STAGE_1/weightReg [15]), .op(n5738) );
  inv_1 U5786 ( .ip(m1Inputs[39]), .op(n6717) );
  nor2_1 U5787 ( .ip1(n5414), .ip2(n6717), .op(n5742) );
  buf_1 U5788 ( .ip(n8175), .op(n7045) );
  nand2_1 U5789 ( .ip1(n7045), .ip2(column[32]), .op(n5760) );
  nor2_1 U5790 ( .ip1(n5593), .ip2(n6728), .op(n5741) );
  fulladder U5791 ( .a(n5269), .b(n5268), .ci(n5267), .co(n5279), .s(n5306) );
  nand2_1 U5792 ( .ip1(n6248), .ip2(m1Inputs[34]), .op(n5312) );
  nor3_1 U5793 ( .ip1(n5593), .ip2(n5312), .ip3(n6691), .op(n5303) );
  nor2_1 U5794 ( .ip1(n5593), .ip2(n6691), .op(n5270) );
  or2_1 U5795 ( .ip1(m1Inputs[36]), .ip2(n5270), .op(n5272) );
  or2_1 U5796 ( .ip1(\STAGE_1/weightReg [1]), .ip2(n5270), .op(n5271) );
  nand2_1 U5797 ( .ip1(n5272), .ip2(n5271), .op(n5273) );
  nor2_1 U5798 ( .ip1(n5274), .ip2(n5273), .op(n5276) );
  nor2_1 U5799 ( .ip1(n5309), .ip2(n5060), .op(n5275) );
  nor2_1 U5800 ( .ip1(n5552), .ip2(n5735), .op(n5298) );
  nor2_1 U5801 ( .ip1(n5295), .ip2(n5060), .op(n5297) );
  nor2_1 U5802 ( .ip1(n6246), .ip2(n5309), .op(n5296) );
  fulladder U5803 ( .a(n5303), .b(n5276), .ci(n5275), .co(n5294), .s(n5305) );
  fulladder U5804 ( .a(n5279), .b(n5278), .ci(n5277), .co(n5287), .s(n5293) );
  xor2_1 U5805 ( .ip1(n5281), .ip2(n5280), .op(n5292) );
  fulladder U5806 ( .a(n5284), .b(n5283), .ci(n5282), .co(n5261), .s(n5285) );
  inv_1 U5807 ( .ip(n5285), .op(n5354) );
  nor2_1 U5808 ( .ip1(n5414), .ip2(n6728), .op(n5286) );
  nor2_1 U5809 ( .ip1(n5287), .ip2(n5286), .op(n5288) );
  nor2_1 U5810 ( .ip1(n5768), .ip2(n5288), .op(n5353) );
  fulladder U5811 ( .a(n5291), .b(n5290), .ci(n5289), .co(n5763), .s(n5352) );
  fulladder U5812 ( .a(n5294), .b(n5293), .ci(n5292), .co(n5348), .s(n5345) );
  and2_1 U5813 ( .ip1(n5349), .ip2(n5348), .op(n5343) );
  nor3_1 U5814 ( .ip1(n5344), .ip2(n5345), .ip3(n5343), .op(n5347) );
  nor3_1 U5815 ( .ip1(n6246), .ip2(n5312), .ip3(n5295), .op(n5313) );
  fulladder U5816 ( .a(n5298), .b(n5297), .ci(n5296), .co(n5304), .s(n5308) );
  nor2_1 U5817 ( .ip1(n5414), .ip2(n6691), .op(n5299) );
  or2_1 U5818 ( .ip1(m1Inputs[34]), .ip2(n5299), .op(n5301) );
  or2_1 U5819 ( .ip1(\STAGE_1/weightReg [2]), .ip2(n5299), .op(n5300) );
  nand2_1 U5820 ( .ip1(n5301), .ip2(n5300), .op(n5302) );
  nor2_1 U5821 ( .ip1(n5303), .ip2(n5302), .op(n5307) );
  fulladder U5822 ( .a(n5306), .b(n5305), .ci(n5304), .co(n5344), .s(n5338) );
  nand2_1 U5823 ( .ip1(n5336), .ip2(n5338), .op(n5341) );
  fulladder U5824 ( .a(n5313), .b(n5308), .ci(n5307), .co(n5336), .s(n5330) );
  nand4_1 U5825 ( .ip1(\STAGE_1/weightReg [1]), .ip2(\STAGE_1/weightReg [2]), 
        .ip3(m1Inputs[32]), .ip4(m1Inputs[33]), .op(n5311) );
  not_ab_or_c_or_d U5826 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[32]), 
        .ip3(n5593), .ip4(n5309), .op(n5318) );
  nand3_1 U5827 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n5318), .ip3(m1Inputs[35]), .op(n5310) );
  nand2_1 U5828 ( .ip1(n5311), .ip2(n5310), .op(n5332) );
  nand2_1 U5829 ( .ip1(n5330), .ip2(n5332), .op(n5335) );
  or2_1 U5830 ( .ip1(n5312), .ip2(n5313), .op(n5316) );
  nand2_1 U5831 ( .ip1(n8001), .ip2(m1Inputs[32]), .op(n5314) );
  or2_1 U5832 ( .ip1(n5314), .ip2(n5313), .op(n5315) );
  nand2_1 U5833 ( .ip1(n5316), .ip2(n5315), .op(n5324) );
  nor2_1 U5834 ( .ip1(n5552), .ip2(n6691), .op(n5317) );
  xor2_1 U5835 ( .ip1(n5318), .ip2(n5317), .op(n5326) );
  nand2_1 U5836 ( .ip1(n5324), .ip2(n5326), .op(n5329) );
  nand2_1 U5837 ( .ip1(n6248), .ip2(m1Inputs[33]), .op(n5323) );
  nand2_1 U5838 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[32]), .op(n5322)
         );
  or2_1 U5839 ( .ip1(m1Inputs[32]), .ip2(m1Inputs[34]), .op(n5320) );
  or2_1 U5840 ( .ip1(n5593), .ip2(m1Inputs[34]), .op(n5319) );
  nand2_1 U5841 ( .ip1(n5320), .ip2(n5319), .op(n5321) );
  not_ab_or_c_or_d U5842 ( .ip1(n5323), .ip2(n5322), .ip3(n5321), .ip4(n5475), 
        .op(n5325) );
  nand2_1 U5843 ( .ip1(n5324), .ip2(n5325), .op(n5328) );
  nand2_1 U5844 ( .ip1(n5326), .ip2(n5325), .op(n5327) );
  nand3_1 U5845 ( .ip1(n5329), .ip2(n5328), .ip3(n5327), .op(n5331) );
  nand2_1 U5846 ( .ip1(n5330), .ip2(n5331), .op(n5334) );
  nand2_1 U5847 ( .ip1(n5332), .ip2(n5331), .op(n5333) );
  nand3_1 U5848 ( .ip1(n5335), .ip2(n5334), .ip3(n5333), .op(n5337) );
  nand2_1 U5849 ( .ip1(n5336), .ip2(n5337), .op(n5340) );
  nand2_1 U5850 ( .ip1(n5338), .ip2(n5337), .op(n5339) );
  nand3_1 U5851 ( .ip1(n5341), .ip2(n5340), .ip3(n5339), .op(n5342) );
  not_ab_or_c_or_d U5852 ( .ip1(n5345), .ip2(n5344), .ip3(n5343), .ip4(n5342), 
        .op(n5346) );
  or2_1 U5853 ( .ip1(n5347), .ip2(n5346), .op(n5351) );
  nor2_1 U5854 ( .ip1(n5349), .ip2(n5348), .op(n5350) );
  nor2_1 U5855 ( .ip1(n5351), .ip2(n5350), .op(n5770) );
  fulladder U5856 ( .a(n5354), .b(n5353), .ci(n5352), .co(n5769), .s(n5349) );
  inv_1 U5857 ( .ip(m1Inputs[21]), .op(n6557) );
  nor2_1 U5858 ( .ip1(n5552), .ip2(n6557), .op(n5412) );
  inv_1 U5859 ( .ip(m1Inputs[18]), .op(n5715) );
  nor2_1 U5860 ( .ip1(n6246), .ip2(n5715), .op(n5411) );
  inv_1 U5861 ( .ip(m1Inputs[16]), .op(n5413) );
  nor2_1 U5862 ( .ip1(n5413), .ip2(n7813), .op(n5410) );
  nand2_1 U5863 ( .ip1(n6280), .ip2(m1Inputs[20]), .op(n5717) );
  nor3_1 U5864 ( .ip1(n5414), .ip2(n5717), .ip3(n6557), .op(n5401) );
  or2_1 U5865 ( .ip1(n5717), .ip2(n5401), .op(n5357) );
  nand2_1 U5866 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[21]), .op(n5355)
         );
  or2_1 U5867 ( .ip1(n5355), .ip2(n5401), .op(n5356) );
  nand2_1 U5868 ( .ip1(n5357), .ip2(n5356), .op(n5389) );
  inv_1 U5869 ( .ip(m1Inputs[17]), .op(n5407) );
  nor2_1 U5870 ( .ip1(n5407), .ip2(n7813), .op(n5380) );
  inv_1 U5871 ( .ip(m1Inputs[22]), .op(n6544) );
  nor2_1 U5872 ( .ip1(n5475), .ip2(n6544), .op(n5379) );
  nor2_1 U5873 ( .ip1(n5413), .ip2(n5669), .op(n5378) );
  and3_1 U5874 ( .ip1(n6248), .ip2(m1Inputs[22]), .ip3(n5398), .op(n5696) );
  inv_1 U5875 ( .ip(m1Inputs[20]), .op(n6573) );
  nand2_1 U5876 ( .ip1(n8001), .ip2(m1Inputs[23]), .op(n6511) );
  nor3_1 U5877 ( .ip1(n5552), .ip2(n6573), .ip3(n6511), .op(n5374) );
  nor2_1 U5878 ( .ip1(n6246), .ip2(n6573), .op(n5358) );
  or2_1 U5879 ( .ip1(m1Inputs[23]), .ip2(n5358), .op(n5360) );
  or2_1 U5880 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n5358), .op(n5359) );
  nand2_1 U5881 ( .ip1(n5360), .ip2(n5359), .op(n5373) );
  nand2_1 U5882 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[21]), .op(n5375)
         );
  nor2_1 U5883 ( .ip1(n5373), .ip2(n5375), .op(n5361) );
  nor2_1 U5884 ( .ip1(n5374), .ip2(n5361), .op(n5686) );
  nand2_1 U5885 ( .ip1(n8064), .ip2(m1Inputs[18]), .op(n5363) );
  nand2_1 U5886 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[19]), .op(n5362)
         );
  xor2_1 U5887 ( .ip1(n5363), .ip2(n5362), .op(n5369) );
  inv_1 U5888 ( .ip(m1Inputs[19]), .op(n6512) );
  nand2_1 U5889 ( .ip1(m1Inputs[18]), .ip2(\STAGE_1/weightReg [4]), .op(n5392)
         );
  nor3_1 U5890 ( .ip1(n6512), .ip2(n7624), .ip3(n5392), .op(n5364) );
  or2_1 U5891 ( .ip1(n5369), .ip2(n5364), .op(n5366) );
  nor2_1 U5892 ( .ip1(n5413), .ip2(n7685), .op(n5368) );
  or2_1 U5893 ( .ip1(n5368), .ip2(n5364), .op(n5365) );
  nand2_1 U5894 ( .ip1(n5366), .ip2(n5365), .op(n5685) );
  nand2_1 U5895 ( .ip1(m1Inputs[18]), .ip2(\STAGE_1/weightReg [6]), .op(n5684)
         );
  inv_1 U5896 ( .ip(n5367), .op(n5693) );
  xnor2_1 U5897 ( .ip1(n5369), .ip2(n5368), .op(n5395) );
  nor3_1 U5898 ( .ip1(n5414), .ip2(n6512), .ip3(n5717), .op(n5387) );
  and2_1 U5899 ( .ip1(\STAGE_1/weightReg [3]), .ip2(n5387), .op(n5372) );
  nand2_1 U5900 ( .ip1(n8001), .ip2(m1Inputs[19]), .op(n5370) );
  mux2_1 U5901 ( .ip1(n5370), .ip2(n8001), .s(n5387), .op(n5391) );
  nor2_1 U5902 ( .ip1(n5392), .ip2(n5391), .op(n5371) );
  nor2_1 U5903 ( .ip1(n5372), .ip2(n5371), .op(n5394) );
  nor2_1 U5904 ( .ip1(n5374), .ip2(n5373), .op(n5376) );
  xor2_1 U5905 ( .ip1(n5376), .ip2(n5375), .op(n5393) );
  inv_1 U5906 ( .ip(n5377), .op(n5692) );
  nor2_1 U5907 ( .ip1(n5407), .ip2(n5669), .op(n5402) );
  fulladder U5908 ( .a(n5380), .b(n5379), .ci(n5378), .co(n5400), .s(n5388) );
  nand2_1 U5909 ( .ip1(m1Inputs[21]), .ip2(\STAGE_1/weightReg [3]), .op(n5382)
         );
  nor2_1 U5910 ( .ip1(n6573), .ip2(n5060), .op(n5381) );
  xor2_1 U5911 ( .ip1(n5382), .ip2(n5381), .op(n5665) );
  nand2_1 U5912 ( .ip1(m1Inputs[17]), .ip2(n7882), .op(n5664) );
  xor2_1 U5913 ( .ip1(n5665), .ip2(n5664), .op(n5683) );
  nor2_1 U5914 ( .ip1(n6512), .ip2(n7624), .op(n5678) );
  inv_1 U5915 ( .ip(m1Inputs[24]), .op(n6532) );
  nor2_1 U5916 ( .ip1(n5552), .ip2(n6532), .op(n5677) );
  nand2_1 U5917 ( .ip1(m1Inputs[16]), .ip2(\STAGE_1/weightReg [15]), .op(n5676) );
  inv_1 U5918 ( .ip(m1Inputs[23]), .op(n6533) );
  nor2_1 U5919 ( .ip1(n5414), .ip2(n6533), .op(n5680) );
  nand2_1 U5920 ( .ip1(n7045), .ip2(column[16]), .op(n5688) );
  nor2_1 U5921 ( .ip1(n5593), .ip2(n6544), .op(n5679) );
  nand2_1 U5922 ( .ip1(n6248), .ip2(m1Inputs[18]), .op(n5430) );
  nor3_1 U5923 ( .ip1(n5593), .ip2(n6512), .ip3(n5430), .op(n5419) );
  nor2_1 U5924 ( .ip1(n5593), .ip2(n6512), .op(n5383) );
  or2_1 U5925 ( .ip1(m1Inputs[20]), .ip2(n5383), .op(n5385) );
  or2_1 U5926 ( .ip1(\STAGE_1/weightReg [1]), .ip2(n5383), .op(n5384) );
  nand2_1 U5927 ( .ip1(n5385), .ip2(n5384), .op(n5386) );
  nor2_1 U5928 ( .ip1(n5387), .ip2(n5386), .op(n5409) );
  nor2_1 U5929 ( .ip1(n5407), .ip2(n5060), .op(n5408) );
  fulladder U5930 ( .a(n5390), .b(n5389), .ci(n5388), .co(n5398), .s(n5404) );
  xor2_1 U5931 ( .ip1(n5392), .ip2(n5391), .op(n5403) );
  fulladder U5932 ( .a(n5395), .b(n5394), .ci(n5393), .co(n5377), .s(n5396) );
  inv_1 U5933 ( .ip(n5396), .op(n5471) );
  nor2_1 U5934 ( .ip1(n5535), .ip2(n6544), .op(n5397) );
  nor2_1 U5935 ( .ip1(n5398), .ip2(n5397), .op(n5399) );
  nor2_1 U5936 ( .ip1(n5696), .ip2(n5399), .op(n5470) );
  fulladder U5937 ( .a(n5402), .b(n5401), .ci(n5400), .co(n5691), .s(n5469) );
  nand2_1 U5938 ( .ip1(n5460), .ip2(n5459), .op(n5468) );
  fulladder U5939 ( .a(n5405), .b(n5404), .ci(n5403), .co(n5460), .s(n5406) );
  inv_1 U5940 ( .ip(n5406), .op(n5466) );
  nor2_1 U5941 ( .ip1(n5552), .ip2(n6573), .op(n5422) );
  nor2_1 U5942 ( .ip1(n6246), .ip2(n5407), .op(n5421) );
  nor2_1 U5943 ( .ip1(n5413), .ip2(n5060), .op(n5420) );
  fulladder U5944 ( .a(n5419), .b(n5409), .ci(n5408), .co(n5405), .s(n5451) );
  fulladder U5945 ( .a(n5412), .b(n5411), .ci(n5410), .co(n5390), .s(n5450) );
  nor3_1 U5946 ( .ip1(n6246), .ip2(n5413), .ip3(n5430), .op(n5431) );
  nor2_1 U5947 ( .ip1(n5414), .ip2(n6512), .op(n5415) );
  or2_1 U5948 ( .ip1(m1Inputs[18]), .ip2(n5415), .op(n5417) );
  or2_1 U5949 ( .ip1(\STAGE_1/weightReg [2]), .ip2(n5415), .op(n5416) );
  nand2_1 U5950 ( .ip1(n5417), .ip2(n5416), .op(n5418) );
  nor2_1 U5951 ( .ip1(n5419), .ip2(n5418), .op(n5424) );
  fulladder U5952 ( .a(n5422), .b(n5421), .ci(n5420), .co(n5452), .s(n5423) );
  fulladder U5953 ( .a(n5431), .b(n5424), .ci(n5423), .co(n5453), .s(n5441) );
  nand2_1 U5954 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[19]), .op(n5427)
         );
  nand4_1 U5955 ( .ip1(\STAGE_1/weightReg [1]), .ip2(\STAGE_1/weightReg [2]), 
        .ip3(m1Inputs[16]), .ip4(m1Inputs[17]), .op(n5426) );
  and2_1 U5956 ( .ip1(n5427), .ip2(n5426), .op(n5425) );
  nand2_1 U5957 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[17]), .op(n5428)
         );
  nor2_1 U5958 ( .ip1(n5425), .ip2(n5428), .op(n5440) );
  nand2_1 U5959 ( .ip1(n5441), .ip2(n5440), .op(n5449) );
  xor2_1 U5960 ( .ip1(n5427), .ip2(n5426), .op(n5429) );
  xor2_1 U5961 ( .ip1(n5429), .ip2(n5428), .op(n5447) );
  or2_1 U5962 ( .ip1(n5430), .ip2(n5431), .op(n5434) );
  nand2_1 U5963 ( .ip1(n8001), .ip2(m1Inputs[16]), .op(n5432) );
  or2_1 U5964 ( .ip1(n5432), .ip2(n5431), .op(n5433) );
  nand2_1 U5965 ( .ip1(n5434), .ip2(n5433), .op(n5443) );
  nand2_1 U5966 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[16]), .op(n5439)
         );
  nand2_1 U5967 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[17]), .op(n5438)
         );
  or2_1 U5968 ( .ip1(m1Inputs[16]), .ip2(m1Inputs[18]), .op(n5436) );
  or2_1 U5969 ( .ip1(n5593), .ip2(m1Inputs[18]), .op(n5435) );
  nand2_1 U5970 ( .ip1(n5436), .ip2(n5435), .op(n5437) );
  not_ab_or_c_or_d U5971 ( .ip1(n5439), .ip2(n5438), .ip3(n5437), .ip4(n5552), 
        .op(n5442) );
  nand2_1 U5972 ( .ip1(n5443), .ip2(n5442), .op(n5446) );
  nor2_1 U5973 ( .ip1(n5441), .ip2(n5440), .op(n5445) );
  nor2_1 U5974 ( .ip1(n5443), .ip2(n5442), .op(n5444) );
  ab_or_c_or_d U5975 ( .ip1(n5447), .ip2(n5446), .ip3(n5445), .ip4(n5444), 
        .op(n5448) );
  nand2_1 U5976 ( .ip1(n5449), .ip2(n5448), .op(n5455) );
  nand2_1 U5977 ( .ip1(n5453), .ip2(n5455), .op(n5458) );
  fulladder U5978 ( .a(n5452), .b(n5451), .ci(n5450), .co(n5462), .s(n5454) );
  nand2_1 U5979 ( .ip1(n5453), .ip2(n5454), .op(n5457) );
  nand2_1 U5980 ( .ip1(n5455), .ip2(n5454), .op(n5456) );
  nand3_1 U5981 ( .ip1(n5458), .ip2(n5457), .ip3(n5456), .op(n5461) );
  nand2_1 U5982 ( .ip1(n5462), .ip2(n5461), .op(n5465) );
  nor2_1 U5983 ( .ip1(n5460), .ip2(n5459), .op(n5464) );
  nor2_1 U5984 ( .ip1(n5462), .ip2(n5461), .op(n5463) );
  ab_or_c_or_d U5985 ( .ip1(n5466), .ip2(n5465), .ip3(n5464), .ip4(n5463), 
        .op(n5467) );
  nand2_1 U5986 ( .ip1(n5468), .ip2(n5467), .op(n5698) );
  fulladder U5987 ( .a(n5471), .b(n5470), .ci(n5469), .co(n5697), .s(n5459) );
  inv_1 U5988 ( .ip(m1Inputs[5]), .op(n6375) );
  nor2_1 U5989 ( .ip1(n5475), .ip2(n6375), .op(n5517) );
  inv_1 U5990 ( .ip(m1Inputs[2]), .op(n5644) );
  nor2_1 U5991 ( .ip1(n6246), .ip2(n5644), .op(n5516) );
  inv_1 U5992 ( .ip(m1Inputs[0]), .op(n5534) );
  nor2_1 U5993 ( .ip1(n5534), .ip2(n7813), .op(n5515) );
  nand2_1 U5994 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[4]), .op(n5646)
         );
  nor3_1 U5995 ( .ip1(n5535), .ip2(n5646), .ip3(n6375), .op(n5526) );
  or2_1 U5996 ( .ip1(n5646), .ip2(n5526), .op(n5474) );
  nand2_1 U5997 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[5]), .op(n5472)
         );
  or2_1 U5998 ( .ip1(n5472), .ip2(n5526), .op(n5473) );
  nand2_1 U5999 ( .ip1(n5474), .ip2(n5473), .op(n5509) );
  inv_1 U6000 ( .ip(m1Inputs[1]), .op(n5551) );
  nor2_1 U6001 ( .ip1(n5551), .ip2(n7813), .op(n5499) );
  inv_1 U6002 ( .ip(m1Inputs[6]), .op(n6362) );
  nor2_1 U6003 ( .ip1(n5552), .ip2(n6362), .op(n5498) );
  nor2_1 U6004 ( .ip1(n5534), .ip2(n5669), .op(n5497) );
  and3_1 U6005 ( .ip1(n6248), .ip2(m1Inputs[6]), .ip3(n5523), .op(n5625) );
  nand2_1 U6006 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[4]), .op(n5476)
         );
  inv_1 U6007 ( .ip(m1Inputs[4]), .op(n6391) );
  nand2_1 U6008 ( .ip1(n8001), .ip2(m1Inputs[7]), .op(n6329) );
  nor3_1 U6009 ( .ip1(n5475), .ip2(n6391), .ip3(n6329), .op(n5480) );
  or2_1 U6010 ( .ip1(n5476), .ip2(n5480), .op(n5479) );
  nand2_1 U6011 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[7]), .op(n5477)
         );
  or2_1 U6012 ( .ip1(n5477), .ip2(n5480), .op(n5478) );
  nand2_1 U6013 ( .ip1(n5479), .ip2(n5478), .op(n5495) );
  or2_1 U6014 ( .ip1(n5495), .ip2(n5480), .op(n5482) );
  nor2_1 U6015 ( .ip1(n5593), .ip2(n6375), .op(n5494) );
  or2_1 U6016 ( .ip1(n5494), .ip2(n5480), .op(n5481) );
  nand2_1 U6017 ( .ip1(n5482), .ip2(n5481), .op(n5615) );
  nand2_1 U6018 ( .ip1(n8064), .ip2(m1Inputs[2]), .op(n5484) );
  nand2_1 U6019 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[3]), .op(n5483)
         );
  xor2_1 U6020 ( .ip1(n5484), .ip2(n5483), .op(n5490) );
  inv_1 U6021 ( .ip(m1Inputs[3]), .op(n6330) );
  nand2_1 U6022 ( .ip1(m1Inputs[2]), .ip2(\STAGE_1/weightReg [4]), .op(n5512)
         );
  nor3_1 U6023 ( .ip1(n6330), .ip2(n7813), .ip3(n5512), .op(n5485) );
  or2_1 U6024 ( .ip1(n5490), .ip2(n5485), .op(n5487) );
  nor2_1 U6025 ( .ip1(n5534), .ip2(n7685), .op(n5489) );
  or2_1 U6026 ( .ip1(n5489), .ip2(n5485), .op(n5486) );
  nand2_1 U6027 ( .ip1(n5487), .ip2(n5486), .op(n5614) );
  nand2_1 U6028 ( .ip1(m1Inputs[2]), .ip2(n8037), .op(n5613) );
  inv_1 U6029 ( .ip(n5488), .op(n5622) );
  xnor2_1 U6030 ( .ip1(n5490), .ip2(n5489), .op(n5520) );
  nor3_1 U6031 ( .ip1(n5535), .ip2(n6330), .ip3(n5646), .op(n5507) );
  and2_1 U6032 ( .ip1(\STAGE_1/weightReg [3]), .ip2(n5507), .op(n5493) );
  nand2_1 U6033 ( .ip1(n8001), .ip2(m1Inputs[3]), .op(n5491) );
  mux2_1 U6034 ( .ip1(n5491), .ip2(\STAGE_1/weightReg [3]), .s(n5507), .op(
        n5511) );
  nor2_1 U6035 ( .ip1(n5512), .ip2(n5511), .op(n5492) );
  nor2_1 U6036 ( .ip1(n5493), .ip2(n5492), .op(n5519) );
  xnor2_1 U6037 ( .ip1(n5495), .ip2(n5494), .op(n5518) );
  inv_1 U6038 ( .ip(n5496), .op(n5621) );
  nor2_1 U6039 ( .ip1(n5551), .ip2(n5669), .op(n5527) );
  fulladder U6040 ( .a(n5499), .b(n5498), .ci(n5497), .co(n5525), .s(n5508) );
  nor2_1 U6041 ( .ip1(n6375), .ip2(n5500), .op(n5502) );
  nand2_1 U6042 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[4]), .op(n5501)
         );
  xor2_1 U6043 ( .ip1(n5502), .ip2(n5501), .op(n5602) );
  nand2_1 U6044 ( .ip1(m1Inputs[1]), .ip2(n7882), .op(n5601) );
  xor2_1 U6045 ( .ip1(n5602), .ip2(n5601), .op(n5612) );
  nor2_1 U6046 ( .ip1(n6330), .ip2(n7813), .op(n5598) );
  inv_1 U6047 ( .ip(m1Inputs[8]), .op(n6350) );
  nor2_1 U6048 ( .ip1(n5552), .ip2(n6350), .op(n5597) );
  nand2_1 U6049 ( .ip1(m1Inputs[0]), .ip2(\STAGE_1/weightReg [15]), .op(n5596)
         );
  inv_1 U6050 ( .ip(m1Inputs[7]), .op(n6351) );
  nor2_1 U6051 ( .ip1(n5535), .ip2(n6351), .op(n5600) );
  nand2_1 U6052 ( .ip1(n7045), .ip2(column[0]), .op(n5617) );
  nor2_1 U6053 ( .ip1(n5593), .ip2(n6362), .op(n5599) );
  nand2_1 U6054 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[2]), .op(n5546)
         );
  nor3_1 U6055 ( .ip1(n5593), .ip2(n6330), .ip3(n5546), .op(n5540) );
  nor2_1 U6056 ( .ip1(n5593), .ip2(n6330), .op(n5503) );
  or2_1 U6057 ( .ip1(m1Inputs[4]), .ip2(n5503), .op(n5505) );
  or2_1 U6058 ( .ip1(\STAGE_1/weightReg [1]), .ip2(n5503), .op(n5504) );
  nand2_1 U6059 ( .ip1(n5505), .ip2(n5504), .op(n5506) );
  nor2_1 U6060 ( .ip1(n5507), .ip2(n5506), .op(n5514) );
  nor2_1 U6061 ( .ip1(n5551), .ip2(n5060), .op(n5513) );
  fulladder U6062 ( .a(n5510), .b(n5509), .ci(n5508), .co(n5523), .s(n5529) );
  xor2_1 U6063 ( .ip1(n5512), .ip2(n5511), .op(n5528) );
  fulladder U6064 ( .a(n5540), .b(n5514), .ci(n5513), .co(n5530), .s(n5543) );
  nor2_1 U6065 ( .ip1(n5552), .ip2(n6391), .op(n5533) );
  nor2_1 U6066 ( .ip1(n6246), .ip2(n5551), .op(n5532) );
  nor2_1 U6067 ( .ip1(n5534), .ip2(n5060), .op(n5531) );
  fulladder U6068 ( .a(n5517), .b(n5516), .ci(n5515), .co(n5510), .s(n5541) );
  fulladder U6069 ( .a(n5520), .b(n5519), .ci(n5518), .co(n5496), .s(n5521) );
  inv_1 U6070 ( .ip(n5521), .op(n5592) );
  nor2_1 U6071 ( .ip1(n5535), .ip2(n6362), .op(n5522) );
  nor2_1 U6072 ( .ip1(n5523), .ip2(n5522), .op(n5524) );
  nor2_1 U6073 ( .ip1(n5625), .ip2(n5524), .op(n5591) );
  fulladder U6074 ( .a(n5527), .b(n5526), .ci(n5525), .co(n5620), .s(n5590) );
  fulladder U6075 ( .a(n5530), .b(n5529), .ci(n5528), .co(n5586), .s(n5582) );
  and2_1 U6076 ( .ip1(n5587), .ip2(n5586), .op(n5581) );
  nor3_1 U6077 ( .ip1(n5582), .ip2(n5583), .ip3(n5581), .op(n5585) );
  fulladder U6078 ( .a(n5533), .b(n5532), .ci(n5531), .co(n5542), .s(n5545) );
  nor3_1 U6079 ( .ip1(n6246), .ip2(n5534), .ip3(n5546), .op(n5547) );
  nor2_1 U6080 ( .ip1(n5535), .ip2(n6330), .op(n5536) );
  or2_1 U6081 ( .ip1(m1Inputs[2]), .ip2(n5536), .op(n5538) );
  or2_1 U6082 ( .ip1(\STAGE_1/weightReg [2]), .ip2(n5536), .op(n5537) );
  nand2_1 U6083 ( .ip1(n5538), .ip2(n5537), .op(n5539) );
  nor2_1 U6084 ( .ip1(n5540), .ip2(n5539), .op(n5544) );
  fulladder U6085 ( .a(n5543), .b(n5542), .ci(n5541), .co(n5583), .s(n5576) );
  nand2_1 U6086 ( .ip1(n5574), .ip2(n5576), .op(n5579) );
  fulladder U6087 ( .a(n5545), .b(n5547), .ci(n5544), .co(n5574), .s(n5568) );
  or2_1 U6088 ( .ip1(n5546), .ip2(n5547), .op(n5550) );
  nand2_1 U6089 ( .ip1(n8001), .ip2(m1Inputs[0]), .op(n5548) );
  or2_1 U6090 ( .ip1(n5548), .ip2(n5547), .op(n5549) );
  nand2_1 U6091 ( .ip1(n5550), .ip2(n5549), .op(n5559) );
  not_ab_or_c_or_d U6092 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[0]), 
        .ip3(n5593), .ip4(n5551), .op(n5565) );
  nor2_1 U6093 ( .ip1(n5552), .ip2(n6330), .op(n5553) );
  xor2_1 U6094 ( .ip1(n5565), .ip2(n5553), .op(n5561) );
  nand2_1 U6095 ( .ip1(n5559), .ip2(n5561), .op(n5564) );
  nand2_1 U6096 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[0]), .op(n5558)
         );
  nand2_1 U6097 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[1]), .op(n5557)
         );
  or2_1 U6098 ( .ip1(m1Inputs[0]), .ip2(m1Inputs[2]), .op(n5555) );
  or2_1 U6099 ( .ip1(n5593), .ip2(m1Inputs[2]), .op(n5554) );
  nand2_1 U6100 ( .ip1(n5555), .ip2(n5554), .op(n5556) );
  not_ab_or_c_or_d U6101 ( .ip1(n5558), .ip2(n5557), .ip3(n5556), .ip4(n5552), 
        .op(n5560) );
  nand2_1 U6102 ( .ip1(n5559), .ip2(n5560), .op(n5563) );
  nand2_1 U6103 ( .ip1(n5561), .ip2(n5560), .op(n5562) );
  nand3_1 U6104 ( .ip1(n5564), .ip2(n5563), .ip3(n5562), .op(n5570) );
  nand2_1 U6105 ( .ip1(n5568), .ip2(n5570), .op(n5573) );
  nand4_1 U6106 ( .ip1(n6248), .ip2(\STAGE_1/weightReg [2]), .ip3(m1Inputs[0]), 
        .ip4(m1Inputs[1]), .op(n5567) );
  nand3_1 U6107 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n5565), .ip3(m1Inputs[3]), 
        .op(n5566) );
  nand2_1 U6108 ( .ip1(n5567), .ip2(n5566), .op(n5569) );
  nand2_1 U6109 ( .ip1(n5568), .ip2(n5569), .op(n5572) );
  nand2_1 U6110 ( .ip1(n5570), .ip2(n5569), .op(n5571) );
  nand3_1 U6111 ( .ip1(n5573), .ip2(n5572), .ip3(n5571), .op(n5575) );
  nand2_1 U6112 ( .ip1(n5574), .ip2(n5575), .op(n5578) );
  nand2_1 U6113 ( .ip1(n5576), .ip2(n5575), .op(n5577) );
  nand3_1 U6114 ( .ip1(n5579), .ip2(n5578), .ip3(n5577), .op(n5580) );
  not_ab_or_c_or_d U6115 ( .ip1(n5583), .ip2(n5582), .ip3(n5581), .ip4(n5580), 
        .op(n5584) );
  or2_1 U6116 ( .ip1(n5585), .ip2(n5584), .op(n5589) );
  nor2_1 U6117 ( .ip1(n5587), .ip2(n5586), .op(n5588) );
  nor2_1 U6118 ( .ip1(n5589), .ip2(n5588), .op(n5627) );
  fulladder U6119 ( .a(n5592), .b(n5591), .ci(n5590), .co(n5626), .s(n5587) );
  nor2_1 U6120 ( .ip1(n6351), .ip2(n5593), .op(n5595) );
  nand2_1 U6121 ( .ip1(m1Inputs[4]), .ip2(\STAGE_1/weightReg [5]), .op(n5594)
         );
  xor2_1 U6122 ( .ip1(n5595), .ip2(n5594), .op(n5648) );
  nand2_1 U6123 ( .ip1(n7045), .ip2(column[1]), .op(n5647) );
  xor2_1 U6124 ( .ip1(n5648), .ip2(n5647), .op(n5654) );
  fulladder U6125 ( .a(n5598), .b(n5597), .ci(n5596), .co(n5653), .s(n5611) );
  fulladder U6126 ( .a(n5600), .b(n5617), .ci(n5599), .co(n5652), .s(n5610) );
  nor2_1 U6127 ( .ip1(n6375), .ip2(n5060), .op(n5636) );
  and3_1 U6128 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[4]), .ip3(n5636), 
        .op(n5604) );
  nor2_1 U6129 ( .ip1(n5602), .ip2(n5601), .op(n5603) );
  nor2_1 U6130 ( .ip1(n5604), .ip2(n5603), .op(n5642) );
  nor2_1 U6131 ( .ip1(n6246), .ip2(n6362), .op(n5637) );
  nand2_1 U6132 ( .ip1(m1Inputs[1]), .ip2(\STAGE_1/weightReg [15]), .op(n5635)
         );
  inv_1 U6133 ( .ip(n5605), .op(n5641) );
  nand2_1 U6134 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[3]), .op(n5607)
         );
  nand2_1 U6135 ( .ip1(m1Inputs[8]), .ip2(n6248), .op(n5606) );
  xor2_1 U6136 ( .ip1(n5607), .ip2(n5606), .op(n5632) );
  nand2_1 U6137 ( .ip1(m1Inputs[2]), .ip2(n7882), .op(n5608) );
  xor2_1 U6138 ( .ip1(n5632), .ip2(n5608), .op(n5640) );
  inv_1 U6139 ( .ip(n5609), .op(n5656) );
  fulladder U6140 ( .a(n5612), .b(n5611), .ci(n5610), .co(n5655), .s(n5623) );
  fulladder U6141 ( .a(n5615), .b(n5614), .ci(n5613), .co(n5616), .s(n5488) );
  nor2_1 U6142 ( .ip1(n5616), .ip2(n5617), .op(n5639) );
  or2_1 U6143 ( .ip1(n5616), .ip2(n5639), .op(n5619) );
  or2_1 U6144 ( .ip1(n5617), .ip2(n5639), .op(n5618) );
  nand2_1 U6145 ( .ip1(n5619), .ip2(n5618), .op(n5662) );
  fulladder U6146 ( .a(n5622), .b(n5621), .ci(n5620), .co(n5661), .s(n5624) );
  fulladder U6147 ( .a(n5625), .b(n5624), .ci(n5623), .co(n5659), .s(n5628) );
  fulladder U6148 ( .a(n5628), .b(n5627), .ci(n5626), .co(n5658), .s(
        \STAGE_1/M1/sum [0]) );
  nand2_1 U6149 ( .ip1(m1Inputs[6]), .ip2(\STAGE_1/weightReg [4]), .op(n5630)
         );
  nand2_1 U6150 ( .ip1(\STAGE_1/weightReg [5]), .ip2(m1Inputs[5]), .op(n5629)
         );
  nand2_1 U6151 ( .ip1(n5630), .ip2(n5629), .op(n5631) );
  nand3_1 U6152 ( .ip1(m1Inputs[6]), .ip2(\STAGE_1/weightReg [5]), .ip3(n5636), 
        .op(n6315) );
  nand2_1 U6153 ( .ip1(n5631), .ip2(n6315), .op(n6317) );
  nand2_1 U6154 ( .ip1(n7045), .ip2(column[2]), .op(n6316) );
  xor2_1 U6155 ( .ip1(n6317), .ip2(n6316), .op(n6334) );
  nand3_1 U6156 ( .ip1(m1Inputs[2]), .ip2(n5632), .ip3(\STAGE_1/weightReg [7]), 
        .op(n5634) );
  nand4_1 U6157 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[3]), .ip3(
        m1Inputs[8]), .ip4(\STAGE_1/weightReg [6]), .op(n5633) );
  nand2_1 U6158 ( .ip1(n5634), .ip2(n5633), .op(n6333) );
  fulladder U6159 ( .a(n5637), .b(n5636), .ci(n5635), .co(n6332), .s(n5605) );
  inv_1 U6160 ( .ip(n5638), .op(n6342) );
  inv_1 U6161 ( .ip(n5639), .op(n6341) );
  fulladder U6162 ( .a(n5642), .b(n5641), .ci(n5640), .co(n6340), .s(n5609) );
  inv_1 U6163 ( .ip(n5643), .op(n6346) );
  nor2_1 U6164 ( .ip1(n5644), .ip2(n8029), .op(n6322) );
  nand2_1 U6165 ( .ip1(n6280), .ip2(m1Inputs[8]), .op(n6321) );
  nand2_1 U6166 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[4]), .op(n6320)
         );
  inv_1 U6167 ( .ip(n5645), .op(n6338) );
  nor3_1 U6168 ( .ip1(n6351), .ip2(n7813), .ip3(n5646), .op(n5650) );
  nor2_1 U6169 ( .ip1(n5648), .ip2(n5647), .op(n5649) );
  nor2_1 U6170 ( .ip1(n5650), .ip2(n5649), .op(n6328) );
  nand2_1 U6171 ( .ip1(m1Inputs[3]), .ip2(\STAGE_1/weightReg [7]), .op(n6327)
         );
  inv_1 U6172 ( .ip(n5651), .op(n6337) );
  fulladder U6173 ( .a(n5654), .b(n5653), .ci(n5652), .co(n6336), .s(n5657) );
  fulladder U6174 ( .a(n5657), .b(n5656), .ci(n5655), .co(n6344), .s(n5663) );
  fulladder U6175 ( .a(n5660), .b(n5659), .ci(n5658), .co(n6348), .s(
        \STAGE_1/M1/sum [1]) );
  fulladder U6176 ( .a(n5663), .b(n5662), .ci(n5661), .co(n6347), .s(n5660) );
  nor2_1 U6177 ( .ip1(n5060), .ip2(n6557), .op(n5707) );
  and3_1 U6178 ( .ip1(n8001), .ip2(m1Inputs[20]), .ip3(n5707), .op(n5667) );
  nor2_1 U6179 ( .ip1(n5665), .ip2(n5664), .op(n5666) );
  nor2_1 U6180 ( .ip1(n5667), .ip2(n5666), .op(n5713) );
  nor2_1 U6181 ( .ip1(n6246), .ip2(n6544), .op(n5708) );
  nand2_1 U6182 ( .ip1(m1Inputs[17]), .ip2(\STAGE_1/weightReg [15]), .op(n5706) );
  inv_1 U6183 ( .ip(n5668), .op(n5712) );
  nand2_1 U6184 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[19]), .op(n5671)
         );
  nand2_1 U6185 ( .ip1(m1Inputs[24]), .ip2(\STAGE_1/weightReg [1]), .op(n5670)
         );
  xor2_1 U6186 ( .ip1(n5671), .ip2(n5670), .op(n5703) );
  nand2_1 U6187 ( .ip1(m1Inputs[18]), .ip2(n7882), .op(n5672) );
  xor2_1 U6188 ( .ip1(n5703), .ip2(n5672), .op(n5711) );
  inv_1 U6189 ( .ip(n5673), .op(n5728) );
  nand2_1 U6190 ( .ip1(m1Inputs[23]), .ip2(\STAGE_1/weightReg [2]), .op(n5675)
         );
  nor2_1 U6191 ( .ip1(n7813), .ip2(n6573), .op(n5674) );
  xor2_1 U6192 ( .ip1(n5675), .ip2(n5674), .op(n5719) );
  nand2_1 U6193 ( .ip1(n7045), .ip2(column[17]), .op(n5718) );
  xor2_1 U6194 ( .ip1(n5719), .ip2(n5718), .op(n5725) );
  fulladder U6195 ( .a(n5678), .b(n5677), .ci(n5676), .co(n5724), .s(n5682) );
  fulladder U6196 ( .a(n5680), .b(n5688), .ci(n5679), .co(n5723), .s(n5681) );
  fulladder U6197 ( .a(n5683), .b(n5682), .ci(n5681), .co(n5726), .s(n5694) );
  fulladder U6198 ( .a(n5686), .b(n5685), .ci(n5684), .co(n5687), .s(n5367) );
  nor2_1 U6199 ( .ip1(n5687), .ip2(n5688), .op(n5710) );
  or2_1 U6200 ( .ip1(n5687), .ip2(n5710), .op(n5690) );
  or2_1 U6201 ( .ip1(n5688), .ip2(n5710), .op(n5689) );
  nand2_1 U6202 ( .ip1(n5690), .ip2(n5689), .op(n5733) );
  fulladder U6203 ( .a(n5693), .b(n5692), .ci(n5691), .co(n5732), .s(n5695) );
  fulladder U6204 ( .a(n5696), .b(n5695), .ci(n5694), .co(n5730), .s(n5699) );
  fulladder U6205 ( .a(n5699), .b(n5698), .ci(n5697), .co(n5729), .s(
        \STAGE_1/M2/sum [0]) );
  nand2_1 U6206 ( .ip1(m1Inputs[22]), .ip2(\STAGE_1/weightReg [4]), .op(n5701)
         );
  nand2_1 U6207 ( .ip1(n8064), .ip2(m1Inputs[21]), .op(n5700) );
  nand2_1 U6208 ( .ip1(n5701), .ip2(n5700), .op(n5702) );
  nand3_1 U6209 ( .ip1(\STAGE_1/weightReg [5]), .ip2(m1Inputs[22]), .ip3(n5707), .op(n6497) );
  nand2_1 U6210 ( .ip1(n5702), .ip2(n6497), .op(n6499) );
  nand2_1 U6211 ( .ip1(n7045), .ip2(column[18]), .op(n6498) );
  xor2_1 U6212 ( .ip1(n6499), .ip2(n6498), .op(n6516) );
  nand3_1 U6213 ( .ip1(m1Inputs[18]), .ip2(n5703), .ip3(\STAGE_1/weightReg [7]), .op(n5705) );
  nand4_1 U6214 ( .ip1(n6248), .ip2(m1Inputs[19]), .ip3(\STAGE_1/weightReg [6]), .ip4(m1Inputs[24]), .op(n5704) );
  nand2_1 U6215 ( .ip1(n5705), .ip2(n5704), .op(n6515) );
  fulladder U6216 ( .a(n5708), .b(n5707), .ci(n5706), .co(n6514), .s(n5668) );
  inv_1 U6217 ( .ip(n5709), .op(n6524) );
  inv_1 U6218 ( .ip(n5710), .op(n6523) );
  fulladder U6219 ( .a(n5713), .b(n5712), .ci(n5711), .co(n6522), .s(n5673) );
  inv_1 U6220 ( .ip(n5714), .op(n6528) );
  nor2_1 U6221 ( .ip1(n5715), .ip2(n8029), .op(n6504) );
  nand2_1 U6222 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[24]), .op(n6503)
         );
  nand2_1 U6223 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[20]), .op(n6502)
         );
  inv_1 U6224 ( .ip(n5716), .op(n6520) );
  nor3_1 U6225 ( .ip1(n7813), .ip2(n6533), .ip3(n5717), .op(n5721) );
  nor2_1 U6226 ( .ip1(n5719), .ip2(n5718), .op(n5720) );
  nor2_1 U6227 ( .ip1(n5721), .ip2(n5720), .op(n6510) );
  nand2_1 U6228 ( .ip1(m1Inputs[19]), .ip2(n7882), .op(n6509) );
  inv_1 U6229 ( .ip(n5722), .op(n6519) );
  fulladder U6230 ( .a(n5725), .b(n5724), .ci(n5723), .co(n6518), .s(n5727) );
  fulladder U6231 ( .a(n5728), .b(n5727), .ci(n5726), .co(n6526), .s(n5734) );
  fulladder U6232 ( .a(n5731), .b(n5730), .ci(n5729), .co(n6530), .s(
        \STAGE_1/M2/sum [1]) );
  fulladder U6233 ( .a(n5734), .b(n5733), .ci(n5732), .co(n6529), .s(n5731) );
  nand2_1 U6234 ( .ip1(m1Inputs[39]), .ip2(\STAGE_1/weightReg [2]), .op(n5737)
         );
  nor2_1 U6235 ( .ip1(n7813), .ip2(n5735), .op(n5736) );
  xor2_1 U6236 ( .ip1(n5737), .ip2(n5736), .op(n5776) );
  nand2_1 U6237 ( .ip1(n7045), .ip2(column[33]), .op(n5775) );
  xor2_1 U6238 ( .ip1(n5776), .ip2(n5775), .op(n5782) );
  fulladder U6239 ( .a(n5740), .b(n5739), .ci(n5738), .co(n5781), .s(n5754) );
  fulladder U6240 ( .a(n5742), .b(n5760), .ci(n5741), .co(n5780), .s(n5753) );
  nor2_1 U6241 ( .ip1(n5060), .ip2(n6749), .op(n5791) );
  and2_1 U6242 ( .ip1(n5791), .ip2(n5743), .op(n5747) );
  nor2_1 U6243 ( .ip1(n5745), .ip2(n5744), .op(n5746) );
  nor2_1 U6244 ( .ip1(n5747), .ip2(n5746), .op(n5797) );
  nor2_1 U6245 ( .ip1(n6246), .ip2(n6728), .op(n5792) );
  nand2_1 U6246 ( .ip1(m1Inputs[33]), .ip2(\STAGE_1/weightReg [15]), .op(n5790) );
  inv_1 U6247 ( .ip(n5748), .op(n5796) );
  nand2_1 U6248 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[35]), .op(n5750)
         );
  nand2_1 U6249 ( .ip1(m1Inputs[40]), .ip2(n6248), .op(n5749) );
  xor2_1 U6250 ( .ip1(n5750), .ip2(n5749), .op(n5787) );
  nand2_1 U6251 ( .ip1(m1Inputs[34]), .ip2(n7882), .op(n5751) );
  xor2_1 U6252 ( .ip1(n5787), .ip2(n5751), .op(n5795) );
  inv_1 U6253 ( .ip(n5752), .op(n5800) );
  fulladder U6254 ( .a(n5755), .b(n5754), .ci(n5753), .co(n5799), .s(n5766) );
  fulladder U6255 ( .a(n5758), .b(n5757), .ci(n5756), .co(n5759), .s(n5251) );
  nor2_1 U6256 ( .ip1(n5759), .ip2(n5760), .op(n5794) );
  or2_1 U6257 ( .ip1(n5759), .ip2(n5794), .op(n5762) );
  or2_1 U6258 ( .ip1(n5760), .ip2(n5794), .op(n5761) );
  nand2_1 U6259 ( .ip1(n5762), .ip2(n5761), .op(n5806) );
  fulladder U6260 ( .a(n5765), .b(n5764), .ci(n5763), .co(n5805), .s(n5767) );
  fulladder U6261 ( .a(n5768), .b(n5767), .ci(n5766), .co(n5803), .s(n5771) );
  fulladder U6262 ( .a(n5771), .b(n5770), .ci(n5769), .co(n5802), .s(
        \STAGE_1/M3/sum [0]) );
  nor2_1 U6263 ( .ip1(n5772), .ip2(n8029), .op(n6689) );
  nand2_1 U6264 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[40]), .op(n6688)
         );
  nand2_1 U6265 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[36]), .op(n6687)
         );
  inv_1 U6266 ( .ip(n5773), .op(n6705) );
  nand2_1 U6267 ( .ip1(n8064), .ip2(m1Inputs[39]), .op(n6743) );
  nor2_1 U6268 ( .ip1(n6743), .ip2(n5774), .op(n5778) );
  nor2_1 U6269 ( .ip1(n5776), .ip2(n5775), .op(n5777) );
  nor2_1 U6270 ( .ip1(n5778), .ip2(n5777), .op(n6693) );
  nand2_1 U6271 ( .ip1(m1Inputs[35]), .ip2(n7882), .op(n6692) );
  inv_1 U6272 ( .ip(n5779), .op(n6704) );
  fulladder U6273 ( .a(n5782), .b(n5781), .ci(n5780), .co(n6703), .s(n5801) );
  nand2_1 U6274 ( .ip1(n8064), .ip2(m1Inputs[38]), .op(n6740) );
  nor3_1 U6275 ( .ip1(n5060), .ip2(n6740), .ip3(n6749), .op(n6686) );
  nor2_1 U6276 ( .ip1(n7813), .ip2(n6749), .op(n5783) );
  or2_1 U6277 ( .ip1(m1Inputs[38]), .ip2(n5783), .op(n5785) );
  or2_1 U6278 ( .ip1(n8078), .ip2(n5783), .op(n5784) );
  nand2_1 U6279 ( .ip1(n5785), .ip2(n5784), .op(n6684) );
  or2_1 U6280 ( .ip1(n6686), .ip2(n6684), .op(n5786) );
  nand2_1 U6281 ( .ip1(n7045), .ip2(column[34]), .op(n6683) );
  xor2_1 U6282 ( .ip1(n5786), .ip2(n6683), .op(n6701) );
  nand3_1 U6283 ( .ip1(m1Inputs[34]), .ip2(n5787), .ip3(\STAGE_1/weightReg [7]), .op(n5789) );
  nand4_1 U6284 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[35]), .ip3(
        \STAGE_1/weightReg [6]), .ip4(m1Inputs[40]), .op(n5788) );
  nand2_1 U6285 ( .ip1(n5789), .ip2(n5788), .op(n6700) );
  fulladder U6286 ( .a(n5792), .b(n5791), .ci(n5790), .co(n6699), .s(n5748) );
  inv_1 U6287 ( .ip(n5793), .op(n6709) );
  inv_1 U6288 ( .ip(n5794), .op(n6708) );
  fulladder U6289 ( .a(n5797), .b(n5796), .ci(n5795), .co(n6707), .s(n5752) );
  inv_1 U6290 ( .ip(n5798), .op(n6712) );
  fulladder U6291 ( .a(n5801), .b(n5800), .ci(n5799), .co(n6711), .s(n5807) );
  fulladder U6292 ( .a(n5804), .b(n5803), .ci(n5802), .co(n6715), .s(
        \STAGE_1/M3/sum [1]) );
  fulladder U6293 ( .a(n5807), .b(n5806), .ci(n5805), .co(n6714), .s(n5804) );
  nand2_1 U6294 ( .ip1(m1Inputs[55]), .ip2(\STAGE_1/weightReg [2]), .op(n5809)
         );
  nor2_1 U6295 ( .ip1(n7624), .ip2(n6947), .op(n5808) );
  xor2_1 U6296 ( .ip1(n5809), .ip2(n5808), .op(n5848) );
  nand2_1 U6297 ( .ip1(n8009), .ip2(column[49]), .op(n5847) );
  xor2_1 U6298 ( .ip1(n5848), .ip2(n5847), .op(n5854) );
  fulladder U6299 ( .a(n5812), .b(n5811), .ci(n5810), .co(n5853), .s(n5826) );
  fulladder U6300 ( .a(n5814), .b(n5832), .ci(n5813), .co(n5852), .s(n5825) );
  nor2_1 U6301 ( .ip1(n5060), .ip2(n6931), .op(n5862) );
  and2_1 U6302 ( .ip1(n5862), .ip2(n5815), .op(n5819) );
  nor2_1 U6303 ( .ip1(n5817), .ip2(n5816), .op(n5818) );
  nor2_1 U6304 ( .ip1(n5819), .ip2(n5818), .op(n5868) );
  nor2_1 U6305 ( .ip1(n6246), .ip2(n6918), .op(n5863) );
  nand2_1 U6306 ( .ip1(m1Inputs[49]), .ip2(\STAGE_1/weightReg [15]), .op(n5861) );
  inv_1 U6307 ( .ip(n5820), .op(n5867) );
  nand2_1 U6308 ( .ip1(m1Inputs[56]), .ip2(\STAGE_1/weightReg [1]), .op(n5822)
         );
  nand2_1 U6309 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[51]), .op(n5821)
         );
  xor2_1 U6310 ( .ip1(n5822), .ip2(n5821), .op(n5858) );
  nand2_1 U6311 ( .ip1(m1Inputs[50]), .ip2(\STAGE_1/weightReg [7]), .op(n5823)
         );
  xor2_1 U6312 ( .ip1(n5858), .ip2(n5823), .op(n5866) );
  inv_1 U6313 ( .ip(n5824), .op(n5871) );
  fulladder U6314 ( .a(n5827), .b(n5826), .ci(n5825), .co(n5870), .s(n5838) );
  fulladder U6315 ( .a(n5830), .b(n5829), .ci(n5828), .co(n5831), .s(n5134) );
  nor2_1 U6316 ( .ip1(n5831), .ip2(n5832), .op(n5865) );
  or2_1 U6317 ( .ip1(n5831), .ip2(n5865), .op(n5834) );
  or2_1 U6318 ( .ip1(n5832), .ip2(n5865), .op(n5833) );
  nand2_1 U6319 ( .ip1(n5834), .ip2(n5833), .op(n5877) );
  fulladder U6320 ( .a(n5837), .b(n5836), .ci(n5835), .co(n5876), .s(n5839) );
  fulladder U6321 ( .a(n5840), .b(n5839), .ci(n5838), .co(n5874), .s(n5843) );
  fulladder U6322 ( .a(n5843), .b(n5842), .ci(n5841), .co(n5873), .s(
        \STAGE_1/M4/sum [0]) );
  nor2_1 U6323 ( .ip1(n5844), .ip2(n8029), .op(n6878) );
  nand2_1 U6324 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[56]), .op(n6877)
         );
  nand2_1 U6325 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[52]), .op(n6876)
         );
  inv_1 U6326 ( .ip(n5845), .op(n6894) );
  nor3_1 U6327 ( .ip1(n7813), .ip2(n6907), .ip3(n5846), .op(n5850) );
  nor2_1 U6328 ( .ip1(n5848), .ip2(n5847), .op(n5849) );
  nor2_1 U6329 ( .ip1(n5850), .ip2(n5849), .op(n6884) );
  nand2_1 U6330 ( .ip1(m1Inputs[51]), .ip2(\STAGE_1/weightReg [7]), .op(n6883)
         );
  inv_1 U6331 ( .ip(n5851), .op(n6893) );
  fulladder U6332 ( .a(n5854), .b(n5853), .ci(n5852), .co(n6892), .s(n5872) );
  nand2_1 U6333 ( .ip1(m1Inputs[54]), .ip2(\STAGE_1/weightReg [4]), .op(n5856)
         );
  nand2_1 U6334 ( .ip1(n8064), .ip2(m1Inputs[53]), .op(n5855) );
  nand2_1 U6335 ( .ip1(n5856), .ip2(n5855), .op(n5857) );
  nand3_1 U6336 ( .ip1(\STAGE_1/weightReg [5]), .ip2(m1Inputs[54]), .ip3(n5862), .op(n6871) );
  nand2_1 U6337 ( .ip1(n5857), .ip2(n6871), .op(n6873) );
  nand2_1 U6338 ( .ip1(n8009), .ip2(column[50]), .op(n6872) );
  xor2_1 U6339 ( .ip1(n6873), .ip2(n6872), .op(n6890) );
  nand3_1 U6340 ( .ip1(m1Inputs[50]), .ip2(n5858), .ip3(\STAGE_1/weightReg [7]), .op(n5860) );
  nand4_1 U6341 ( .ip1(m1Inputs[51]), .ip2(\STAGE_1/weightReg [1]), .ip3(n8037), .ip4(m1Inputs[56]), .op(n5859) );
  nand2_1 U6342 ( .ip1(n5860), .ip2(n5859), .op(n6889) );
  fulladder U6343 ( .a(n5863), .b(n5862), .ci(n5861), .co(n6888), .s(n5820) );
  inv_1 U6344 ( .ip(n5864), .op(n6898) );
  inv_1 U6345 ( .ip(n5865), .op(n6897) );
  fulladder U6346 ( .a(n5868), .b(n5867), .ci(n5866), .co(n6896), .s(n5824) );
  inv_1 U6347 ( .ip(n5869), .op(n6901) );
  fulladder U6348 ( .a(n5872), .b(n5871), .ci(n5870), .co(n6900), .s(n5878) );
  fulladder U6349 ( .a(n5875), .b(n5874), .ci(n5873), .co(n6904), .s(
        \STAGE_1/M4/sum [1]) );
  fulladder U6350 ( .a(n5878), .b(n5877), .ci(n5876), .co(n6903), .s(n5875) );
  nand2_1 U6351 ( .ip1(m1Inputs[71]), .ip2(n6280), .op(n5881) );
  nor2_1 U6352 ( .ip1(n7813), .ip2(n5879), .op(n5880) );
  xor2_1 U6353 ( .ip1(n5881), .ip2(n5880), .op(n5935) );
  nand2_1 U6354 ( .ip1(n8009), .ip2(column[65]), .op(n5934) );
  xor2_1 U6355 ( .ip1(n5935), .ip2(n5934), .op(n5941) );
  fulladder U6356 ( .a(n5884), .b(n5883), .ci(n5882), .co(n5940), .s(n5897) );
  fulladder U6357 ( .a(n5886), .b(n5903), .ci(n5885), .co(n5939), .s(n5896) );
  nor2_1 U6358 ( .ip1(n5060), .ip2(n7122), .op(n5923) );
  and3_1 U6359 ( .ip1(n8001), .ip2(m1Inputs[68]), .ip3(n5923), .op(n5890) );
  nor2_1 U6360 ( .ip1(n5888), .ip2(n5887), .op(n5889) );
  nor2_1 U6361 ( .ip1(n5890), .ip2(n5889), .op(n5929) );
  nor2_1 U6362 ( .ip1(n6246), .ip2(n7101), .op(n5924) );
  nand2_1 U6363 ( .ip1(m1Inputs[65]), .ip2(\STAGE_1/weightReg [15]), .op(n5922) );
  inv_1 U6364 ( .ip(n5891), .op(n5928) );
  nand2_1 U6365 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[67]), .op(n5893)
         );
  nand2_1 U6366 ( .ip1(m1Inputs[72]), .ip2(n6248), .op(n5892) );
  xor2_1 U6367 ( .ip1(n5893), .ip2(n5892), .op(n5918) );
  nand2_1 U6368 ( .ip1(m1Inputs[66]), .ip2(\STAGE_1/weightReg [7]), .op(n5894)
         );
  xor2_1 U6369 ( .ip1(n5918), .ip2(n5894), .op(n5927) );
  inv_1 U6370 ( .ip(n5895), .op(n5943) );
  fulladder U6371 ( .a(n5898), .b(n5897), .ci(n5896), .co(n5942), .s(n5909) );
  fulladder U6372 ( .a(n5901), .b(n5900), .ci(n5899), .co(n5902), .s(n5020) );
  nor2_1 U6373 ( .ip1(n5902), .ip2(n5903), .op(n5926) );
  or2_1 U6374 ( .ip1(n5902), .ip2(n5926), .op(n5905) );
  or2_1 U6375 ( .ip1(n5903), .ip2(n5926), .op(n5904) );
  nand2_1 U6376 ( .ip1(n5905), .ip2(n5904), .op(n5949) );
  fulladder U6377 ( .a(n5908), .b(n5907), .ci(n5906), .co(n5948), .s(n5910) );
  fulladder U6378 ( .a(n5911), .b(n5910), .ci(n5909), .co(n5946), .s(n5914) );
  fulladder U6379 ( .a(n5914), .b(n5913), .ci(n5912), .co(n5945), .s(
        \STAGE_1/M5/sum [0]) );
  nand2_1 U6380 ( .ip1(m1Inputs[70]), .ip2(n8078), .op(n5916) );
  nand2_1 U6381 ( .ip1(n8064), .ip2(m1Inputs[69]), .op(n5915) );
  nand2_1 U6382 ( .ip1(n5916), .ip2(n5915), .op(n5917) );
  nand3_1 U6383 ( .ip1(\STAGE_1/weightReg [5]), .ip2(m1Inputs[70]), .ip3(n5923), .op(n7055) );
  nand2_1 U6384 ( .ip1(n5917), .ip2(n7055), .op(n7057) );
  nand2_1 U6385 ( .ip1(n8009), .ip2(column[66]), .op(n7056) );
  xor2_1 U6386 ( .ip1(n7057), .ip2(n7056), .op(n7074) );
  nand3_1 U6387 ( .ip1(m1Inputs[66]), .ip2(n5918), .ip3(\STAGE_1/weightReg [7]), .op(n5921) );
  nand2_1 U6388 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[72]), .op(n7094)
         );
  or2_1 U6389 ( .ip1(n7094), .ip2(n5919), .op(n5920) );
  nand2_1 U6390 ( .ip1(n5921), .ip2(n5920), .op(n7073) );
  fulladder U6391 ( .a(n5924), .b(n5923), .ci(n5922), .co(n7072), .s(n5891) );
  inv_1 U6392 ( .ip(n5925), .op(n7082) );
  inv_1 U6393 ( .ip(n5926), .op(n7081) );
  fulladder U6394 ( .a(n5929), .b(n5928), .ci(n5927), .co(n7080), .s(n5895) );
  inv_1 U6395 ( .ip(n5930), .op(n7086) );
  nor2_1 U6396 ( .ip1(n5931), .ip2(n8029), .op(n7062) );
  nand2_1 U6397 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[72]), .op(n7061)
         );
  nand2_1 U6398 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[68]), .op(n7060)
         );
  inv_1 U6399 ( .ip(n5932), .op(n7078) );
  nand2_1 U6400 ( .ip1(n8064), .ip2(m1Inputs[71]), .op(n7116) );
  nor2_1 U6401 ( .ip1(n7116), .ip2(n5933), .op(n5937) );
  nor2_1 U6402 ( .ip1(n5935), .ip2(n5934), .op(n5936) );
  nor2_1 U6403 ( .ip1(n5937), .ip2(n5936), .op(n7068) );
  nand2_1 U6404 ( .ip1(m1Inputs[67]), .ip2(\STAGE_1/weightReg [7]), .op(n7067)
         );
  inv_1 U6405 ( .ip(n5938), .op(n7077) );
  fulladder U6406 ( .a(n5941), .b(n5940), .ci(n5939), .co(n7076), .s(n5944) );
  fulladder U6407 ( .a(n5944), .b(n5943), .ci(n5942), .co(n7084), .s(n5950) );
  fulladder U6408 ( .a(n5947), .b(n5946), .ci(n5945), .co(n7088), .s(
        \STAGE_1/M5/sum [1]) );
  fulladder U6409 ( .a(n5950), .b(n5949), .ci(n5948), .co(n7087), .s(n5947) );
  nand2_1 U6410 ( .ip1(m1Inputs[84]), .ip2(\STAGE_1/weightReg [5]), .op(n5952)
         );
  nand2_1 U6411 ( .ip1(m1Inputs[87]), .ip2(n6280), .op(n5951) );
  xor2_1 U6412 ( .ip1(n5952), .ip2(n5951), .op(n5991) );
  nand2_1 U6413 ( .ip1(n8009), .ip2(column[81]), .op(n5992) );
  xor2_1 U6414 ( .ip1(n5991), .ip2(n5992), .op(n5999) );
  fulladder U6415 ( .a(n5954), .b(n5953), .ci(n5977), .co(n5955), .s(n5970) );
  inv_1 U6416 ( .ip(n5955), .op(n5998) );
  fulladder U6417 ( .a(n5958), .b(n5957), .ci(n5956), .co(n5997), .s(n4913) );
  inv_1 U6418 ( .ip(n5959), .op(n6017) );
  nor2_1 U6419 ( .ip1(n6246), .ip2(n7293), .op(n6012) );
  nand2_1 U6420 ( .ip1(m1Inputs[81]), .ip2(\STAGE_1/weightReg [15]), .op(n6010) );
  inv_1 U6421 ( .ip(n5960), .op(n6003) );
  or2_1 U6422 ( .ip1(n5961), .ip2(n5962), .op(n5965) );
  or2_1 U6423 ( .ip1(n5963), .ip2(n5962), .op(n5964) );
  nand2_1 U6424 ( .ip1(n5965), .ip2(n5964), .op(n6002) );
  nand2_1 U6425 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[83]), .op(n5967)
         );
  nand2_1 U6426 ( .ip1(m1Inputs[88]), .ip2(n6248), .op(n5966) );
  xor2_1 U6427 ( .ip1(n5967), .ip2(n5966), .op(n6007) );
  nand2_1 U6428 ( .ip1(m1Inputs[82]), .ip2(\STAGE_1/weightReg [7]), .op(n5968)
         );
  xor2_1 U6429 ( .ip1(n6007), .ip2(n5968), .op(n6001) );
  inv_1 U6430 ( .ip(n5969), .op(n6016) );
  fulladder U6431 ( .a(n5972), .b(n5971), .ci(n5970), .co(n6015), .s(n5983) );
  fulladder U6432 ( .a(n5975), .b(n5974), .ci(n5973), .co(n5976), .s(n4898) );
  nor2_1 U6433 ( .ip1(n5976), .ip2(n5977), .op(n6004) );
  or2_1 U6434 ( .ip1(n5976), .ip2(n6004), .op(n5979) );
  or2_1 U6435 ( .ip1(n5977), .ip2(n6004), .op(n5978) );
  nand2_1 U6436 ( .ip1(n5979), .ip2(n5978), .op(n6022) );
  fulladder U6437 ( .a(n5982), .b(n5981), .ci(n5980), .co(n6021), .s(n5984) );
  fulladder U6438 ( .a(n5985), .b(n5984), .ci(n5983), .co(n6019), .s(n5988) );
  fulladder U6439 ( .a(n5988), .b(n5987), .ci(n5986), .co(n6018), .s(
        \STAGE_1/M6/sum [0]) );
  nor2_1 U6440 ( .ip1(n5989), .ip2(n7628), .op(n7251) );
  nand2_1 U6441 ( .ip1(n6280), .ip2(m1Inputs[88]), .op(n7250) );
  nand2_1 U6442 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[84]), .op(n7249)
         );
  nor3_1 U6443 ( .ip1(n7813), .ip2(n7279), .ip3(n5990), .op(n5993) );
  or2_1 U6444 ( .ip1(n5991), .ip2(n5993), .op(n5996) );
  inv_1 U6445 ( .ip(n5992), .op(n5994) );
  or2_1 U6446 ( .ip1(n5994), .ip2(n5993), .op(n5995) );
  nand2_1 U6447 ( .ip1(n5996), .ip2(n5995), .op(n7255) );
  nand2_1 U6448 ( .ip1(m1Inputs[83]), .ip2(\STAGE_1/weightReg [7]), .op(n7254)
         );
  fulladder U6449 ( .a(n5999), .b(n5998), .ci(n5997), .co(n7269), .s(n5959) );
  inv_1 U6450 ( .ip(n6000), .op(n7275) );
  fulladder U6451 ( .a(n6003), .b(n6002), .ci(n6001), .co(n7268), .s(n5969) );
  inv_1 U6452 ( .ip(n6004), .op(n7267) );
  nand2_1 U6453 ( .ip1(m1Inputs[86]), .ip2(n8078), .op(n6005) );
  nand2_1 U6454 ( .ip1(n8064), .ip2(m1Inputs[85]), .op(n7257) );
  nand2_1 U6455 ( .ip1(n6005), .ip2(n7257), .op(n6006) );
  nand3_1 U6456 ( .ip1(\STAGE_1/weightReg [5]), .ip2(m1Inputs[86]), .ip3(n6011), .op(n7244) );
  nand2_1 U6457 ( .ip1(n6006), .ip2(n7244), .op(n7246) );
  nand2_1 U6458 ( .ip1(n8009), .ip2(column[82]), .op(n7245) );
  xor2_1 U6459 ( .ip1(n7246), .ip2(n7245), .op(n7264) );
  nand3_1 U6460 ( .ip1(m1Inputs[82]), .ip2(n6007), .ip3(\STAGE_1/weightReg [7]), .op(n6009) );
  nand4_1 U6461 ( .ip1(n6248), .ip2(m1Inputs[83]), .ip3(\STAGE_1/weightReg [6]), .ip4(m1Inputs[88]), .op(n6008) );
  nand2_1 U6462 ( .ip1(n6009), .ip2(n6008), .op(n7263) );
  fulladder U6463 ( .a(n6012), .b(n6011), .ci(n6010), .co(n7262), .s(n5960) );
  inv_1 U6464 ( .ip(n6013), .op(n7266) );
  inv_1 U6465 ( .ip(n6014), .op(n7274) );
  fulladder U6466 ( .a(n6017), .b(n6016), .ci(n6015), .co(n7273), .s(n6023) );
  fulladder U6467 ( .a(n6020), .b(n6019), .ci(n6018), .co(n7277), .s(
        \STAGE_1/M6/sum [1]) );
  fulladder U6468 ( .a(n6023), .b(n6022), .ci(n6021), .co(n7276), .s(n6020) );
  nand2_1 U6469 ( .ip1(m1Inputs[103]), .ip2(\STAGE_1/weightReg [2]), .op(n6026) );
  nor2_1 U6470 ( .ip1(n7813), .ip2(n6024), .op(n6025) );
  xor2_1 U6471 ( .ip1(n6026), .ip2(n6025), .op(n6066) );
  nand2_1 U6472 ( .ip1(n8009), .ip2(column[97]), .op(n6065) );
  xor2_1 U6473 ( .ip1(n6066), .ip2(n6065), .op(n6072) );
  fulladder U6474 ( .a(n6029), .b(n6028), .ci(n6027), .co(n6071), .s(n6044) );
  fulladder U6475 ( .a(n6031), .b(n6050), .ci(n6030), .co(n6070), .s(n6043) );
  nor2_1 U6476 ( .ip1(n5060), .ip2(n7496), .op(n6080) );
  and2_1 U6477 ( .ip1(n6080), .ip2(n6032), .op(n6034) );
  or2_1 U6478 ( .ip1(n6033), .ip2(n6034), .op(n6037) );
  or2_1 U6479 ( .ip1(n6035), .ip2(n6034), .op(n6036) );
  nand2_1 U6480 ( .ip1(n6037), .ip2(n6036), .op(n6086) );
  nor2_1 U6481 ( .ip1(n6246), .ip2(n7475), .op(n6081) );
  nand2_1 U6482 ( .ip1(m1Inputs[97]), .ip2(\STAGE_1/weightReg [15]), .op(n6079) );
  inv_1 U6483 ( .ip(n6038), .op(n6085) );
  nand2_1 U6484 ( .ip1(n8037), .ip2(m1Inputs[99]), .op(n6040) );
  nand2_1 U6485 ( .ip1(m1Inputs[104]), .ip2(n6248), .op(n6039) );
  xor2_1 U6486 ( .ip1(n6040), .ip2(n6039), .op(n6076) );
  nand2_1 U6487 ( .ip1(m1Inputs[98]), .ip2(\STAGE_1/weightReg [7]), .op(n6041)
         );
  xor2_1 U6488 ( .ip1(n6076), .ip2(n6041), .op(n6084) );
  inv_1 U6489 ( .ip(n6042), .op(n6089) );
  fulladder U6490 ( .a(n6045), .b(n6044), .ci(n6043), .co(n6088), .s(n6056) );
  fulladder U6491 ( .a(n6048), .b(n6047), .ci(n6046), .co(n6049), .s(n4779) );
  nor2_1 U6492 ( .ip1(n6049), .ip2(n6050), .op(n6083) );
  or2_1 U6493 ( .ip1(n6049), .ip2(n6083), .op(n6052) );
  or2_1 U6494 ( .ip1(n6050), .ip2(n6083), .op(n6051) );
  nand2_1 U6495 ( .ip1(n6052), .ip2(n6051), .op(n6095) );
  fulladder U6496 ( .a(n6055), .b(n6054), .ci(n6053), .co(n6094), .s(n6057) );
  fulladder U6497 ( .a(n6058), .b(n6057), .ci(n6056), .co(n6092), .s(n6061) );
  fulladder U6498 ( .a(n6061), .b(n6060), .ci(n6059), .co(n6091), .s(
        \STAGE_1/M7/sum [0]) );
  nor2_1 U6499 ( .ip1(n6062), .ip2(n7628), .op(n7436) );
  nand2_1 U6500 ( .ip1(n6280), .ip2(m1Inputs[104]), .op(n7435) );
  nand2_1 U6501 ( .ip1(n8037), .ip2(m1Inputs[100]), .op(n7434) );
  inv_1 U6502 ( .ip(n6063), .op(n7452) );
  nand2_1 U6503 ( .ip1(n8064), .ip2(m1Inputs[103]), .op(n7490) );
  nor2_1 U6504 ( .ip1(n7490), .ip2(n6064), .op(n6068) );
  nor2_1 U6505 ( .ip1(n6066), .ip2(n6065), .op(n6067) );
  nor2_1 U6506 ( .ip1(n6068), .ip2(n6067), .op(n7442) );
  nand2_1 U6507 ( .ip1(m1Inputs[99]), .ip2(\STAGE_1/weightReg [7]), .op(n7441)
         );
  inv_1 U6508 ( .ip(n6069), .op(n7451) );
  fulladder U6509 ( .a(n6072), .b(n6071), .ci(n6070), .co(n7450), .s(n6090) );
  nand2_1 U6510 ( .ip1(m1Inputs[102]), .ip2(n8078), .op(n6074) );
  nand2_1 U6511 ( .ip1(n8064), .ip2(m1Inputs[101]), .op(n6073) );
  nand2_1 U6512 ( .ip1(n6074), .ip2(n6073), .op(n6075) );
  nand3_1 U6513 ( .ip1(\STAGE_1/weightReg [5]), .ip2(m1Inputs[102]), .ip3(
        n6080), .op(n7429) );
  nand2_1 U6514 ( .ip1(n6075), .ip2(n7429), .op(n7431) );
  nand2_1 U6515 ( .ip1(n8009), .ip2(column[98]), .op(n7430) );
  xor2_1 U6516 ( .ip1(n7431), .ip2(n7430), .op(n7448) );
  nand3_1 U6517 ( .ip1(m1Inputs[98]), .ip2(n6076), .ip3(n7882), .op(n6078) );
  nand4_1 U6518 ( .ip1(n6248), .ip2(m1Inputs[99]), .ip3(n8037), .ip4(
        m1Inputs[104]), .op(n6077) );
  nand2_1 U6519 ( .ip1(n6078), .ip2(n6077), .op(n7447) );
  fulladder U6520 ( .a(n6081), .b(n6080), .ci(n6079), .co(n7446), .s(n6038) );
  inv_1 U6521 ( .ip(n6082), .op(n7456) );
  inv_1 U6522 ( .ip(n6083), .op(n7455) );
  fulladder U6523 ( .a(n6086), .b(n6085), .ci(n6084), .co(n7454), .s(n6042) );
  inv_1 U6524 ( .ip(n6087), .op(n7459) );
  fulladder U6525 ( .a(n6090), .b(n6089), .ci(n6088), .co(n7458), .s(n6096) );
  fulladder U6526 ( .a(n6093), .b(n6092), .ci(n6091), .co(n7462), .s(
        \STAGE_1/M7/sum [1]) );
  fulladder U6527 ( .a(n6096), .b(n6095), .ci(n6094), .co(n7461), .s(n6093) );
  or2_1 U6528 ( .ip1(n6097), .ip2(n6098), .op(n6101) );
  or2_1 U6529 ( .ip1(n6099), .ip2(n6098), .op(n6100) );
  nand2_1 U6530 ( .ip1(n6101), .ip2(n6100), .op(n6148) );
  nor2_1 U6531 ( .ip1(n6246), .ip2(n7663), .op(n6143) );
  nand2_1 U6532 ( .ip1(m1Inputs[113]), .ip2(\STAGE_1/weightReg [15]), .op(
        n6141) );
  inv_1 U6533 ( .ip(n6102), .op(n6147) );
  nand2_1 U6534 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[115]), .op(n6104) );
  nand2_1 U6535 ( .ip1(m1Inputs[120]), .ip2(n6248), .op(n6103) );
  xor2_1 U6536 ( .ip1(n6104), .ip2(n6103), .op(n6138) );
  nand2_1 U6537 ( .ip1(m1Inputs[114]), .ip2(\STAGE_1/weightReg [7]), .op(n6105) );
  xor2_1 U6538 ( .ip1(n6138), .ip2(n6105), .op(n6146) );
  inv_1 U6539 ( .ip(n6106), .op(n6163) );
  nand2_1 U6540 ( .ip1(m1Inputs[119]), .ip2(\STAGE_1/weightReg [2]), .op(n6109) );
  nor2_1 U6541 ( .ip1(n7813), .ip2(n6107), .op(n6108) );
  xor2_1 U6542 ( .ip1(n6109), .ip2(n6108), .op(n6154) );
  nand2_1 U6543 ( .ip1(n8175), .ip2(column[113]), .op(n6153) );
  xor2_1 U6544 ( .ip1(n6154), .ip2(n6153), .op(n6160) );
  fulladder U6545 ( .a(n6112), .b(n6111), .ci(n6110), .co(n6159), .s(n6117) );
  fulladder U6546 ( .a(n6114), .b(n6122), .ci(n6113), .co(n6158), .s(n6115) );
  fulladder U6547 ( .a(n6117), .b(n6116), .ci(n6115), .co(n6161), .s(n6128) );
  fulladder U6548 ( .a(n6120), .b(n6119), .ci(n6118), .co(n6121), .s(n4660) );
  nor2_1 U6549 ( .ip1(n6121), .ip2(n6122), .op(n6145) );
  or2_1 U6550 ( .ip1(n6121), .ip2(n6145), .op(n6124) );
  or2_1 U6551 ( .ip1(n6122), .ip2(n6145), .op(n6123) );
  nand2_1 U6552 ( .ip1(n6124), .ip2(n6123), .op(n6168) );
  fulladder U6553 ( .a(n6127), .b(n6126), .ci(n6125), .co(n6167), .s(n6129) );
  fulladder U6554 ( .a(n6130), .b(n6129), .ci(n6128), .co(n6165), .s(n6133) );
  fulladder U6555 ( .a(n6133), .b(n6132), .ci(n6131), .co(n6164), .s(
        \STAGE_1/M8/sum [0]) );
  nand2_1 U6556 ( .ip1(\STAGE_1/weightReg [5]), .ip2(m1Inputs[118]), .op(n7675) );
  nor3_1 U6557 ( .ip1(n5060), .ip2(n7675), .ip3(n7684), .op(n7619) );
  nor2_1 U6558 ( .ip1(n7813), .ip2(n7684), .op(n6134) );
  or2_1 U6559 ( .ip1(m1Inputs[118]), .ip2(n6134), .op(n6136) );
  or2_1 U6560 ( .ip1(n8078), .ip2(n6134), .op(n6135) );
  nand2_1 U6561 ( .ip1(n6136), .ip2(n6135), .op(n7617) );
  or2_1 U6562 ( .ip1(n7619), .ip2(n7617), .op(n6137) );
  nand2_1 U6563 ( .ip1(n8175), .ip2(column[114]), .op(n7616) );
  xor2_1 U6564 ( .ip1(n6137), .ip2(n7616), .op(n7636) );
  nand3_1 U6565 ( .ip1(m1Inputs[114]), .ip2(n6138), .ip3(
        \STAGE_1/weightReg [7]), .op(n6140) );
  nand4_1 U6566 ( .ip1(n6248), .ip2(m1Inputs[115]), .ip3(
        \STAGE_1/weightReg [6]), .ip4(m1Inputs[120]), .op(n6139) );
  nand2_1 U6567 ( .ip1(n6140), .ip2(n6139), .op(n7635) );
  fulladder U6568 ( .a(n6143), .b(n6142), .ci(n6141), .co(n7634), .s(n6102) );
  inv_1 U6569 ( .ip(n6144), .op(n7644) );
  inv_1 U6570 ( .ip(n6145), .op(n7643) );
  fulladder U6571 ( .a(n6148), .b(n6147), .ci(n6146), .co(n7642), .s(n6106) );
  inv_1 U6572 ( .ip(n6149), .op(n7648) );
  nor2_1 U6573 ( .ip1(n6150), .ip2(n7628), .op(n7622) );
  nand2_1 U6574 ( .ip1(n6280), .ip2(m1Inputs[120]), .op(n7621) );
  nand2_1 U6575 ( .ip1(n8037), .ip2(m1Inputs[116]), .op(n7620) );
  inv_1 U6576 ( .ip(n6151), .op(n7640) );
  nand2_1 U6577 ( .ip1(n8064), .ip2(m1Inputs[119]), .op(n7678) );
  nor2_1 U6578 ( .ip1(n7678), .ip2(n6152), .op(n6156) );
  nor2_1 U6579 ( .ip1(n6154), .ip2(n6153), .op(n6155) );
  nor2_1 U6580 ( .ip1(n6156), .ip2(n6155), .op(n7632) );
  nand2_1 U6581 ( .ip1(m1Inputs[115]), .ip2(\STAGE_1/weightReg [7]), .op(n7630) );
  inv_1 U6582 ( .ip(n6157), .op(n7639) );
  fulladder U6583 ( .a(n6160), .b(n6159), .ci(n6158), .co(n7638), .s(n6162) );
  fulladder U6584 ( .a(n6163), .b(n6162), .ci(n6161), .co(n7646), .s(n6169) );
  fulladder U6585 ( .a(n6166), .b(n6165), .ci(n6164), .co(n7650), .s(
        \STAGE_1/M8/sum [1]) );
  fulladder U6586 ( .a(n6169), .b(n6168), .ci(n6167), .co(n7649), .s(n6166) );
  nor2_1 U6587 ( .ip1(n5060), .ip2(n7865), .op(n6213) );
  and3_1 U6588 ( .ip1(n8001), .ip2(m1Inputs[132]), .ip3(n6213), .op(n6171) );
  or2_1 U6589 ( .ip1(n6170), .ip2(n6171), .op(n6174) );
  or2_1 U6590 ( .ip1(n6172), .ip2(n6171), .op(n6173) );
  nand2_1 U6591 ( .ip1(n6174), .ip2(n6173), .op(n6219) );
  nor2_1 U6592 ( .ip1(n6246), .ip2(n7849), .op(n6214) );
  nand2_1 U6593 ( .ip1(m1Inputs[129]), .ip2(\STAGE_1/weightReg [15]), .op(
        n6212) );
  inv_1 U6594 ( .ip(n6175), .op(n6218) );
  nand2_1 U6595 ( .ip1(n8037), .ip2(m1Inputs[131]), .op(n6177) );
  nand2_1 U6596 ( .ip1(m1Inputs[136]), .ip2(n6248), .op(n6176) );
  xor2_1 U6597 ( .ip1(n6177), .ip2(n6176), .op(n6209) );
  nand2_1 U6598 ( .ip1(m1Inputs[130]), .ip2(n7882), .op(n6178) );
  xor2_1 U6599 ( .ip1(n6209), .ip2(n6178), .op(n6217) );
  inv_1 U6600 ( .ip(n6179), .op(n6234) );
  nand2_1 U6601 ( .ip1(m1Inputs[135]), .ip2(\STAGE_1/weightReg [2]), .op(n6181) );
  nor2_1 U6602 ( .ip1(n7813), .ip2(n7881), .op(n6180) );
  xor2_1 U6603 ( .ip1(n6181), .ip2(n6180), .op(n6225) );
  nand2_1 U6604 ( .ip1(n8175), .ip2(column[129]), .op(n6224) );
  xor2_1 U6605 ( .ip1(n6225), .ip2(n6224), .op(n6231) );
  fulladder U6606 ( .a(n6184), .b(n6183), .ci(n6182), .co(n6230), .s(n6188) );
  fulladder U6607 ( .a(n6186), .b(n6194), .ci(n6185), .co(n6229), .s(n6187) );
  fulladder U6608 ( .a(n6189), .b(n6188), .ci(n6187), .co(n6232), .s(n6200) );
  fulladder U6609 ( .a(n6192), .b(n6191), .ci(n6190), .co(n6193), .s(n4542) );
  nor2_1 U6610 ( .ip1(n6193), .ip2(n6194), .op(n6216) );
  or2_1 U6611 ( .ip1(n6193), .ip2(n6216), .op(n6196) );
  or2_1 U6612 ( .ip1(n6194), .ip2(n6216), .op(n6195) );
  nand2_1 U6613 ( .ip1(n6196), .ip2(n6195), .op(n6239) );
  fulladder U6614 ( .a(n6199), .b(n6198), .ci(n6197), .co(n6238), .s(n6201) );
  fulladder U6615 ( .a(n6202), .b(n6201), .ci(n6200), .co(n6236), .s(n6205) );
  fulladder U6616 ( .a(n6205), .b(n6204), .ci(n6203), .co(n6235), .s(
        \STAGE_1/M9/sum [0]) );
  nand2_1 U6617 ( .ip1(m1Inputs[134]), .ip2(n8078), .op(n6207) );
  nand2_1 U6618 ( .ip1(\STAGE_1/weightReg [5]), .ip2(m1Inputs[133]), .op(n6206) );
  nand2_1 U6619 ( .ip1(n6207), .ip2(n6206), .op(n6208) );
  nand3_1 U6620 ( .ip1(\STAGE_1/weightReg [5]), .ip2(m1Inputs[134]), .ip3(
        n6213), .op(n7804) );
  nand2_1 U6621 ( .ip1(n6208), .ip2(n7804), .op(n7806) );
  nand2_1 U6622 ( .ip1(n8175), .ip2(column[130]), .op(n7805) );
  xor2_1 U6623 ( .ip1(n7806), .ip2(n7805), .op(n7824) );
  nand3_1 U6624 ( .ip1(m1Inputs[130]), .ip2(n6209), .ip3(
        \STAGE_1/weightReg [7]), .op(n6211) );
  nand4_1 U6625 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[131]), .ip3(
        \STAGE_1/weightReg [6]), .ip4(m1Inputs[136]), .op(n6210) );
  nand2_1 U6626 ( .ip1(n6211), .ip2(n6210), .op(n7823) );
  fulladder U6627 ( .a(n6214), .b(n6213), .ci(n6212), .co(n7822), .s(n6175) );
  inv_1 U6628 ( .ip(n6215), .op(n7832) );
  inv_1 U6629 ( .ip(n6216), .op(n7831) );
  fulladder U6630 ( .a(n6219), .b(n6218), .ci(n6217), .co(n7830), .s(n6179) );
  inv_1 U6631 ( .ip(n6220), .op(n7836) );
  inv_1 U6632 ( .ip(\STAGE_1/weightReg [15]), .op(n8029) );
  nor2_1 U6633 ( .ip1(n6221), .ip2(n8029), .op(n7811) );
  nand2_1 U6634 ( .ip1(n6280), .ip2(m1Inputs[136]), .op(n7810) );
  nand2_1 U6635 ( .ip1(n8037), .ip2(m1Inputs[132]), .op(n7809) );
  inv_1 U6636 ( .ip(n6222), .op(n7828) );
  nor3_1 U6637 ( .ip1(n7813), .ip2(n7841), .ip3(n6223), .op(n6227) );
  nor2_1 U6638 ( .ip1(n6225), .ip2(n6224), .op(n6226) );
  nor2_1 U6639 ( .ip1(n6227), .ip2(n6226), .op(n7818) );
  nand2_1 U6640 ( .ip1(m1Inputs[131]), .ip2(\STAGE_1/weightReg [7]), .op(n7817) );
  inv_1 U6641 ( .ip(n6228), .op(n7827) );
  fulladder U6642 ( .a(n6231), .b(n6230), .ci(n6229), .co(n7826), .s(n6233) );
  fulladder U6643 ( .a(n6234), .b(n6233), .ci(n6232), .co(n7834), .s(n6240) );
  fulladder U6644 ( .a(n6237), .b(n6236), .ci(n6235), .co(n7838), .s(
        \STAGE_1/M9/sum [1]) );
  fulladder U6645 ( .a(n6240), .b(n6239), .ci(n6238), .co(n7837), .s(n6237) );
  or2_1 U6646 ( .ip1(n6241), .ip2(n6242), .op(n6245) );
  or2_1 U6647 ( .ip1(n6243), .ip2(n6242), .op(n6244) );
  nand2_1 U6648 ( .ip1(n6245), .ip2(n6244), .op(n6304) );
  nor2_1 U6649 ( .ip1(n6246), .ip2(n8046), .op(n6299) );
  nand2_1 U6650 ( .ip1(m1Inputs[145]), .ip2(\STAGE_1/weightReg [15]), .op(
        n6297) );
  inv_1 U6651 ( .ip(n6247), .op(n6303) );
  nand2_1 U6652 ( .ip1(n8037), .ip2(m1Inputs[147]), .op(n6250) );
  nand2_1 U6653 ( .ip1(m1Inputs[152]), .ip2(n6248), .op(n6249) );
  xor2_1 U6654 ( .ip1(n6250), .ip2(n6249), .op(n6293) );
  nand2_1 U6655 ( .ip1(m1Inputs[146]), .ip2(\STAGE_1/weightReg [7]), .op(n6251) );
  xor2_1 U6656 ( .ip1(n6293), .ip2(n6251), .op(n6302) );
  inv_1 U6657 ( .ip(n6252), .op(n6308) );
  nand2_1 U6658 ( .ip1(m1Inputs[151]), .ip2(\STAGE_1/weightReg [2]), .op(n6254) );
  nor2_1 U6659 ( .ip1(n7813), .ip2(n8077), .op(n6253) );
  xor2_1 U6660 ( .ip1(n6254), .ip2(n6253), .op(n6284) );
  nand2_1 U6661 ( .ip1(n8175), .ip2(column[145]), .op(n6283) );
  xor2_1 U6662 ( .ip1(n6284), .ip2(n6283), .op(n6290) );
  fulladder U6663 ( .a(n6257), .b(n6256), .ci(n6255), .co(n6289), .s(n6261) );
  fulladder U6664 ( .a(n6259), .b(n6267), .ci(n6258), .co(n6288), .s(n6260) );
  fulladder U6665 ( .a(n6262), .b(n6261), .ci(n6260), .co(n6306), .s(n6273) );
  fulladder U6666 ( .a(n6265), .b(n6264), .ci(n6263), .co(n6266), .s(n4423) );
  nor2_1 U6667 ( .ip1(n6266), .ip2(n6267), .op(n6301) );
  or2_1 U6668 ( .ip1(n6266), .ip2(n6301), .op(n6269) );
  or2_1 U6669 ( .ip1(n6267), .ip2(n6301), .op(n6268) );
  nand2_1 U6670 ( .ip1(n6269), .ip2(n6268), .op(n6313) );
  fulladder U6671 ( .a(n6272), .b(n6271), .ci(n6270), .co(n6312), .s(n6274) );
  fulladder U6672 ( .a(n6275), .b(n6274), .ci(n6273), .co(n6310), .s(n6278) );
  fulladder U6673 ( .a(n6278), .b(n6277), .ci(n6276), .co(n6309), .s(
        \STAGE_1/M10/sum [0]) );
  nor2_1 U6674 ( .ip1(n6279), .ip2(n8029), .op(n7998) );
  nand2_1 U6675 ( .ip1(n6280), .ip2(m1Inputs[152]), .op(n7997) );
  nand2_1 U6676 ( .ip1(n8037), .ip2(m1Inputs[148]), .op(n7996) );
  inv_1 U6677 ( .ip(n6281), .op(n8017) );
  nor3_1 U6678 ( .ip1(n7813), .ip2(n8031), .ip3(n6282), .op(n6286) );
  nor2_1 U6679 ( .ip1(n6284), .ip2(n6283), .op(n6285) );
  nor2_1 U6680 ( .ip1(n6286), .ip2(n6285), .op(n8003) );
  nand2_1 U6681 ( .ip1(m1Inputs[147]), .ip2(\STAGE_1/weightReg [7]), .op(n8002) );
  inv_1 U6682 ( .ip(n6287), .op(n8016) );
  fulladder U6683 ( .a(n6290), .b(n6289), .ci(n6288), .co(n8015), .s(n6307) );
  nand2_1 U6684 ( .ip1(m1Inputs[150]), .ip2(\STAGE_1/weightReg [4]), .op(n6291) );
  nand2_1 U6685 ( .ip1(\STAGE_1/weightReg [5]), .ip2(m1Inputs[149]), .op(n8005) );
  nand2_1 U6686 ( .ip1(n6291), .ip2(n8005), .op(n6292) );
  nand3_1 U6687 ( .ip1(\STAGE_1/weightReg [5]), .ip2(m1Inputs[150]), .ip3(
        n6298), .op(n7991) );
  nand2_1 U6688 ( .ip1(n6292), .ip2(n7991), .op(n7993) );
  nand2_1 U6689 ( .ip1(n8175), .ip2(column[146]), .op(n7992) );
  xor2_1 U6690 ( .ip1(n7993), .ip2(n7992), .op(n8013) );
  nand3_1 U6691 ( .ip1(m1Inputs[146]), .ip2(n6293), .ip3(
        \STAGE_1/weightReg [7]), .op(n6296) );
  nand2_1 U6692 ( .ip1(n8037), .ip2(m1Inputs[152]), .op(n8039) );
  or2_1 U6693 ( .ip1(n8039), .ip2(n6294), .op(n6295) );
  nand2_1 U6694 ( .ip1(n6296), .ip2(n6295), .op(n8012) );
  fulladder U6695 ( .a(n6299), .b(n6298), .ci(n6297), .co(n8011), .s(n6247) );
  inv_1 U6696 ( .ip(n6300), .op(n8021) );
  inv_1 U6697 ( .ip(n6301), .op(n8020) );
  fulladder U6698 ( .a(n6304), .b(n6303), .ci(n6302), .co(n8019), .s(n6252) );
  inv_1 U6699 ( .ip(n6305), .op(n8024) );
  fulladder U6700 ( .a(n6308), .b(n6307), .ci(n6306), .co(n8023), .s(n6314) );
  fulladder U6701 ( .a(n6311), .b(n6310), .ci(n6309), .co(n8027), .s(
        \STAGE_1/M10/sum [1]) );
  fulladder U6702 ( .a(n6314), .b(n6313), .ci(n6312), .co(n8026), .s(n6311) );
  nand2_1 U6703 ( .ip1(m1Inputs[7]), .ip2(\STAGE_1/weightReg [4]), .op(n6417)
         );
  inv_1 U6704 ( .ip(n6315), .op(n6319) );
  nor2_1 U6705 ( .ip1(n6317), .ip2(n6316), .op(n6318) );
  nor2_1 U6706 ( .ip1(n6319), .ip2(n6318), .op(n6416) );
  fulladder U6707 ( .a(n6322), .b(n6321), .ci(n6320), .co(n6415), .s(n5645) );
  inv_1 U6708 ( .ip(n6323), .op(n6431) );
  nand2_1 U6709 ( .ip1(m1Inputs[6]), .ip2(\STAGE_1/weightReg [5]), .op(n6376)
         );
  nand2_1 U6710 ( .ip1(n8037), .ip2(m1Inputs[6]), .op(n6378) );
  nor3_1 U6711 ( .ip1(n6378), .ip2(n7813), .ip3(n6375), .op(n6400) );
  or2_1 U6712 ( .ip1(n6376), .ip2(n6400), .op(n6326) );
  nand2_1 U6713 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[5]), .op(n6324)
         );
  or2_1 U6714 ( .ip1(n6324), .ip2(n6400), .op(n6325) );
  nand2_1 U6715 ( .ip1(n6326), .ip2(n6325), .op(n6398) );
  nand2_1 U6716 ( .ip1(n7045), .ip2(column[3]), .op(n6399) );
  xor2_1 U6717 ( .ip1(n6398), .ip2(n6399), .op(n6427) );
  fulladder U6718 ( .a(n6329), .b(n6328), .ci(n6327), .co(n6426), .s(n5651) );
  nand2_1 U6719 ( .ip1(\STAGE_1/weightReg [7]), .ip2(m1Inputs[4]), .op(n6406)
         );
  nor2_1 U6720 ( .ip1(n6330), .ip2(n8029), .op(n6405) );
  nand2_1 U6721 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[8]), .op(n6404)
         );
  inv_1 U6722 ( .ip(n6331), .op(n6430) );
  fulladder U6723 ( .a(n6334), .b(n6333), .ci(n6332), .co(n6429), .s(n5638) );
  inv_1 U6724 ( .ip(n6335), .op(n6443) );
  fulladder U6725 ( .a(n6338), .b(n6337), .ci(n6336), .co(n6339), .s(n6345) );
  inv_1 U6726 ( .ip(n6339), .op(n6442) );
  fulladder U6727 ( .a(n6342), .b(n6341), .ci(n6340), .co(n6441), .s(n5643) );
  inv_1 U6728 ( .ip(n6343), .op(n6439) );
  fulladder U6729 ( .a(n6346), .b(n6345), .ci(n6344), .co(n6438), .s(n6349) );
  fulladder U6730 ( .a(n6349), .b(n6348), .ci(n6347), .co(n6437), .s(
        \STAGE_1/M1/sum [2]) );
  inv_1 U6731 ( .ip(column[12]), .op(n6484) );
  nor2_1 U6732 ( .ip1(n8180), .ip2(n6484), .op(n6490) );
  nor2_1 U6733 ( .ip1(n6350), .ip2(n8029), .op(n6446) );
  nand2_1 U6734 ( .ip1(n7882), .ip2(m1Inputs[8]), .op(n6354) );
  nor2_1 U6735 ( .ip1(n6351), .ip2(n8029), .op(n6353) );
  nand2_1 U6736 ( .ip1(n7045), .ip2(column[7]), .op(n6352) );
  nand2_1 U6737 ( .ip1(n7045), .ip2(column[8]), .op(n6444) );
  fulladder U6738 ( .a(n6354), .b(n6353), .ci(n6352), .co(n6445), .s(n6371) );
  nand2_1 U6739 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[7]), .op(n6377)
         );
  nor2_1 U6740 ( .ip1(n6354), .ip2(n6377), .op(n6359) );
  buf_1 U6741 ( .ip(n8175), .op(n8051) );
  nand2_1 U6742 ( .ip1(\STAGE_1/weightReg [7]), .ip2(m1Inputs[7]), .op(n6363)
         );
  or2_1 U6743 ( .ip1(n6363), .ip2(n6359), .op(n6357) );
  nand2_1 U6744 ( .ip1(m1Inputs[8]), .ip2(n8037), .op(n6355) );
  or2_1 U6745 ( .ip1(n6355), .ip2(n6359), .op(n6356) );
  nand2_1 U6746 ( .ip1(n6357), .ip2(n6356), .op(n6361) );
  and3_1 U6747 ( .ip1(n8051), .ip2(column[6]), .ip3(n6361), .op(n6358) );
  nor2_1 U6748 ( .ip1(n6359), .ip2(n6358), .op(n6370) );
  nand2_1 U6749 ( .ip1(n7045), .ip2(column[6]), .op(n6360) );
  xor2_1 U6750 ( .ip1(n6361), .ip2(n6360), .op(n6374) );
  nor2_1 U6751 ( .ip1(n6362), .ip2(n7628), .op(n6373) );
  nor2_1 U6752 ( .ip1(n6363), .ip2(n6378), .op(n6368) );
  or2_1 U6753 ( .ip1(n6377), .ip2(n6368), .op(n6366) );
  nand2_1 U6754 ( .ip1(\STAGE_1/weightReg [7]), .ip2(m1Inputs[6]), .op(n6364)
         );
  or2_1 U6755 ( .ip1(n6364), .ip2(n6368), .op(n6365) );
  nand2_1 U6756 ( .ip1(n6366), .ip2(n6365), .op(n6387) );
  and3_1 U6757 ( .ip1(n8051), .ip2(column[5]), .ip3(n6387), .op(n6367) );
  nor2_1 U6758 ( .ip1(n6368), .ip2(n6367), .op(n6372) );
  fulladder U6759 ( .a(n6371), .b(n6370), .ci(n6369), .co(n6465), .s(n6470) );
  fulladder U6760 ( .a(n6374), .b(n6373), .ci(n6372), .co(n6369), .s(n6394) );
  nand2_1 U6761 ( .ip1(m1Inputs[8]), .ip2(\STAGE_1/weightReg [5]), .op(n6390)
         );
  nor2_1 U6762 ( .ip1(n6375), .ip2(n8029), .op(n6389) );
  nor2_1 U6763 ( .ip1(n6377), .ip2(n6376), .op(n6382) );
  or2_1 U6764 ( .ip1(n6378), .ip2(n6382), .op(n6381) );
  nand2_1 U6765 ( .ip1(m1Inputs[7]), .ip2(\STAGE_1/weightReg [5]), .op(n6379)
         );
  or2_1 U6766 ( .ip1(n6379), .ip2(n6382), .op(n6380) );
  nand2_1 U6767 ( .ip1(n6381), .ip2(n6380), .op(n6408) );
  or2_1 U6768 ( .ip1(n6408), .ip2(n6382), .op(n6385) );
  nand2_1 U6769 ( .ip1(n7045), .ip2(column[4]), .op(n6407) );
  inv_1 U6770 ( .ip(n6407), .op(n6383) );
  or2_1 U6771 ( .ip1(n6383), .ip2(n6382), .op(n6384) );
  nand2_1 U6772 ( .ip1(n6385), .ip2(n6384), .op(n6388) );
  nand2_1 U6773 ( .ip1(n7045), .ip2(column[5]), .op(n6386) );
  xor2_1 U6774 ( .ip1(n6387), .ip2(n6386), .op(n6397) );
  fulladder U6775 ( .a(n6390), .b(n6389), .ci(n6388), .co(n6393), .s(n6396) );
  nor2_1 U6776 ( .ip1(n6391), .ip2(n8029), .op(n6411) );
  nand2_1 U6777 ( .ip1(\STAGE_1/weightReg [7]), .ip2(m1Inputs[5]), .op(n6410)
         );
  nand2_1 U6778 ( .ip1(m1Inputs[8]), .ip2(\STAGE_1/weightReg [4]), .op(n6409)
         );
  fulladder U6779 ( .a(n6394), .b(n6393), .ci(n6392), .co(n6469), .s(n6474) );
  fulladder U6780 ( .a(n6397), .b(n6396), .ci(n6395), .co(n6392), .s(n6420) );
  or2_1 U6781 ( .ip1(n6398), .ip2(n6400), .op(n6403) );
  inv_1 U6782 ( .ip(n6399), .op(n6401) );
  or2_1 U6783 ( .ip1(n6401), .ip2(n6400), .op(n6402) );
  nand2_1 U6784 ( .ip1(n6403), .ip2(n6402), .op(n6414) );
  fulladder U6785 ( .a(n6406), .b(n6405), .ci(n6404), .co(n6413), .s(n6425) );
  xor2_1 U6786 ( .ip1(n6408), .ip2(n6407), .op(n6412) );
  fulladder U6787 ( .a(n6411), .b(n6410), .ci(n6409), .co(n6395), .s(n6423) );
  fulladder U6788 ( .a(n6414), .b(n6413), .ci(n6412), .co(n6419), .s(n6422) );
  fulladder U6789 ( .a(n6417), .b(n6416), .ci(n6415), .co(n6421), .s(n6323) );
  fulladder U6790 ( .a(n6420), .b(n6419), .ci(n6418), .co(n6473), .s(n6478) );
  fulladder U6791 ( .a(n6423), .b(n6422), .ci(n6421), .co(n6418), .s(n6424) );
  inv_1 U6792 ( .ip(n6424), .op(n6435) );
  fulladder U6793 ( .a(n6427), .b(n6426), .ci(n6425), .co(n6428), .s(n6331) );
  inv_1 U6794 ( .ip(n6428), .op(n6434) );
  fulladder U6795 ( .a(n6431), .b(n6430), .ci(n6429), .co(n6433), .s(n6335) );
  inv_1 U6796 ( .ip(n6432), .op(n6477) );
  fulladder U6797 ( .a(n6435), .b(n6434), .ci(n6433), .co(n6432), .s(n6436) );
  inv_1 U6798 ( .ip(n6436), .op(n6482) );
  fulladder U6799 ( .a(n6439), .b(n6438), .ci(n6437), .co(n6440), .s(
        \STAGE_1/M1/sum [3]) );
  inv_1 U6800 ( .ip(n6440), .op(n6481) );
  fulladder U6801 ( .a(n6443), .b(n6442), .ci(n6441), .co(n6480), .s(n6343) );
  fulladder U6802 ( .a(n6446), .b(n6445), .ci(n6444), .co(n6457), .s(n6466) );
  nand2_1 U6803 ( .ip1(n7045), .ip2(column[9]), .op(n6462) );
  nor3_1 U6804 ( .ip1(n6458), .ip2(n6457), .ip3(n6462), .op(n6453) );
  nand3_1 U6805 ( .ip1(column[11]), .ip2(n6453), .ip3(column[10]), .op(n6448)
         );
  and2_1 U6806 ( .ip1(n8051), .ip2(column[11]), .op(n6452) );
  nand2_1 U6807 ( .ip1(n7045), .ip2(column[10]), .op(n6456) );
  nand4_1 U6808 ( .ip1(n6458), .ip2(n6457), .ip3(n6456), .ip4(n6462), .op(
        n6449) );
  nor2_1 U6809 ( .ip1(n6452), .ip2(n6449), .op(n6487) );
  inv_1 U6810 ( .ip(n6487), .op(n6447) );
  nand2_1 U6811 ( .ip1(n6448), .ip2(n6447), .op(n6485) );
  xor2_1 U6812 ( .ip1(n6490), .ip2(n6485), .op(\STAGE_1/M1/sum [12]) );
  nand2_1 U6813 ( .ip1(column[10]), .ip2(n6453), .op(n6450) );
  nand2_1 U6814 ( .ip1(n6450), .ip2(n6449), .op(n6451) );
  xor2_1 U6815 ( .ip1(n6452), .ip2(n6451), .op(\STAGE_1/M1/sum [11]) );
  and3_1 U6816 ( .ip1(n6458), .ip2(n6457), .ip3(n6462), .op(n6454) );
  nor2_1 U6817 ( .ip1(n6454), .ip2(n6453), .op(n6455) );
  xor2_1 U6818 ( .ip1(n6456), .ip2(n6455), .op(\STAGE_1/M1/sum [10]) );
  inv_1 U6819 ( .ip(n6462), .op(n6463) );
  nand2_1 U6820 ( .ip1(n6458), .ip2(n6457), .op(n6460) );
  or2_1 U6821 ( .ip1(n6458), .ip2(n6457), .op(n6459) );
  nand2_1 U6822 ( .ip1(n6460), .ip2(n6459), .op(n6461) );
  mux2_1 U6823 ( .ip1(n6463), .ip2(n6462), .s(n6461), .op(\STAGE_1/M1/sum [9])
         );
  fulladder U6824 ( .a(n6466), .b(n6465), .ci(n6464), .co(n6458), .s(n6467) );
  inv_1 U6825 ( .ip(n6467), .op(\STAGE_1/M1/sum [8]) );
  fulladder U6826 ( .a(n6470), .b(n6469), .ci(n6468), .co(n6464), .s(n6471) );
  inv_1 U6827 ( .ip(n6471), .op(\STAGE_1/M1/sum [7]) );
  fulladder U6828 ( .a(n6474), .b(n6473), .ci(n6472), .co(n6468), .s(n6475) );
  inv_1 U6829 ( .ip(n6475), .op(\STAGE_1/M1/sum [6]) );
  fulladder U6830 ( .a(n6478), .b(n6477), .ci(n6476), .co(n6472), .s(n6479) );
  inv_1 U6831 ( .ip(n6479), .op(\STAGE_1/M1/sum [5]) );
  fulladder U6832 ( .a(n6482), .b(n6481), .ci(n6480), .co(n6476), .s(n6483) );
  inv_1 U6833 ( .ip(n6483), .op(\STAGE_1/M1/sum [4]) );
  nor3_1 U6834 ( .ip1(n8180), .ip2(n6485), .ip3(n6484), .op(n6486) );
  nor2_1 U6835 ( .ip1(n6487), .ip2(n6486), .op(n6489) );
  nand2_1 U6836 ( .ip1(n8009), .ip2(column[13]), .op(n6488) );
  inv_1 U6837 ( .ip(n6488), .op(n6494) );
  fulladder U6838 ( .a(n6490), .b(n6489), .ci(n6488), .co(n6493), .s(
        \STAGE_1/M1/sum [13]) );
  nand2_1 U6839 ( .ip1(n7045), .ip2(column[14]), .op(n6492) );
  nor2_1 U6840 ( .ip1(column[14]), .ip2(column[15]), .op(n6491) );
  not_ab_or_c_or_d U6841 ( .ip1(column[14]), .ip2(column[15]), .ip3(n6491), 
        .ip4(n8180), .op(n6496) );
  fulladder U6842 ( .a(n6494), .b(n6493), .ci(n6492), .co(n6495), .s(
        \STAGE_1/M1/sum [14]) );
  xnor2_1 U6843 ( .ip1(n6496), .ip2(n6495), .op(\STAGE_1/M1/sum [15]) );
  nand2_1 U6844 ( .ip1(n8078), .ip2(m1Inputs[23]), .op(n6599) );
  inv_1 U6845 ( .ip(n6497), .op(n6501) );
  nor2_1 U6846 ( .ip1(n6499), .ip2(n6498), .op(n6500) );
  nor2_1 U6847 ( .ip1(n6501), .ip2(n6500), .op(n6598) );
  fulladder U6848 ( .a(n6504), .b(n6503), .ci(n6502), .co(n6597), .s(n5716) );
  inv_1 U6849 ( .ip(n6505), .op(n6613) );
  nand2_1 U6850 ( .ip1(n8064), .ip2(m1Inputs[22]), .op(n6558) );
  nand2_1 U6851 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[22]), .op(n6560)
         );
  nor3_1 U6852 ( .ip1(n7813), .ip2(n6560), .ip3(n6557), .op(n6582) );
  or2_1 U6853 ( .ip1(n6558), .ip2(n6582), .op(n6508) );
  nand2_1 U6854 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[21]), .op(n6506)
         );
  or2_1 U6855 ( .ip1(n6506), .ip2(n6582), .op(n6507) );
  nand2_1 U6856 ( .ip1(n6508), .ip2(n6507), .op(n6580) );
  nand2_1 U6857 ( .ip1(n7045), .ip2(column[19]), .op(n6581) );
  xor2_1 U6858 ( .ip1(n6580), .ip2(n6581), .op(n6609) );
  fulladder U6859 ( .a(n6511), .b(n6510), .ci(n6509), .co(n6608), .s(n5722) );
  inv_1 U6860 ( .ip(n7685), .op(n7882) );
  nand2_1 U6861 ( .ip1(n7882), .ip2(m1Inputs[20]), .op(n6588) );
  nor2_1 U6862 ( .ip1(n6512), .ip2(n8029), .op(n6587) );
  nand2_1 U6863 ( .ip1(n8001), .ip2(m1Inputs[24]), .op(n6586) );
  inv_1 U6864 ( .ip(n6513), .op(n6612) );
  fulladder U6865 ( .a(n6516), .b(n6515), .ci(n6514), .co(n6611), .s(n5709) );
  inv_1 U6866 ( .ip(n6517), .op(n6625) );
  fulladder U6867 ( .a(n6520), .b(n6519), .ci(n6518), .co(n6521), .s(n6527) );
  inv_1 U6868 ( .ip(n6521), .op(n6624) );
  fulladder U6869 ( .a(n6524), .b(n6523), .ci(n6522), .co(n6623), .s(n5714) );
  inv_1 U6870 ( .ip(n6525), .op(n6621) );
  fulladder U6871 ( .a(n6528), .b(n6527), .ci(n6526), .co(n6620), .s(n6531) );
  fulladder U6872 ( .a(n6531), .b(n6530), .ci(n6529), .co(n6619), .s(
        \STAGE_1/M2/sum [2]) );
  and2_1 U6873 ( .ip1(n8051), .ip2(column[29]), .op(n6679) );
  nand2_1 U6874 ( .ip1(n7045), .ip2(column[27]), .op(n6640) );
  nor2_1 U6875 ( .ip1(n6532), .ip2(n8029), .op(n6628) );
  nand2_1 U6876 ( .ip1(n7882), .ip2(m1Inputs[24]), .op(n6536) );
  nor2_1 U6877 ( .ip1(n6533), .ip2(n8029), .op(n6535) );
  nand2_1 U6878 ( .ip1(n7045), .ip2(column[23]), .op(n6534) );
  nand2_1 U6879 ( .ip1(n7045), .ip2(column[24]), .op(n6626) );
  fulladder U6880 ( .a(n6536), .b(n6535), .ci(n6534), .co(n6627), .s(n6553) );
  nand2_1 U6881 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[23]), .op(n6559)
         );
  nor2_1 U6882 ( .ip1(n6536), .ip2(n6559), .op(n6541) );
  nand2_1 U6883 ( .ip1(n7882), .ip2(m1Inputs[23]), .op(n6545) );
  or2_1 U6884 ( .ip1(n6545), .ip2(n6541), .op(n6539) );
  nand2_1 U6885 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[24]), .op(n6537)
         );
  or2_1 U6886 ( .ip1(n6537), .ip2(n6541), .op(n6538) );
  nand2_1 U6887 ( .ip1(n6539), .ip2(n6538), .op(n6543) );
  and3_1 U6888 ( .ip1(n8051), .ip2(column[22]), .ip3(n6543), .op(n6540) );
  nor2_1 U6889 ( .ip1(n6541), .ip2(n6540), .op(n6552) );
  nand2_1 U6890 ( .ip1(n7045), .ip2(column[22]), .op(n6542) );
  xor2_1 U6891 ( .ip1(n6543), .ip2(n6542), .op(n6556) );
  nor2_1 U6892 ( .ip1(n6544), .ip2(n8029), .op(n6555) );
  nor2_1 U6893 ( .ip1(n6545), .ip2(n6560), .op(n6550) );
  or2_1 U6894 ( .ip1(n6559), .ip2(n6550), .op(n6548) );
  nand2_1 U6895 ( .ip1(n7882), .ip2(m1Inputs[22]), .op(n6546) );
  or2_1 U6896 ( .ip1(n6546), .ip2(n6550), .op(n6547) );
  nand2_1 U6897 ( .ip1(n6548), .ip2(n6547), .op(n6569) );
  and3_1 U6898 ( .ip1(n8051), .ip2(column[21]), .ip3(n6569), .op(n6549) );
  nor2_1 U6899 ( .ip1(n6550), .ip2(n6549), .op(n6554) );
  fulladder U6900 ( .a(n6553), .b(n6552), .ci(n6551), .co(n6655), .s(n6660) );
  fulladder U6901 ( .a(n6556), .b(n6555), .ci(n6554), .co(n6551), .s(n6576) );
  nand2_1 U6902 ( .ip1(n8064), .ip2(m1Inputs[24]), .op(n6572) );
  nor2_1 U6903 ( .ip1(n6557), .ip2(n8029), .op(n6571) );
  nor2_1 U6904 ( .ip1(n6559), .ip2(n6558), .op(n6564) );
  or2_1 U6905 ( .ip1(n6560), .ip2(n6564), .op(n6563) );
  nand2_1 U6906 ( .ip1(n8064), .ip2(m1Inputs[23]), .op(n6561) );
  or2_1 U6907 ( .ip1(n6561), .ip2(n6564), .op(n6562) );
  nand2_1 U6908 ( .ip1(n6563), .ip2(n6562), .op(n6590) );
  or2_1 U6909 ( .ip1(n6590), .ip2(n6564), .op(n6567) );
  nand2_1 U6910 ( .ip1(n7045), .ip2(column[20]), .op(n6589) );
  inv_1 U6911 ( .ip(n6589), .op(n6565) );
  or2_1 U6912 ( .ip1(n6565), .ip2(n6564), .op(n6566) );
  nand2_1 U6913 ( .ip1(n6567), .ip2(n6566), .op(n6570) );
  nand2_1 U6914 ( .ip1(n7045), .ip2(column[21]), .op(n6568) );
  xor2_1 U6915 ( .ip1(n6569), .ip2(n6568), .op(n6579) );
  fulladder U6916 ( .a(n6572), .b(n6571), .ci(n6570), .co(n6575), .s(n6578) );
  nor2_1 U6917 ( .ip1(n6573), .ip2(n8029), .op(n6593) );
  nand2_1 U6918 ( .ip1(n7882), .ip2(m1Inputs[21]), .op(n6592) );
  nand2_1 U6919 ( .ip1(n8078), .ip2(m1Inputs[24]), .op(n6591) );
  fulladder U6920 ( .a(n6576), .b(n6575), .ci(n6574), .co(n6659), .s(n6664) );
  fulladder U6921 ( .a(n6579), .b(n6578), .ci(n6577), .co(n6574), .s(n6602) );
  or2_1 U6922 ( .ip1(n6580), .ip2(n6582), .op(n6585) );
  inv_1 U6923 ( .ip(n6581), .op(n6583) );
  or2_1 U6924 ( .ip1(n6583), .ip2(n6582), .op(n6584) );
  nand2_1 U6925 ( .ip1(n6585), .ip2(n6584), .op(n6596) );
  fulladder U6926 ( .a(n6588), .b(n6587), .ci(n6586), .co(n6595), .s(n6607) );
  xor2_1 U6927 ( .ip1(n6590), .ip2(n6589), .op(n6594) );
  fulladder U6928 ( .a(n6593), .b(n6592), .ci(n6591), .co(n6577), .s(n6605) );
  fulladder U6929 ( .a(n6596), .b(n6595), .ci(n6594), .co(n6601), .s(n6604) );
  fulladder U6930 ( .a(n6599), .b(n6598), .ci(n6597), .co(n6603), .s(n6505) );
  fulladder U6931 ( .a(n6602), .b(n6601), .ci(n6600), .co(n6663), .s(n6668) );
  fulladder U6932 ( .a(n6605), .b(n6604), .ci(n6603), .co(n6600), .s(n6606) );
  inv_1 U6933 ( .ip(n6606), .op(n6617) );
  fulladder U6934 ( .a(n6609), .b(n6608), .ci(n6607), .co(n6610), .s(n6513) );
  inv_1 U6935 ( .ip(n6610), .op(n6616) );
  fulladder U6936 ( .a(n6613), .b(n6612), .ci(n6611), .co(n6615), .s(n6517) );
  inv_1 U6937 ( .ip(n6614), .op(n6667) );
  fulladder U6938 ( .a(n6617), .b(n6616), .ci(n6615), .co(n6614), .s(n6618) );
  inv_1 U6939 ( .ip(n6618), .op(n6672) );
  fulladder U6940 ( .a(n6621), .b(n6620), .ci(n6619), .co(n6622), .s(
        \STAGE_1/M2/sum [3]) );
  inv_1 U6941 ( .ip(n6622), .op(n6671) );
  fulladder U6942 ( .a(n6625), .b(n6624), .ci(n6623), .co(n6670), .s(n6525) );
  fulladder U6943 ( .a(n6628), .b(n6627), .ci(n6626), .co(n6647), .s(n6656) );
  nand2_1 U6944 ( .ip1(n7045), .ip2(column[25]), .op(n6652) );
  nor3_1 U6945 ( .ip1(n6648), .ip2(n6647), .ip3(n6652), .op(n6642) );
  nand2_1 U6946 ( .ip1(column[26]), .ip2(n6642), .op(n6637) );
  nor2_1 U6947 ( .ip1(n6640), .ip2(n6637), .op(n6631) );
  nand2_1 U6948 ( .ip1(column[28]), .ip2(n6631), .op(n6675) );
  and2_1 U6949 ( .ip1(n8051), .ip2(column[28]), .op(n6635) );
  and2_1 U6950 ( .ip1(n8051), .ip2(column[26]), .op(n6646) );
  nand3_1 U6951 ( .ip1(n6648), .ip2(n6647), .ip3(n6652), .op(n6643) );
  nor2_1 U6952 ( .ip1(n6646), .ip2(n6643), .op(n6636) );
  nand2_1 U6953 ( .ip1(n6636), .ip2(n6640), .op(n6632) );
  nor2_1 U6954 ( .ip1(n6635), .ip2(n6632), .op(n6674) );
  inv_1 U6955 ( .ip(n6674), .op(n6629) );
  nand2_1 U6956 ( .ip1(n6675), .ip2(n6629), .op(n6630) );
  xor2_1 U6957 ( .ip1(n6679), .ip2(n6630), .op(\STAGE_1/M2/sum [13]) );
  inv_1 U6958 ( .ip(n6631), .op(n6633) );
  nand2_1 U6959 ( .ip1(n6633), .ip2(n6632), .op(n6634) );
  xor2_1 U6960 ( .ip1(n6635), .ip2(n6634), .op(\STAGE_1/M2/sum [12]) );
  inv_1 U6961 ( .ip(n6640), .op(n6641) );
  inv_1 U6962 ( .ip(n6636), .op(n6638) );
  nand2_1 U6963 ( .ip1(n6638), .ip2(n6637), .op(n6639) );
  mux2_1 U6964 ( .ip1(n6641), .ip2(n6640), .s(n6639), .op(\STAGE_1/M2/sum [11]) );
  inv_1 U6965 ( .ip(n6642), .op(n6644) );
  nand2_1 U6966 ( .ip1(n6644), .ip2(n6643), .op(n6645) );
  xor2_1 U6967 ( .ip1(n6646), .ip2(n6645), .op(\STAGE_1/M2/sum [10]) );
  inv_1 U6968 ( .ip(n6652), .op(n6653) );
  nand2_1 U6969 ( .ip1(n6648), .ip2(n6647), .op(n6650) );
  or2_1 U6970 ( .ip1(n6648), .ip2(n6647), .op(n6649) );
  nand2_1 U6971 ( .ip1(n6650), .ip2(n6649), .op(n6651) );
  mux2_1 U6972 ( .ip1(n6653), .ip2(n6652), .s(n6651), .op(\STAGE_1/M2/sum [9])
         );
  fulladder U6973 ( .a(n6656), .b(n6655), .ci(n6654), .co(n6648), .s(n6657) );
  inv_1 U6974 ( .ip(n6657), .op(\STAGE_1/M2/sum [8]) );
  fulladder U6975 ( .a(n6660), .b(n6659), .ci(n6658), .co(n6654), .s(n6661) );
  inv_1 U6976 ( .ip(n6661), .op(\STAGE_1/M2/sum [7]) );
  fulladder U6977 ( .a(n6664), .b(n6663), .ci(n6662), .co(n6658), .s(n6665) );
  inv_1 U6978 ( .ip(n6665), .op(\STAGE_1/M2/sum [6]) );
  fulladder U6979 ( .a(n6668), .b(n6667), .ci(n6666), .co(n6662), .s(n6669) );
  inv_1 U6980 ( .ip(n6669), .op(\STAGE_1/M2/sum [5]) );
  fulladder U6981 ( .a(n6672), .b(n6671), .ci(n6670), .co(n6666), .s(n6673) );
  inv_1 U6982 ( .ip(n6673), .op(\STAGE_1/M2/sum [4]) );
  nand2_1 U6983 ( .ip1(n7045), .ip2(column[30]), .op(n6680) );
  or2_1 U6984 ( .ip1(n6679), .ip2(n6674), .op(n6676) );
  nand2_1 U6985 ( .ip1(n6676), .ip2(n6675), .op(n6678) );
  nor2_1 U6986 ( .ip1(column[30]), .ip2(column[31]), .op(n6677) );
  not_ab_or_c_or_d U6987 ( .ip1(column[30]), .ip2(column[31]), .ip3(n6677), 
        .ip4(n8180), .op(n6682) );
  fulladder U6988 ( .a(n6680), .b(n6679), .ci(n6678), .co(n6681), .s(
        \STAGE_1/M2/sum [14]) );
  xnor2_1 U6989 ( .ip1(n6682), .ip2(n6681), .op(\STAGE_1/M2/sum [15]) );
  nand2_1 U6990 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[39]), .op(n6788)
         );
  nor2_1 U6991 ( .ip1(n6684), .ip2(n6683), .op(n6685) );
  nor2_1 U6992 ( .ip1(n6686), .ip2(n6685), .op(n6787) );
  fulladder U6993 ( .a(n6689), .b(n6688), .ci(n6687), .co(n6786), .s(n5773) );
  inv_1 U6994 ( .ip(n6690), .op(n6802) );
  nand2_1 U6995 ( .ip1(n7882), .ip2(m1Inputs[36]), .op(n6776) );
  nor2_1 U6996 ( .ip1(n6691), .ip2(n8029), .op(n6775) );
  nand2_1 U6997 ( .ip1(n8001), .ip2(m1Inputs[40]), .op(n6774) );
  fulladder U6998 ( .a(n6694), .b(n6693), .ci(n6692), .co(n6797), .s(n5779) );
  nand2_1 U6999 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[38]), .op(n6742)
         );
  nor3_1 U7000 ( .ip1(n7813), .ip2(n6742), .ip3(n6749), .op(n6770) );
  or2_1 U7001 ( .ip1(n6740), .ip2(n6770), .op(n6697) );
  nand2_1 U7002 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[37]), .op(n6695)
         );
  or2_1 U7003 ( .ip1(n6695), .ip2(n6770), .op(n6696) );
  nand2_1 U7004 ( .ip1(n6697), .ip2(n6696), .op(n6768) );
  nand2_1 U7005 ( .ip1(n7045), .ip2(column[35]), .op(n6769) );
  xor2_1 U7006 ( .ip1(n6768), .ip2(n6769), .op(n6796) );
  inv_1 U7007 ( .ip(n6698), .op(n6801) );
  fulladder U7008 ( .a(n6701), .b(n6700), .ci(n6699), .co(n6800), .s(n5793) );
  inv_1 U7009 ( .ip(n6702), .op(n6814) );
  fulladder U7010 ( .a(n6705), .b(n6704), .ci(n6703), .co(n6706), .s(n6713) );
  inv_1 U7011 ( .ip(n6706), .op(n6813) );
  fulladder U7012 ( .a(n6709), .b(n6708), .ci(n6707), .co(n6812), .s(n5798) );
  inv_1 U7013 ( .ip(n6710), .op(n6810) );
  fulladder U7014 ( .a(n6713), .b(n6712), .ci(n6711), .co(n6809), .s(n6716) );
  fulladder U7015 ( .a(n6716), .b(n6715), .ci(n6714), .co(n6808), .s(
        \STAGE_1/M3/sum [2]) );
  and2_1 U7016 ( .ip1(n8051), .ip2(column[45]), .op(n6867) );
  nor2_1 U7017 ( .ip1(n6748), .ip2(n8029), .op(n6817) );
  nand2_1 U7018 ( .ip1(n7882), .ip2(m1Inputs[40]), .op(n6720) );
  nor2_1 U7019 ( .ip1(n6717), .ip2(n8029), .op(n6719) );
  nand2_1 U7020 ( .ip1(n7045), .ip2(column[39]), .op(n6718) );
  nand2_1 U7021 ( .ip1(n7045), .ip2(column[40]), .op(n6815) );
  fulladder U7022 ( .a(n6720), .b(n6719), .ci(n6718), .co(n6816), .s(n6736) );
  nand2_1 U7023 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[39]), .op(n6741)
         );
  nor2_1 U7024 ( .ip1(n6720), .ip2(n6741), .op(n6725) );
  nand2_1 U7025 ( .ip1(n8037), .ip2(m1Inputs[40]), .op(n6721) );
  or2_1 U7026 ( .ip1(n6721), .ip2(n6725), .op(n6723) );
  nand2_1 U7027 ( .ip1(n7882), .ip2(m1Inputs[39]), .op(n6729) );
  or2_1 U7028 ( .ip1(n6729), .ip2(n6725), .op(n6722) );
  nand2_1 U7029 ( .ip1(n6723), .ip2(n6722), .op(n6727) );
  and3_1 U7030 ( .ip1(n8051), .ip2(column[38]), .ip3(n6727), .op(n6724) );
  nor2_1 U7031 ( .ip1(n6725), .ip2(n6724), .op(n6735) );
  nand2_1 U7032 ( .ip1(n7045), .ip2(column[38]), .op(n6726) );
  xor2_1 U7033 ( .ip1(n6727), .ip2(n6726), .op(n6739) );
  nor2_1 U7034 ( .ip1(n6728), .ip2(n7628), .op(n6738) );
  nor2_1 U7035 ( .ip1(n6729), .ip2(n6742), .op(n6733) );
  or2_1 U7036 ( .ip1(n6741), .ip2(n6733), .op(n6732) );
  nand2_1 U7037 ( .ip1(n7882), .ip2(m1Inputs[38]), .op(n6730) );
  or2_1 U7038 ( .ip1(n6730), .ip2(n6733), .op(n6731) );
  nand2_1 U7039 ( .ip1(n6732), .ip2(n6731), .op(n6754) );
  and3_1 U7040 ( .ip1(n8051), .ip2(column[37]), .ip3(n6754), .op(n6756) );
  nor2_1 U7041 ( .ip1(n6733), .ip2(n6756), .op(n6737) );
  fulladder U7042 ( .a(n6736), .b(n6735), .ci(n6734), .co(n6843), .s(n6848) );
  fulladder U7043 ( .a(n6739), .b(n6738), .ci(n6737), .co(n6734), .s(n6763) );
  nand2_1 U7044 ( .ip1(n8064), .ip2(m1Inputs[40]), .op(n6752) );
  nor2_1 U7045 ( .ip1(n6749), .ip2(n8029), .op(n6751) );
  nor2_1 U7046 ( .ip1(n6741), .ip2(n6740), .op(n6747) );
  or2_1 U7047 ( .ip1(n6742), .ip2(n6747), .op(n6745) );
  or2_1 U7048 ( .ip1(n6743), .ip2(n6747), .op(n6744) );
  nand2_1 U7049 ( .ip1(n6745), .ip2(n6744), .op(n6778) );
  and3_1 U7050 ( .ip1(n8051), .ip2(column[36]), .ip3(n6778), .op(n6746) );
  nor2_1 U7051 ( .ip1(n6747), .ip2(n6746), .op(n6750) );
  nor2_1 U7052 ( .ip1(n5060), .ip2(n6748), .op(n6781) );
  nor2_1 U7053 ( .ip1(n7685), .ip2(n6749), .op(n6780) );
  nand2_1 U7054 ( .ip1(m1Inputs[36]), .ip2(\STAGE_1/weightReg [15]), .op(n6779) );
  fulladder U7055 ( .a(n6752), .b(n6751), .ci(n6750), .co(n6762), .s(n6753) );
  inv_1 U7056 ( .ip(n6753), .op(n6765) );
  inv_1 U7057 ( .ip(n6754), .op(n6755) );
  or2_1 U7058 ( .ip1(n6755), .ip2(n6756), .op(n6759) );
  nand2_1 U7059 ( .ip1(n7045), .ip2(column[37]), .op(n6757) );
  or2_1 U7060 ( .ip1(n6757), .ip2(n6756), .op(n6758) );
  nand2_1 U7061 ( .ip1(n6759), .ip2(n6758), .op(n6764) );
  inv_1 U7062 ( .ip(n6760), .op(n6761) );
  fulladder U7063 ( .a(n6763), .b(n6762), .ci(n6761), .co(n6847), .s(n6852) );
  fulladder U7064 ( .a(n6766), .b(n6765), .ci(n6764), .co(n6760), .s(n6767) );
  inv_1 U7065 ( .ip(n6767), .op(n6791) );
  or2_1 U7066 ( .ip1(n6768), .ip2(n6770), .op(n6773) );
  inv_1 U7067 ( .ip(n6769), .op(n6771) );
  or2_1 U7068 ( .ip1(n6771), .ip2(n6770), .op(n6772) );
  nand2_1 U7069 ( .ip1(n6773), .ip2(n6772), .op(n6785) );
  fulladder U7070 ( .a(n6776), .b(n6775), .ci(n6774), .co(n6784), .s(n6798) );
  nand2_1 U7071 ( .ip1(n7045), .ip2(column[36]), .op(n6777) );
  xor2_1 U7072 ( .ip1(n6778), .ip2(n6777), .op(n6783) );
  fulladder U7073 ( .a(n6781), .b(n6780), .ci(n6779), .co(n6766), .s(n6782) );
  inv_1 U7074 ( .ip(n6782), .op(n6794) );
  fulladder U7075 ( .a(n6785), .b(n6784), .ci(n6783), .co(n6790), .s(n6793) );
  fulladder U7076 ( .a(n6788), .b(n6787), .ci(n6786), .co(n6792), .s(n6690) );
  fulladder U7077 ( .a(n6791), .b(n6790), .ci(n6789), .co(n6851), .s(n6856) );
  fulladder U7078 ( .a(n6794), .b(n6793), .ci(n6792), .co(n6789), .s(n6795) );
  inv_1 U7079 ( .ip(n6795), .op(n6806) );
  fulladder U7080 ( .a(n6798), .b(n6797), .ci(n6796), .co(n6799), .s(n6698) );
  inv_1 U7081 ( .ip(n6799), .op(n6805) );
  fulladder U7082 ( .a(n6802), .b(n6801), .ci(n6800), .co(n6804), .s(n6702) );
  inv_1 U7083 ( .ip(n6803), .op(n6855) );
  fulladder U7084 ( .a(n6806), .b(n6805), .ci(n6804), .co(n6803), .s(n6807) );
  inv_1 U7085 ( .ip(n6807), .op(n6860) );
  fulladder U7086 ( .a(n6810), .b(n6809), .ci(n6808), .co(n6811), .s(
        \STAGE_1/M3/sum [3]) );
  inv_1 U7087 ( .ip(n6811), .op(n6859) );
  fulladder U7088 ( .a(n6814), .b(n6813), .ci(n6812), .co(n6858), .s(n6710) );
  fulladder U7089 ( .a(n6817), .b(n6816), .ci(n6815), .co(n6835), .s(n6844) );
  nand2_1 U7090 ( .ip1(n7045), .ip2(column[41]), .op(n6840) );
  nor3_1 U7091 ( .ip1(n6836), .ip2(n6835), .ip3(n6840), .op(n6831) );
  nand2_1 U7092 ( .ip1(n7045), .ip2(column[43]), .op(n6830) );
  inv_1 U7093 ( .ip(n6830), .op(n6829) );
  nand3_1 U7094 ( .ip1(column[42]), .ip2(n6831), .ip3(n6829), .op(n6822) );
  inv_1 U7095 ( .ip(n6822), .op(n6818) );
  nand2_1 U7096 ( .ip1(column[44]), .ip2(n6818), .op(n6863) );
  and2_1 U7097 ( .ip1(n8051), .ip2(column[44]), .op(n6824) );
  nand2_1 U7098 ( .ip1(n7045), .ip2(column[42]), .op(n6834) );
  and4_1 U7099 ( .ip1(n6836), .ip2(n6835), .ip3(n6834), .ip4(n6840), .op(n6825) );
  nand2_1 U7100 ( .ip1(n6825), .ip2(n6830), .op(n6821) );
  nor2_1 U7101 ( .ip1(n6824), .ip2(n6821), .op(n6862) );
  inv_1 U7102 ( .ip(n6862), .op(n6819) );
  nand2_1 U7103 ( .ip1(n6863), .ip2(n6819), .op(n6820) );
  xor2_1 U7104 ( .ip1(n6867), .ip2(n6820), .op(\STAGE_1/M3/sum [13]) );
  nand2_1 U7105 ( .ip1(n6822), .ip2(n6821), .op(n6823) );
  xor2_1 U7106 ( .ip1(n6824), .ip2(n6823), .op(\STAGE_1/M3/sum [12]) );
  or2_1 U7107 ( .ip1(column[42]), .ip2(n6825), .op(n6827) );
  or2_1 U7108 ( .ip1(n6831), .ip2(n6825), .op(n6826) );
  nand2_1 U7109 ( .ip1(n6827), .ip2(n6826), .op(n6828) );
  mux2_1 U7110 ( .ip1(n6830), .ip2(n6829), .s(n6828), .op(\STAGE_1/M3/sum [11]) );
  and3_1 U7111 ( .ip1(n6836), .ip2(n6835), .ip3(n6840), .op(n6832) );
  nor2_1 U7112 ( .ip1(n6832), .ip2(n6831), .op(n6833) );
  xor2_1 U7113 ( .ip1(n6834), .ip2(n6833), .op(\STAGE_1/M3/sum [10]) );
  inv_1 U7114 ( .ip(n6840), .op(n6841) );
  nand2_1 U7115 ( .ip1(n6836), .ip2(n6835), .op(n6838) );
  or2_1 U7116 ( .ip1(n6836), .ip2(n6835), .op(n6837) );
  nand2_1 U7117 ( .ip1(n6838), .ip2(n6837), .op(n6839) );
  mux2_1 U7118 ( .ip1(n6841), .ip2(n6840), .s(n6839), .op(\STAGE_1/M3/sum [9])
         );
  fulladder U7119 ( .a(n6844), .b(n6843), .ci(n6842), .co(n6836), .s(n6845) );
  inv_1 U7120 ( .ip(n6845), .op(\STAGE_1/M3/sum [8]) );
  fulladder U7121 ( .a(n6848), .b(n6847), .ci(n6846), .co(n6842), .s(n6849) );
  inv_1 U7122 ( .ip(n6849), .op(\STAGE_1/M3/sum [7]) );
  fulladder U7123 ( .a(n6852), .b(n6851), .ci(n6850), .co(n6846), .s(n6853) );
  inv_1 U7124 ( .ip(n6853), .op(\STAGE_1/M3/sum [6]) );
  fulladder U7125 ( .a(n6856), .b(n6855), .ci(n6854), .co(n6850), .s(n6857) );
  inv_1 U7126 ( .ip(n6857), .op(\STAGE_1/M3/sum [5]) );
  fulladder U7127 ( .a(n6860), .b(n6859), .ci(n6858), .co(n6854), .s(n6861) );
  inv_1 U7128 ( .ip(n6861), .op(\STAGE_1/M3/sum [4]) );
  nand2_1 U7129 ( .ip1(n7045), .ip2(column[46]), .op(n6868) );
  or2_1 U7130 ( .ip1(n6867), .ip2(n6862), .op(n6864) );
  nand2_1 U7131 ( .ip1(n6864), .ip2(n6863), .op(n6866) );
  nor2_1 U7132 ( .ip1(column[46]), .ip2(column[47]), .op(n6865) );
  not_ab_or_c_or_d U7133 ( .ip1(column[46]), .ip2(column[47]), .ip3(n6865), 
        .ip4(n8180), .op(n6870) );
  fulladder U7134 ( .a(n6868), .b(n6867), .ci(n6866), .co(n6869), .s(
        \STAGE_1/M3/sum [14]) );
  xnor2_1 U7135 ( .ip1(n6870), .ip2(n6869), .op(\STAGE_1/M3/sum [15]) );
  nand2_1 U7136 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[55]), .op(n6973)
         );
  inv_1 U7137 ( .ip(n6871), .op(n6875) );
  nor2_1 U7138 ( .ip1(n6873), .ip2(n6872), .op(n6874) );
  nor2_1 U7139 ( .ip1(n6875), .ip2(n6874), .op(n6972) );
  fulladder U7140 ( .a(n6878), .b(n6877), .ci(n6876), .co(n6971), .s(n5845) );
  inv_1 U7141 ( .ip(n6879), .op(n6987) );
  nand2_1 U7142 ( .ip1(n8064), .ip2(m1Inputs[54]), .op(n6932) );
  nand2_1 U7143 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[54]), .op(n6934)
         );
  nor3_1 U7144 ( .ip1(n7813), .ip2(n6934), .ip3(n6931), .op(n6956) );
  or2_1 U7145 ( .ip1(n6932), .ip2(n6956), .op(n6882) );
  nand2_1 U7146 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[53]), .op(n6880)
         );
  or2_1 U7147 ( .ip1(n6880), .ip2(n6956), .op(n6881) );
  nand2_1 U7148 ( .ip1(n6882), .ip2(n6881), .op(n6954) );
  nand2_1 U7149 ( .ip1(n8009), .ip2(column[51]), .op(n6955) );
  xor2_1 U7150 ( .ip1(n6954), .ip2(n6955), .op(n6983) );
  fulladder U7151 ( .a(n6885), .b(n6884), .ci(n6883), .co(n6982), .s(n5851) );
  nand2_1 U7152 ( .ip1(n7882), .ip2(m1Inputs[52]), .op(n6962) );
  nor2_1 U7153 ( .ip1(n6886), .ip2(n8029), .op(n6961) );
  nand2_1 U7154 ( .ip1(n8001), .ip2(m1Inputs[56]), .op(n6960) );
  inv_1 U7155 ( .ip(n6887), .op(n6986) );
  fulladder U7156 ( .a(n6890), .b(n6889), .ci(n6888), .co(n6985), .s(n5864) );
  inv_1 U7157 ( .ip(n6891), .op(n6999) );
  fulladder U7158 ( .a(n6894), .b(n6893), .ci(n6892), .co(n6895), .s(n6902) );
  inv_1 U7159 ( .ip(n6895), .op(n6998) );
  fulladder U7160 ( .a(n6898), .b(n6897), .ci(n6896), .co(n6997), .s(n5869) );
  inv_1 U7161 ( .ip(n6899), .op(n6995) );
  fulladder U7162 ( .a(n6902), .b(n6901), .ci(n6900), .co(n6994), .s(n6905) );
  fulladder U7163 ( .a(n6905), .b(n6904), .ci(n6903), .co(n6993), .s(
        \STAGE_1/M4/sum [2]) );
  and2_1 U7164 ( .ip1(n8051), .ip2(column[60]), .op(n7048) );
  nor2_1 U7165 ( .ip1(n6906), .ip2(n7628), .op(n7002) );
  nand2_1 U7166 ( .ip1(n7882), .ip2(m1Inputs[56]), .op(n6910) );
  nor2_1 U7167 ( .ip1(n6907), .ip2(n7628), .op(n6909) );
  nand2_1 U7168 ( .ip1(n8009), .ip2(column[55]), .op(n6908) );
  nand2_1 U7169 ( .ip1(n8009), .ip2(column[56]), .op(n7000) );
  fulladder U7170 ( .a(n6910), .b(n6909), .ci(n6908), .co(n7001), .s(n6927) );
  nand2_1 U7171 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[55]), .op(n6933)
         );
  nor2_1 U7172 ( .ip1(n6910), .ip2(n6933), .op(n6915) );
  nand2_1 U7173 ( .ip1(\STAGE_1/weightReg [7]), .ip2(m1Inputs[55]), .op(n6919)
         );
  or2_1 U7174 ( .ip1(n6919), .ip2(n6915), .op(n6913) );
  nand2_1 U7175 ( .ip1(n8037), .ip2(m1Inputs[56]), .op(n6911) );
  or2_1 U7176 ( .ip1(n6911), .ip2(n6915), .op(n6912) );
  nand2_1 U7177 ( .ip1(n6913), .ip2(n6912), .op(n6917) );
  and3_1 U7178 ( .ip1(n8051), .ip2(column[54]), .ip3(n6917), .op(n6914) );
  nor2_1 U7179 ( .ip1(n6915), .ip2(n6914), .op(n6926) );
  nand2_1 U7180 ( .ip1(n7045), .ip2(column[54]), .op(n6916) );
  xor2_1 U7181 ( .ip1(n6917), .ip2(n6916), .op(n6930) );
  nor2_1 U7182 ( .ip1(n6918), .ip2(n7628), .op(n6929) );
  nor2_1 U7183 ( .ip1(n6919), .ip2(n6934), .op(n6924) );
  or2_1 U7184 ( .ip1(n6933), .ip2(n6924), .op(n6922) );
  nand2_1 U7185 ( .ip1(n7882), .ip2(m1Inputs[54]), .op(n6920) );
  or2_1 U7186 ( .ip1(n6920), .ip2(n6924), .op(n6921) );
  nand2_1 U7187 ( .ip1(n6922), .ip2(n6921), .op(n6943) );
  and3_1 U7188 ( .ip1(n8051), .ip2(column[53]), .ip3(n6943), .op(n6923) );
  nor2_1 U7189 ( .ip1(n6924), .ip2(n6923), .op(n6928) );
  fulladder U7190 ( .a(n6927), .b(n6926), .ci(n6925), .co(n7023), .s(n7028) );
  fulladder U7191 ( .a(n6930), .b(n6929), .ci(n6928), .co(n6925), .s(n6950) );
  nand2_1 U7192 ( .ip1(n8064), .ip2(m1Inputs[56]), .op(n6946) );
  nor2_1 U7193 ( .ip1(n6931), .ip2(n8029), .op(n6945) );
  nor2_1 U7194 ( .ip1(n6933), .ip2(n6932), .op(n6938) );
  or2_1 U7195 ( .ip1(n6934), .ip2(n6938), .op(n6937) );
  nand2_1 U7196 ( .ip1(n8064), .ip2(m1Inputs[55]), .op(n6935) );
  or2_1 U7197 ( .ip1(n6935), .ip2(n6938), .op(n6936) );
  nand2_1 U7198 ( .ip1(n6937), .ip2(n6936), .op(n6964) );
  or2_1 U7199 ( .ip1(n6964), .ip2(n6938), .op(n6941) );
  nand2_1 U7200 ( .ip1(n7045), .ip2(column[52]), .op(n6963) );
  inv_1 U7201 ( .ip(n6963), .op(n6939) );
  or2_1 U7202 ( .ip1(n6939), .ip2(n6938), .op(n6940) );
  nand2_1 U7203 ( .ip1(n6941), .ip2(n6940), .op(n6944) );
  nand2_1 U7204 ( .ip1(n7045), .ip2(column[53]), .op(n6942) );
  xor2_1 U7205 ( .ip1(n6943), .ip2(n6942), .op(n6953) );
  fulladder U7206 ( .a(n6946), .b(n6945), .ci(n6944), .co(n6949), .s(n6952) );
  nor2_1 U7207 ( .ip1(n6947), .ip2(n8029), .op(n6967) );
  nand2_1 U7208 ( .ip1(n7882), .ip2(m1Inputs[53]), .op(n6966) );
  nand2_1 U7209 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[56]), .op(n6965)
         );
  fulladder U7210 ( .a(n6950), .b(n6949), .ci(n6948), .co(n7027), .s(n7032) );
  fulladder U7211 ( .a(n6953), .b(n6952), .ci(n6951), .co(n6948), .s(n6976) );
  or2_1 U7212 ( .ip1(n6954), .ip2(n6956), .op(n6959) );
  inv_1 U7213 ( .ip(n6955), .op(n6957) );
  or2_1 U7214 ( .ip1(n6957), .ip2(n6956), .op(n6958) );
  nand2_1 U7215 ( .ip1(n6959), .ip2(n6958), .op(n6970) );
  fulladder U7216 ( .a(n6962), .b(n6961), .ci(n6960), .co(n6969), .s(n6981) );
  xor2_1 U7217 ( .ip1(n6964), .ip2(n6963), .op(n6968) );
  fulladder U7218 ( .a(n6967), .b(n6966), .ci(n6965), .co(n6951), .s(n6979) );
  fulladder U7219 ( .a(n6970), .b(n6969), .ci(n6968), .co(n6975), .s(n6978) );
  fulladder U7220 ( .a(n6973), .b(n6972), .ci(n6971), .co(n6977), .s(n6879) );
  fulladder U7221 ( .a(n6976), .b(n6975), .ci(n6974), .co(n7031), .s(n7036) );
  fulladder U7222 ( .a(n6979), .b(n6978), .ci(n6977), .co(n6974), .s(n6980) );
  inv_1 U7223 ( .ip(n6980), .op(n6991) );
  fulladder U7224 ( .a(n6983), .b(n6982), .ci(n6981), .co(n6984), .s(n6887) );
  inv_1 U7225 ( .ip(n6984), .op(n6990) );
  fulladder U7226 ( .a(n6987), .b(n6986), .ci(n6985), .co(n6989), .s(n6891) );
  inv_1 U7227 ( .ip(n6988), .op(n7035) );
  fulladder U7228 ( .a(n6991), .b(n6990), .ci(n6989), .co(n6988), .s(n6992) );
  inv_1 U7229 ( .ip(n6992), .op(n7040) );
  fulladder U7230 ( .a(n6995), .b(n6994), .ci(n6993), .co(n6996), .s(
        \STAGE_1/M4/sum [3]) );
  inv_1 U7231 ( .ip(n6996), .op(n7039) );
  fulladder U7232 ( .a(n6999), .b(n6998), .ci(n6997), .co(n7038), .s(n6899) );
  fulladder U7233 ( .a(n7002), .b(n7001), .ci(n7000), .co(n7015), .s(n7024) );
  nand2_1 U7234 ( .ip1(n8009), .ip2(column[57]), .op(n7020) );
  inv_1 U7235 ( .ip(column[58]), .op(n7003) );
  nor4_1 U7236 ( .ip1(n7016), .ip2(n7015), .ip3(n7020), .ip4(n7003), .op(n7006) );
  nand2_1 U7237 ( .ip1(column[59]), .ip2(n7006), .op(n7043) );
  and2_1 U7238 ( .ip1(n8051), .ip2(column[59]), .op(n7010) );
  nand2_1 U7239 ( .ip1(n8009), .ip2(column[58]), .op(n7014) );
  nand4_1 U7240 ( .ip1(n7016), .ip2(n7015), .ip3(n7014), .ip4(n7020), .op(
        n7007) );
  nor2_1 U7241 ( .ip1(n7010), .ip2(n7007), .op(n7042) );
  inv_1 U7242 ( .ip(n7042), .op(n7004) );
  nand2_1 U7243 ( .ip1(n7043), .ip2(n7004), .op(n7005) );
  xor2_1 U7244 ( .ip1(n7048), .ip2(n7005), .op(\STAGE_1/M4/sum [12]) );
  inv_1 U7245 ( .ip(n7006), .op(n7008) );
  nand2_1 U7246 ( .ip1(n7008), .ip2(n7007), .op(n7009) );
  xor2_1 U7247 ( .ip1(n7010), .ip2(n7009), .op(\STAGE_1/M4/sum [11]) );
  and3_1 U7248 ( .ip1(n7016), .ip2(n7015), .ip3(n7020), .op(n7012) );
  nor3_1 U7249 ( .ip1(n7016), .ip2(n7015), .ip3(n7020), .op(n7011) );
  nor2_1 U7250 ( .ip1(n7012), .ip2(n7011), .op(n7013) );
  xor2_1 U7251 ( .ip1(n7014), .ip2(n7013), .op(\STAGE_1/M4/sum [10]) );
  inv_1 U7252 ( .ip(n7020), .op(n7021) );
  nand2_1 U7253 ( .ip1(n7016), .ip2(n7015), .op(n7018) );
  or2_1 U7254 ( .ip1(n7016), .ip2(n7015), .op(n7017) );
  nand2_1 U7255 ( .ip1(n7018), .ip2(n7017), .op(n7019) );
  mux2_1 U7256 ( .ip1(n7021), .ip2(n7020), .s(n7019), .op(\STAGE_1/M4/sum [9])
         );
  fulladder U7257 ( .a(n7024), .b(n7023), .ci(n7022), .co(n7016), .s(n7025) );
  inv_1 U7258 ( .ip(n7025), .op(\STAGE_1/M4/sum [8]) );
  fulladder U7259 ( .a(n7028), .b(n7027), .ci(n7026), .co(n7022), .s(n7029) );
  inv_1 U7260 ( .ip(n7029), .op(\STAGE_1/M4/sum [7]) );
  fulladder U7261 ( .a(n7032), .b(n7031), .ci(n7030), .co(n7026), .s(n7033) );
  inv_1 U7262 ( .ip(n7033), .op(\STAGE_1/M4/sum [6]) );
  fulladder U7263 ( .a(n7036), .b(n7035), .ci(n7034), .co(n7030), .s(n7037) );
  inv_1 U7264 ( .ip(n7037), .op(\STAGE_1/M4/sum [5]) );
  fulladder U7265 ( .a(n7040), .b(n7039), .ci(n7038), .co(n7034), .s(n7041) );
  inv_1 U7266 ( .ip(n7041), .op(\STAGE_1/M4/sum [4]) );
  or2_1 U7267 ( .ip1(n7048), .ip2(n7042), .op(n7044) );
  nand2_1 U7268 ( .ip1(n7044), .ip2(n7043), .op(n7047) );
  nand2_1 U7269 ( .ip1(n7045), .ip2(column[61]), .op(n7046) );
  nand2_1 U7270 ( .ip1(n7045), .ip2(column[62]), .op(n7052) );
  inv_1 U7271 ( .ip(n7046), .op(n7051) );
  fulladder U7272 ( .a(n7048), .b(n7047), .ci(n7046), .co(n7050), .s(
        \STAGE_1/M4/sum [13]) );
  nor2_1 U7273 ( .ip1(column[62]), .ip2(column[63]), .op(n7049) );
  not_ab_or_c_or_d U7274 ( .ip1(column[62]), .ip2(column[63]), .ip3(n7049), 
        .ip4(n8180), .op(n7054) );
  fulladder U7275 ( .a(n7052), .b(n7051), .ci(n7050), .co(n7053), .s(
        \STAGE_1/M4/sum [14]) );
  xnor2_1 U7276 ( .ip1(n7054), .ip2(n7053), .op(\STAGE_1/M4/sum [15]) );
  nand2_1 U7277 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[71]), .op(n7161)
         );
  inv_1 U7278 ( .ip(n7055), .op(n7059) );
  nor2_1 U7279 ( .ip1(n7057), .ip2(n7056), .op(n7058) );
  nor2_1 U7280 ( .ip1(n7059), .ip2(n7058), .op(n7160) );
  fulladder U7281 ( .a(n7062), .b(n7061), .ci(n7060), .co(n7159), .s(n5932) );
  inv_1 U7282 ( .ip(n7063), .op(n7175) );
  nand2_1 U7283 ( .ip1(n8064), .ip2(m1Inputs[70]), .op(n7113) );
  nand2_1 U7284 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[70]), .op(n7115)
         );
  nor3_1 U7285 ( .ip1(n7813), .ip2(n7115), .ip3(n7122), .op(n7143) );
  or2_1 U7286 ( .ip1(n7113), .ip2(n7143), .op(n7066) );
  nand2_1 U7287 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[69]), .op(n7064)
         );
  or2_1 U7288 ( .ip1(n7064), .ip2(n7143), .op(n7065) );
  nand2_1 U7289 ( .ip1(n7066), .ip2(n7065), .op(n7141) );
  nand2_1 U7290 ( .ip1(n8009), .ip2(column[67]), .op(n7142) );
  xor2_1 U7291 ( .ip1(n7141), .ip2(n7142), .op(n7171) );
  fulladder U7292 ( .a(n7069), .b(n7068), .ci(n7067), .co(n7170), .s(n5938) );
  nand2_1 U7293 ( .ip1(\STAGE_1/weightReg [7]), .ip2(m1Inputs[68]), .op(n7149)
         );
  nor2_1 U7294 ( .ip1(n7070), .ip2(n8029), .op(n7148) );
  nand2_1 U7295 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[72]), .op(n7147)
         );
  inv_1 U7296 ( .ip(n7071), .op(n7174) );
  fulladder U7297 ( .a(n7074), .b(n7073), .ci(n7072), .co(n7173), .s(n5925) );
  inv_1 U7298 ( .ip(n7075), .op(n7187) );
  fulladder U7299 ( .a(n7078), .b(n7077), .ci(n7076), .co(n7079), .s(n7085) );
  inv_1 U7300 ( .ip(n7079), .op(n7186) );
  fulladder U7301 ( .a(n7082), .b(n7081), .ci(n7080), .co(n7185), .s(n5930) );
  inv_1 U7302 ( .ip(n7083), .op(n7183) );
  fulladder U7303 ( .a(n7086), .b(n7085), .ci(n7084), .co(n7182), .s(n7089) );
  fulladder U7304 ( .a(n7089), .b(n7088), .ci(n7087), .co(n7181), .s(
        \STAGE_1/M5/sum [2]) );
  inv_1 U7305 ( .ip(column[77]), .op(n7234) );
  nor2_1 U7306 ( .ip1(n8180), .ip2(n7234), .op(n7240) );
  nor2_1 U7307 ( .ip1(n7121), .ip2(n8029), .op(n7190) );
  nand2_1 U7308 ( .ip1(\STAGE_1/weightReg [7]), .ip2(m1Inputs[72]), .op(n7093)
         );
  nor2_1 U7309 ( .ip1(n7090), .ip2(n7628), .op(n7092) );
  nand2_1 U7310 ( .ip1(n8009), .ip2(column[71]), .op(n7091) );
  nand2_1 U7311 ( .ip1(n8009), .ip2(column[72]), .op(n7188) );
  fulladder U7312 ( .a(n7093), .b(n7092), .ci(n7091), .co(n7189), .s(n7109) );
  nand2_1 U7313 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[71]), .op(n7114)
         );
  nor2_1 U7314 ( .ip1(n7093), .ip2(n7114), .op(n7098) );
  or2_1 U7315 ( .ip1(n7094), .ip2(n7098), .op(n7096) );
  nand2_1 U7316 ( .ip1(n7882), .ip2(m1Inputs[71]), .op(n7102) );
  or2_1 U7317 ( .ip1(n7102), .ip2(n7098), .op(n7095) );
  nand2_1 U7318 ( .ip1(n7096), .ip2(n7095), .op(n7100) );
  and3_1 U7319 ( .ip1(n8051), .ip2(column[70]), .ip3(n7100), .op(n7097) );
  nor2_1 U7320 ( .ip1(n7098), .ip2(n7097), .op(n7108) );
  nand2_1 U7321 ( .ip1(n8009), .ip2(column[70]), .op(n7099) );
  xor2_1 U7322 ( .ip1(n7100), .ip2(n7099), .op(n7112) );
  nor2_1 U7323 ( .ip1(n7101), .ip2(n7628), .op(n7111) );
  nor2_1 U7324 ( .ip1(n7102), .ip2(n7115), .op(n7106) );
  or2_1 U7325 ( .ip1(n7114), .ip2(n7106), .op(n7105) );
  nand2_1 U7326 ( .ip1(\STAGE_1/weightReg [7]), .ip2(m1Inputs[70]), .op(n7103)
         );
  or2_1 U7327 ( .ip1(n7103), .ip2(n7106), .op(n7104) );
  nand2_1 U7328 ( .ip1(n7105), .ip2(n7104), .op(n7127) );
  and3_1 U7329 ( .ip1(n8051), .ip2(column[69]), .ip3(n7127), .op(n7129) );
  nor2_1 U7330 ( .ip1(n7106), .ip2(n7129), .op(n7110) );
  fulladder U7331 ( .a(n7109), .b(n7108), .ci(n7107), .co(n7215), .s(n7220) );
  fulladder U7332 ( .a(n7112), .b(n7111), .ci(n7110), .co(n7107), .s(n7136) );
  nand2_1 U7333 ( .ip1(n8064), .ip2(m1Inputs[72]), .op(n7125) );
  nor2_1 U7334 ( .ip1(n7122), .ip2(n8029), .op(n7124) );
  nor2_1 U7335 ( .ip1(n7114), .ip2(n7113), .op(n7120) );
  or2_1 U7336 ( .ip1(n7115), .ip2(n7120), .op(n7118) );
  or2_1 U7337 ( .ip1(n7116), .ip2(n7120), .op(n7117) );
  nand2_1 U7338 ( .ip1(n7118), .ip2(n7117), .op(n7151) );
  and3_1 U7339 ( .ip1(n8051), .ip2(column[68]), .ip3(n7151), .op(n7119) );
  nor2_1 U7340 ( .ip1(n7120), .ip2(n7119), .op(n7123) );
  nor2_1 U7341 ( .ip1(n5060), .ip2(n7121), .op(n7154) );
  nor2_1 U7342 ( .ip1(n7685), .ip2(n7122), .op(n7153) );
  nand2_1 U7343 ( .ip1(m1Inputs[68]), .ip2(\STAGE_1/weightReg [15]), .op(n7152) );
  fulladder U7344 ( .a(n7125), .b(n7124), .ci(n7123), .co(n7135), .s(n7126) );
  inv_1 U7345 ( .ip(n7126), .op(n7138) );
  inv_1 U7346 ( .ip(n7127), .op(n7128) );
  or2_1 U7347 ( .ip1(n7128), .ip2(n7129), .op(n7132) );
  nand2_1 U7348 ( .ip1(n8009), .ip2(column[69]), .op(n7130) );
  or2_1 U7349 ( .ip1(n7130), .ip2(n7129), .op(n7131) );
  nand2_1 U7350 ( .ip1(n7132), .ip2(n7131), .op(n7137) );
  inv_1 U7351 ( .ip(n7133), .op(n7134) );
  fulladder U7352 ( .a(n7136), .b(n7135), .ci(n7134), .co(n7219), .s(n7224) );
  fulladder U7353 ( .a(n7139), .b(n7138), .ci(n7137), .co(n7133), .s(n7140) );
  inv_1 U7354 ( .ip(n7140), .op(n7164) );
  or2_1 U7355 ( .ip1(n7141), .ip2(n7143), .op(n7146) );
  inv_1 U7356 ( .ip(n7142), .op(n7144) );
  or2_1 U7357 ( .ip1(n7144), .ip2(n7143), .op(n7145) );
  nand2_1 U7358 ( .ip1(n7146), .ip2(n7145), .op(n7158) );
  fulladder U7359 ( .a(n7149), .b(n7148), .ci(n7147), .co(n7157), .s(n7169) );
  nand2_1 U7360 ( .ip1(n8009), .ip2(column[68]), .op(n7150) );
  xor2_1 U7361 ( .ip1(n7151), .ip2(n7150), .op(n7156) );
  fulladder U7362 ( .a(n7154), .b(n7153), .ci(n7152), .co(n7139), .s(n7155) );
  inv_1 U7363 ( .ip(n7155), .op(n7167) );
  fulladder U7364 ( .a(n7158), .b(n7157), .ci(n7156), .co(n7163), .s(n7166) );
  fulladder U7365 ( .a(n7161), .b(n7160), .ci(n7159), .co(n7165), .s(n7063) );
  fulladder U7366 ( .a(n7164), .b(n7163), .ci(n7162), .co(n7223), .s(n7228) );
  fulladder U7367 ( .a(n7167), .b(n7166), .ci(n7165), .co(n7162), .s(n7168) );
  inv_1 U7368 ( .ip(n7168), .op(n7179) );
  fulladder U7369 ( .a(n7171), .b(n7170), .ci(n7169), .co(n7172), .s(n7071) );
  inv_1 U7370 ( .ip(n7172), .op(n7178) );
  fulladder U7371 ( .a(n7175), .b(n7174), .ci(n7173), .co(n7177), .s(n7075) );
  inv_1 U7372 ( .ip(n7176), .op(n7227) );
  fulladder U7373 ( .a(n7179), .b(n7178), .ci(n7177), .co(n7176), .s(n7180) );
  inv_1 U7374 ( .ip(n7180), .op(n7232) );
  fulladder U7375 ( .a(n7183), .b(n7182), .ci(n7181), .co(n7184), .s(
        \STAGE_1/M5/sum [3]) );
  inv_1 U7376 ( .ip(n7184), .op(n7231) );
  fulladder U7377 ( .a(n7187), .b(n7186), .ci(n7185), .co(n7230), .s(n7083) );
  fulladder U7378 ( .a(n7190), .b(n7189), .ci(n7188), .co(n7207), .s(n7216) );
  nand2_1 U7379 ( .ip1(n8009), .ip2(column[73]), .op(n7212) );
  nor3_1 U7380 ( .ip1(n7208), .ip2(n7207), .ip3(n7212), .op(n7202) );
  and2_1 U7381 ( .ip1(column[74]), .ip2(n7202), .op(n7198) );
  nand2_1 U7382 ( .ip1(column[75]), .ip2(n7198), .op(n7195) );
  inv_1 U7383 ( .ip(n7195), .op(n7191) );
  nand2_1 U7384 ( .ip1(column[76]), .ip2(n7191), .op(n7193) );
  and2_1 U7385 ( .ip1(n8175), .ip2(column[76]), .op(n7197) );
  and2_1 U7386 ( .ip1(n8051), .ip2(column[74]), .op(n7206) );
  nand3_1 U7387 ( .ip1(n7208), .ip2(n7207), .ip3(n7212), .op(n7203) );
  nor2_1 U7388 ( .ip1(n7206), .ip2(n7203), .op(n7199) );
  nand2_1 U7389 ( .ip1(n8009), .ip2(column[75]), .op(n7201) );
  nand2_1 U7390 ( .ip1(n7199), .ip2(n7201), .op(n7194) );
  nor2_1 U7391 ( .ip1(n7197), .ip2(n7194), .op(n7237) );
  inv_1 U7392 ( .ip(n7237), .op(n7192) );
  nand2_1 U7393 ( .ip1(n7193), .ip2(n7192), .op(n7235) );
  xor2_1 U7394 ( .ip1(n7240), .ip2(n7235), .op(\STAGE_1/M5/sum [13]) );
  nand2_1 U7395 ( .ip1(n7195), .ip2(n7194), .op(n7196) );
  xor2_1 U7396 ( .ip1(n7197), .ip2(n7196), .op(\STAGE_1/M5/sum [12]) );
  nor2_1 U7397 ( .ip1(n7199), .ip2(n7198), .op(n7200) );
  xor2_1 U7398 ( .ip1(n7201), .ip2(n7200), .op(\STAGE_1/M5/sum [11]) );
  inv_1 U7399 ( .ip(n7202), .op(n7204) );
  nand2_1 U7400 ( .ip1(n7204), .ip2(n7203), .op(n7205) );
  xor2_1 U7401 ( .ip1(n7206), .ip2(n7205), .op(\STAGE_1/M5/sum [10]) );
  inv_1 U7402 ( .ip(n7212), .op(n7213) );
  nand2_1 U7403 ( .ip1(n7208), .ip2(n7207), .op(n7210) );
  or2_1 U7404 ( .ip1(n7208), .ip2(n7207), .op(n7209) );
  nand2_1 U7405 ( .ip1(n7210), .ip2(n7209), .op(n7211) );
  mux2_1 U7406 ( .ip1(n7213), .ip2(n7212), .s(n7211), .op(\STAGE_1/M5/sum [9])
         );
  fulladder U7407 ( .a(n7216), .b(n7215), .ci(n7214), .co(n7208), .s(n7217) );
  inv_1 U7408 ( .ip(n7217), .op(\STAGE_1/M5/sum [8]) );
  fulladder U7409 ( .a(n7220), .b(n7219), .ci(n7218), .co(n7214), .s(n7221) );
  inv_1 U7410 ( .ip(n7221), .op(\STAGE_1/M5/sum [7]) );
  fulladder U7411 ( .a(n7224), .b(n7223), .ci(n7222), .co(n7218), .s(n7225) );
  inv_1 U7412 ( .ip(n7225), .op(\STAGE_1/M5/sum [6]) );
  fulladder U7413 ( .a(n7228), .b(n7227), .ci(n7226), .co(n7222), .s(n7229) );
  inv_1 U7414 ( .ip(n7229), .op(\STAGE_1/M5/sum [5]) );
  fulladder U7415 ( .a(n7232), .b(n7231), .ci(n7230), .co(n7226), .s(n7233) );
  inv_1 U7416 ( .ip(n7233), .op(\STAGE_1/M5/sum [4]) );
  nand2_1 U7417 ( .ip1(n8009), .ip2(column[78]), .op(n7241) );
  nor3_1 U7418 ( .ip1(n8180), .ip2(n7235), .ip3(n7234), .op(n7236) );
  nor2_1 U7419 ( .ip1(n7237), .ip2(n7236), .op(n7239) );
  nor2_1 U7420 ( .ip1(column[78]), .ip2(column[79]), .op(n7238) );
  not_ab_or_c_or_d U7421 ( .ip1(column[78]), .ip2(column[79]), .ip3(n7238), 
        .ip4(n8180), .op(n7243) );
  fulladder U7422 ( .a(n7241), .b(n7240), .ci(n7239), .co(n7242), .s(
        \STAGE_1/M5/sum [14]) );
  xnor2_1 U7423 ( .ip1(n7243), .ip2(n7242), .op(\STAGE_1/M5/sum [15]) );
  nand2_1 U7424 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[87]), .op(n7348)
         );
  inv_1 U7425 ( .ip(n7244), .op(n7248) );
  nor2_1 U7426 ( .ip1(n7246), .ip2(n7245), .op(n7247) );
  nor2_1 U7427 ( .ip1(n7248), .ip2(n7247), .op(n7347) );
  fulladder U7428 ( .a(n7251), .b(n7250), .ci(n7249), .co(n7346), .s(n7271) );
  inv_1 U7429 ( .ip(n7252), .op(n7362) );
  nand2_1 U7430 ( .ip1(\STAGE_1/weightReg [7]), .ip2(m1Inputs[84]), .op(n7337)
         );
  nor2_1 U7431 ( .ip1(n7253), .ip2(n7628), .op(n7336) );
  nand2_1 U7432 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[88]), .op(n7335)
         );
  fulladder U7433 ( .a(n7256), .b(n7255), .ci(n7254), .co(n7357), .s(n7270) );
  nand2_1 U7434 ( .ip1(n8064), .ip2(m1Inputs[86]), .op(n7307) );
  nand2_1 U7435 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[86]), .op(n7309)
         );
  nor2_1 U7436 ( .ip1(n7309), .ip2(n7257), .op(n7331) );
  or2_1 U7437 ( .ip1(n7307), .ip2(n7331), .op(n7260) );
  nand2_1 U7438 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[85]), .op(n7258)
         );
  or2_1 U7439 ( .ip1(n7258), .ip2(n7331), .op(n7259) );
  nand2_1 U7440 ( .ip1(n7260), .ip2(n7259), .op(n7329) );
  nand2_1 U7441 ( .ip1(n8009), .ip2(column[83]), .op(n7330) );
  xor2_1 U7442 ( .ip1(n7329), .ip2(n7330), .op(n7356) );
  inv_1 U7443 ( .ip(n7261), .op(n7361) );
  fulladder U7444 ( .a(n7264), .b(n7263), .ci(n7262), .co(n7360), .s(n6013) );
  inv_1 U7445 ( .ip(n7265), .op(n7374) );
  fulladder U7446 ( .a(n7268), .b(n7267), .ci(n7266), .co(n7373), .s(n6014) );
  fulladder U7447 ( .a(n7271), .b(n7270), .ci(n7269), .co(n7372), .s(n6000) );
  inv_1 U7448 ( .ip(n7272), .op(n7370) );
  fulladder U7449 ( .a(n7275), .b(n7274), .ci(n7273), .co(n7369), .s(n7278) );
  fulladder U7450 ( .a(n7278), .b(n7277), .ci(n7276), .co(n7368), .s(
        \STAGE_1/M6/sum [2]) );
  inv_1 U7451 ( .ip(column[93]), .op(n7419) );
  nor2_1 U7452 ( .ip1(n8180), .ip2(n7419), .op(n7425) );
  and2_1 U7453 ( .ip1(m1Inputs[88]), .ip2(\STAGE_1/weightReg [15]), .op(n7282)
         );
  nand2_1 U7454 ( .ip1(n7882), .ip2(m1Inputs[88]), .op(n7285) );
  nor2_1 U7455 ( .ip1(n7279), .ip2(n8029), .op(n7284) );
  nand2_1 U7456 ( .ip1(n8009), .ip2(column[87]), .op(n7283) );
  nand2_1 U7457 ( .ip1(n8009), .ip2(column[88]), .op(n7280) );
  fulladder U7458 ( .a(n7282), .b(n7281), .ci(n7280), .co(n7396), .s(n7401) );
  fulladder U7459 ( .a(n7285), .b(n7284), .ci(n7283), .co(n7281), .s(n7302) );
  nand2_1 U7460 ( .ip1(\STAGE_1/weightReg [6]), .ip2(m1Inputs[87]), .op(n7308)
         );
  nor2_1 U7461 ( .ip1(n7285), .ip2(n7308), .op(n7290) );
  nand2_1 U7462 ( .ip1(\STAGE_1/weightReg [7]), .ip2(m1Inputs[87]), .op(n7294)
         );
  or2_1 U7463 ( .ip1(n7294), .ip2(n7290), .op(n7288) );
  nand2_1 U7464 ( .ip1(n8037), .ip2(m1Inputs[88]), .op(n7286) );
  or2_1 U7465 ( .ip1(n7286), .ip2(n7290), .op(n7287) );
  nand2_1 U7466 ( .ip1(n7288), .ip2(n7287), .op(n7292) );
  and3_1 U7467 ( .ip1(n8051), .ip2(column[86]), .ip3(n7292), .op(n7289) );
  nor2_1 U7468 ( .ip1(n7290), .ip2(n7289), .op(n7301) );
  nand2_1 U7469 ( .ip1(n8009), .ip2(column[86]), .op(n7291) );
  xor2_1 U7470 ( .ip1(n7292), .ip2(n7291), .op(n7305) );
  nor2_1 U7471 ( .ip1(n7293), .ip2(n7628), .op(n7304) );
  nor2_1 U7472 ( .ip1(n7294), .ip2(n7309), .op(n7299) );
  or2_1 U7473 ( .ip1(n7308), .ip2(n7299), .op(n7297) );
  nand2_1 U7474 ( .ip1(\STAGE_1/weightReg [7]), .ip2(m1Inputs[86]), .op(n7295)
         );
  or2_1 U7475 ( .ip1(n7295), .ip2(n7299), .op(n7296) );
  nand2_1 U7476 ( .ip1(n7297), .ip2(n7296), .op(n7318) );
  and3_1 U7477 ( .ip1(n8051), .ip2(column[85]), .ip3(n7318), .op(n7298) );
  nor2_1 U7478 ( .ip1(n7299), .ip2(n7298), .op(n7303) );
  fulladder U7479 ( .a(n7302), .b(n7301), .ci(n7300), .co(n7400), .s(n7405) );
  fulladder U7480 ( .a(n7305), .b(n7304), .ci(n7303), .co(n7300), .s(n7325) );
  nand2_1 U7481 ( .ip1(n8064), .ip2(m1Inputs[88]), .op(n7321) );
  nor2_1 U7482 ( .ip1(n7306), .ip2(n8029), .op(n7320) );
  nor2_1 U7483 ( .ip1(n7308), .ip2(n7307), .op(n7313) );
  or2_1 U7484 ( .ip1(n7309), .ip2(n7313), .op(n7312) );
  nand2_1 U7485 ( .ip1(n8064), .ip2(m1Inputs[87]), .op(n7310) );
  or2_1 U7486 ( .ip1(n7310), .ip2(n7313), .op(n7311) );
  nand2_1 U7487 ( .ip1(n7312), .ip2(n7311), .op(n7339) );
  or2_1 U7488 ( .ip1(n7339), .ip2(n7313), .op(n7316) );
  nand2_1 U7489 ( .ip1(n8009), .ip2(column[84]), .op(n7338) );
  inv_1 U7490 ( .ip(n7338), .op(n7314) );
  or2_1 U7491 ( .ip1(n7314), .ip2(n7313), .op(n7315) );
  nand2_1 U7492 ( .ip1(n7316), .ip2(n7315), .op(n7319) );
  nand2_1 U7493 ( .ip1(n8009), .ip2(column[85]), .op(n7317) );
  xor2_1 U7494 ( .ip1(n7318), .ip2(n7317), .op(n7328) );
  fulladder U7495 ( .a(n7321), .b(n7320), .ci(n7319), .co(n7324), .s(n7327) );
  nor2_1 U7496 ( .ip1(n7322), .ip2(n8029), .op(n7342) );
  nand2_1 U7497 ( .ip1(\STAGE_1/weightReg [7]), .ip2(m1Inputs[85]), .op(n7341)
         );
  nand2_1 U7498 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[88]), .op(n7340)
         );
  fulladder U7499 ( .a(n7325), .b(n7324), .ci(n7323), .co(n7404), .s(n7409) );
  fulladder U7500 ( .a(n7328), .b(n7327), .ci(n7326), .co(n7323), .s(n7351) );
  or2_1 U7501 ( .ip1(n7329), .ip2(n7331), .op(n7334) );
  inv_1 U7502 ( .ip(n7330), .op(n7332) );
  or2_1 U7503 ( .ip1(n7332), .ip2(n7331), .op(n7333) );
  nand2_1 U7504 ( .ip1(n7334), .ip2(n7333), .op(n7345) );
  fulladder U7505 ( .a(n7337), .b(n7336), .ci(n7335), .co(n7344), .s(n7358) );
  xor2_1 U7506 ( .ip1(n7339), .ip2(n7338), .op(n7343) );
  fulladder U7507 ( .a(n7342), .b(n7341), .ci(n7340), .co(n7326), .s(n7354) );
  fulladder U7508 ( .a(n7345), .b(n7344), .ci(n7343), .co(n7350), .s(n7353) );
  fulladder U7509 ( .a(n7348), .b(n7347), .ci(n7346), .co(n7352), .s(n7252) );
  fulladder U7510 ( .a(n7351), .b(n7350), .ci(n7349), .co(n7408), .s(n7413) );
  fulladder U7511 ( .a(n7354), .b(n7353), .ci(n7352), .co(n7349), .s(n7355) );
  inv_1 U7512 ( .ip(n7355), .op(n7366) );
  fulladder U7513 ( .a(n7358), .b(n7357), .ci(n7356), .co(n7359), .s(n7261) );
  inv_1 U7514 ( .ip(n7359), .op(n7365) );
  fulladder U7515 ( .a(n7362), .b(n7361), .ci(n7360), .co(n7364), .s(n7265) );
  inv_1 U7516 ( .ip(n7363), .op(n7412) );
  fulladder U7517 ( .a(n7366), .b(n7365), .ci(n7364), .co(n7363), .s(n7367) );
  inv_1 U7518 ( .ip(n7367), .op(n7417) );
  fulladder U7519 ( .a(n7370), .b(n7369), .ci(n7368), .co(n7371), .s(
        \STAGE_1/M6/sum [3]) );
  inv_1 U7520 ( .ip(n7371), .op(n7416) );
  fulladder U7521 ( .a(n7374), .b(n7373), .ci(n7372), .co(n7415), .s(n7272) );
  nand2_1 U7522 ( .ip1(n8009), .ip2(column[89]), .op(n7397) );
  nor3_1 U7523 ( .ip1(n7396), .ip2(n7394), .ip3(n7397), .op(n7389) );
  nand3_1 U7524 ( .ip1(column[91]), .ip2(column[90]), .ip3(n7389), .op(n7377)
         );
  inv_1 U7525 ( .ip(n7377), .op(n7375) );
  nand2_1 U7526 ( .ip1(n7375), .ip2(column[92]), .op(n7379) );
  inv_1 U7527 ( .ip(n7396), .op(n7395) );
  nand2_1 U7528 ( .ip1(column[92]), .ip2(n8175), .op(n7381) );
  and2_1 U7529 ( .ip1(n8175), .ip2(column[90]), .op(n7393) );
  nand3_1 U7530 ( .ip1(n7396), .ip2(n7394), .ip3(n7397), .op(n7391) );
  nor2_1 U7531 ( .ip1(n7393), .ip2(n7391), .op(n7384) );
  nand2_1 U7532 ( .ip1(n8009), .ip2(column[91]), .op(n7387) );
  nand2_1 U7533 ( .ip1(n7384), .ip2(n7387), .op(n7376) );
  nand2_1 U7534 ( .ip1(n7377), .ip2(n7376), .op(n7380) );
  nand2_1 U7535 ( .ip1(n7381), .ip2(n7380), .op(n7383) );
  nor2_1 U7536 ( .ip1(n7395), .ip2(n7383), .op(n7422) );
  inv_1 U7537 ( .ip(n7422), .op(n7378) );
  nand2_1 U7538 ( .ip1(n7379), .ip2(n7378), .op(n7420) );
  xor2_1 U7539 ( .ip1(n7425), .ip2(n7420), .op(\STAGE_1/M6/sum [13]) );
  or2_1 U7540 ( .ip1(n7381), .ip2(n7380), .op(n7382) );
  nand2_1 U7541 ( .ip1(n7383), .ip2(n7382), .op(\STAGE_1/M6/sum [12]) );
  or2_1 U7542 ( .ip1(n7389), .ip2(n7384), .op(n7386) );
  or2_1 U7543 ( .ip1(column[90]), .ip2(n7384), .op(n7385) );
  nand2_1 U7544 ( .ip1(n7386), .ip2(n7385), .op(n7388) );
  xor2_1 U7545 ( .ip1(n7388), .ip2(n7387), .op(\STAGE_1/M6/sum [11]) );
  inv_1 U7546 ( .ip(n7389), .op(n7390) );
  nand2_1 U7547 ( .ip1(n7391), .ip2(n7390), .op(n7392) );
  xor2_1 U7548 ( .ip1(n7393), .ip2(n7392), .op(\STAGE_1/M6/sum [10]) );
  mux2_1 U7549 ( .ip1(n7396), .ip2(n7395), .s(n7394), .op(n7398) );
  xor2_1 U7550 ( .ip1(n7398), .ip2(n7397), .op(\STAGE_1/M6/sum [9]) );
  fulladder U7551 ( .a(n7401), .b(n7400), .ci(n7399), .co(n7394), .s(n7402) );
  inv_1 U7552 ( .ip(n7402), .op(\STAGE_1/M6/sum [8]) );
  fulladder U7553 ( .a(n7405), .b(n7404), .ci(n7403), .co(n7399), .s(n7406) );
  inv_1 U7554 ( .ip(n7406), .op(\STAGE_1/M6/sum [7]) );
  fulladder U7555 ( .a(n7409), .b(n7408), .ci(n7407), .co(n7403), .s(n7410) );
  inv_1 U7556 ( .ip(n7410), .op(\STAGE_1/M6/sum [6]) );
  fulladder U7557 ( .a(n7413), .b(n7412), .ci(n7411), .co(n7407), .s(n7414) );
  inv_1 U7558 ( .ip(n7414), .op(\STAGE_1/M6/sum [5]) );
  fulladder U7559 ( .a(n7417), .b(n7416), .ci(n7415), .co(n7411), .s(n7418) );
  inv_1 U7560 ( .ip(n7418), .op(\STAGE_1/M6/sum [4]) );
  nand2_1 U7561 ( .ip1(n8009), .ip2(column[94]), .op(n7426) );
  nor3_1 U7562 ( .ip1(n8180), .ip2(n7420), .ip3(n7419), .op(n7421) );
  nor2_1 U7563 ( .ip1(n7422), .ip2(n7421), .op(n7424) );
  nor2_1 U7564 ( .ip1(column[94]), .ip2(column[95]), .op(n7423) );
  not_ab_or_c_or_d U7565 ( .ip1(column[94]), .ip2(column[95]), .ip3(n7423), 
        .ip4(n8180), .op(n7428) );
  fulladder U7566 ( .a(n7426), .b(n7425), .ci(n7424), .co(n7427), .s(
        \STAGE_1/M6/sum [14]) );
  xnor2_1 U7567 ( .ip1(n7428), .ip2(n7427), .op(\STAGE_1/M6/sum [15]) );
  nand2_1 U7568 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[103]), .op(n7535) );
  inv_1 U7569 ( .ip(n7429), .op(n7433) );
  nor2_1 U7570 ( .ip1(n7431), .ip2(n7430), .op(n7432) );
  nor2_1 U7571 ( .ip1(n7433), .ip2(n7432), .op(n7534) );
  fulladder U7572 ( .a(n7436), .b(n7435), .ci(n7434), .co(n7533), .s(n6063) );
  inv_1 U7573 ( .ip(n7437), .op(n7549) );
  nand2_1 U7574 ( .ip1(n8064), .ip2(m1Inputs[102]), .op(n7487) );
  nand2_1 U7575 ( .ip1(n8037), .ip2(m1Inputs[102]), .op(n7489) );
  nor3_1 U7576 ( .ip1(n7813), .ip2(n7489), .ip3(n7496), .op(n7517) );
  or2_1 U7577 ( .ip1(n7487), .ip2(n7517), .op(n7440) );
  nand2_1 U7578 ( .ip1(n8037), .ip2(m1Inputs[101]), .op(n7438) );
  or2_1 U7579 ( .ip1(n7438), .ip2(n7517), .op(n7439) );
  nand2_1 U7580 ( .ip1(n7440), .ip2(n7439), .op(n7515) );
  nand2_1 U7581 ( .ip1(n8009), .ip2(column[99]), .op(n7516) );
  xor2_1 U7582 ( .ip1(n7515), .ip2(n7516), .op(n7545) );
  fulladder U7583 ( .a(n7443), .b(n7442), .ci(n7441), .co(n7544), .s(n6069) );
  nand2_1 U7584 ( .ip1(\STAGE_1/weightReg [7]), .ip2(m1Inputs[100]), .op(n7523) );
  nor2_1 U7585 ( .ip1(n7444), .ip2(n7628), .op(n7522) );
  nand2_1 U7586 ( .ip1(n8001), .ip2(m1Inputs[104]), .op(n7521) );
  inv_1 U7587 ( .ip(n7445), .op(n7548) );
  fulladder U7588 ( .a(n7448), .b(n7447), .ci(n7446), .co(n7547), .s(n6082) );
  inv_1 U7589 ( .ip(n7449), .op(n7561) );
  fulladder U7590 ( .a(n7452), .b(n7451), .ci(n7450), .co(n7453), .s(n7460) );
  inv_1 U7591 ( .ip(n7453), .op(n7560) );
  fulladder U7592 ( .a(n7456), .b(n7455), .ci(n7454), .co(n7559), .s(n6087) );
  inv_1 U7593 ( .ip(n7457), .op(n7557) );
  fulladder U7594 ( .a(n7460), .b(n7459), .ci(n7458), .co(n7556), .s(n7463) );
  fulladder U7595 ( .a(n7463), .b(n7462), .ci(n7461), .co(n7555), .s(
        \STAGE_1/M7/sum [2]) );
  and2_1 U7596 ( .ip1(n8051), .ip2(column[108]), .op(n7609) );
  nor2_1 U7597 ( .ip1(n7495), .ip2(n7628), .op(n7564) );
  nand2_1 U7598 ( .ip1(n7882), .ip2(m1Inputs[104]), .op(n7467) );
  nor2_1 U7599 ( .ip1(n7464), .ip2(n7628), .op(n7466) );
  nand2_1 U7600 ( .ip1(n8175), .ip2(column[103]), .op(n7465) );
  nand2_1 U7601 ( .ip1(n8175), .ip2(column[104]), .op(n7562) );
  fulladder U7602 ( .a(n7467), .b(n7466), .ci(n7465), .co(n7563), .s(n7483) );
  nand2_1 U7603 ( .ip1(n8037), .ip2(m1Inputs[103]), .op(n7488) );
  nor2_1 U7604 ( .ip1(n7467), .ip2(n7488), .op(n7472) );
  nand2_1 U7605 ( .ip1(n8037), .ip2(m1Inputs[104]), .op(n7468) );
  or2_1 U7606 ( .ip1(n7468), .ip2(n7472), .op(n7470) );
  nand2_1 U7607 ( .ip1(\STAGE_1/weightReg [7]), .ip2(m1Inputs[103]), .op(n7476) );
  or2_1 U7608 ( .ip1(n7476), .ip2(n7472), .op(n7469) );
  nand2_1 U7609 ( .ip1(n7470), .ip2(n7469), .op(n7474) );
  and3_1 U7610 ( .ip1(n8051), .ip2(column[102]), .ip3(n7474), .op(n7471) );
  nor2_1 U7611 ( .ip1(n7472), .ip2(n7471), .op(n7482) );
  nand2_1 U7612 ( .ip1(n8009), .ip2(column[102]), .op(n7473) );
  xor2_1 U7613 ( .ip1(n7474), .ip2(n7473), .op(n7486) );
  nor2_1 U7614 ( .ip1(n7475), .ip2(n7628), .op(n7485) );
  nor2_1 U7615 ( .ip1(n7476), .ip2(n7489), .op(n7480) );
  or2_1 U7616 ( .ip1(n7488), .ip2(n7480), .op(n7479) );
  nand2_1 U7617 ( .ip1(\STAGE_1/weightReg [7]), .ip2(m1Inputs[102]), .op(n7477) );
  or2_1 U7618 ( .ip1(n7477), .ip2(n7480), .op(n7478) );
  nand2_1 U7619 ( .ip1(n7479), .ip2(n7478), .op(n7501) );
  and3_1 U7620 ( .ip1(n8051), .ip2(column[101]), .ip3(n7501), .op(n7503) );
  nor2_1 U7621 ( .ip1(n7480), .ip2(n7503), .op(n7484) );
  fulladder U7622 ( .a(n7483), .b(n7482), .ci(n7481), .co(n7585), .s(n7590) );
  fulladder U7623 ( .a(n7486), .b(n7485), .ci(n7484), .co(n7481), .s(n7510) );
  nand2_1 U7624 ( .ip1(n8064), .ip2(m1Inputs[104]), .op(n7499) );
  nor2_1 U7625 ( .ip1(n7496), .ip2(n7628), .op(n7498) );
  nor2_1 U7626 ( .ip1(n7488), .ip2(n7487), .op(n7494) );
  or2_1 U7627 ( .ip1(n7489), .ip2(n7494), .op(n7492) );
  or2_1 U7628 ( .ip1(n7490), .ip2(n7494), .op(n7491) );
  nand2_1 U7629 ( .ip1(n7492), .ip2(n7491), .op(n7525) );
  and3_1 U7630 ( .ip1(n8051), .ip2(column[100]), .ip3(n7525), .op(n7493) );
  nor2_1 U7631 ( .ip1(n7494), .ip2(n7493), .op(n7497) );
  nor2_1 U7632 ( .ip1(n5060), .ip2(n7495), .op(n7528) );
  nor2_1 U7633 ( .ip1(n7685), .ip2(n7496), .op(n7527) );
  nand2_1 U7634 ( .ip1(m1Inputs[100]), .ip2(\STAGE_1/weightReg [15]), .op(
        n7526) );
  fulladder U7635 ( .a(n7499), .b(n7498), .ci(n7497), .co(n7509), .s(n7500) );
  inv_1 U7636 ( .ip(n7500), .op(n7512) );
  inv_1 U7637 ( .ip(n7501), .op(n7502) );
  or2_1 U7638 ( .ip1(n7502), .ip2(n7503), .op(n7506) );
  nand2_1 U7639 ( .ip1(n8009), .ip2(column[101]), .op(n7504) );
  or2_1 U7640 ( .ip1(n7504), .ip2(n7503), .op(n7505) );
  nand2_1 U7641 ( .ip1(n7506), .ip2(n7505), .op(n7511) );
  inv_1 U7642 ( .ip(n7507), .op(n7508) );
  fulladder U7643 ( .a(n7510), .b(n7509), .ci(n7508), .co(n7589), .s(n7594) );
  fulladder U7644 ( .a(n7513), .b(n7512), .ci(n7511), .co(n7507), .s(n7514) );
  inv_1 U7645 ( .ip(n7514), .op(n7538) );
  or2_1 U7646 ( .ip1(n7515), .ip2(n7517), .op(n7520) );
  inv_1 U7647 ( .ip(n7516), .op(n7518) );
  or2_1 U7648 ( .ip1(n7518), .ip2(n7517), .op(n7519) );
  nand2_1 U7649 ( .ip1(n7520), .ip2(n7519), .op(n7532) );
  fulladder U7650 ( .a(n7523), .b(n7522), .ci(n7521), .co(n7531), .s(n7543) );
  nand2_1 U7651 ( .ip1(n8009), .ip2(column[100]), .op(n7524) );
  xor2_1 U7652 ( .ip1(n7525), .ip2(n7524), .op(n7530) );
  fulladder U7653 ( .a(n7528), .b(n7527), .ci(n7526), .co(n7513), .s(n7529) );
  inv_1 U7654 ( .ip(n7529), .op(n7541) );
  fulladder U7655 ( .a(n7532), .b(n7531), .ci(n7530), .co(n7537), .s(n7540) );
  fulladder U7656 ( .a(n7535), .b(n7534), .ci(n7533), .co(n7539), .s(n7437) );
  fulladder U7657 ( .a(n7538), .b(n7537), .ci(n7536), .co(n7593), .s(n7598) );
  fulladder U7658 ( .a(n7541), .b(n7540), .ci(n7539), .co(n7536), .s(n7542) );
  inv_1 U7659 ( .ip(n7542), .op(n7553) );
  fulladder U7660 ( .a(n7545), .b(n7544), .ci(n7543), .co(n7546), .s(n7445) );
  inv_1 U7661 ( .ip(n7546), .op(n7552) );
  fulladder U7662 ( .a(n7549), .b(n7548), .ci(n7547), .co(n7551), .s(n7449) );
  inv_1 U7663 ( .ip(n7550), .op(n7597) );
  fulladder U7664 ( .a(n7553), .b(n7552), .ci(n7551), .co(n7550), .s(n7554) );
  inv_1 U7665 ( .ip(n7554), .op(n7602) );
  fulladder U7666 ( .a(n7557), .b(n7556), .ci(n7555), .co(n7558), .s(
        \STAGE_1/M7/sum [3]) );
  inv_1 U7667 ( .ip(n7558), .op(n7601) );
  fulladder U7668 ( .a(n7561), .b(n7560), .ci(n7559), .co(n7600), .s(n7457) );
  fulladder U7669 ( .a(n7564), .b(n7563), .ci(n7562), .co(n7577), .s(n7586) );
  nand2_1 U7670 ( .ip1(n8175), .ip2(column[105]), .op(n7582) );
  inv_1 U7671 ( .ip(column[106]), .op(n7565) );
  nor4_1 U7672 ( .ip1(n7578), .ip2(n7577), .ip3(n7582), .ip4(n7565), .op(n7568) );
  nand2_1 U7673 ( .ip1(column[107]), .ip2(n7568), .op(n7605) );
  and2_1 U7674 ( .ip1(n8051), .ip2(column[107]), .op(n7572) );
  nand2_1 U7675 ( .ip1(n8175), .ip2(column[106]), .op(n7576) );
  nand4_1 U7676 ( .ip1(n7578), .ip2(n7577), .ip3(n7576), .ip4(n7582), .op(
        n7569) );
  nor2_1 U7677 ( .ip1(n7572), .ip2(n7569), .op(n7604) );
  inv_1 U7678 ( .ip(n7604), .op(n7566) );
  nand2_1 U7679 ( .ip1(n7605), .ip2(n7566), .op(n7567) );
  xor2_1 U7680 ( .ip1(n7609), .ip2(n7567), .op(\STAGE_1/M7/sum [12]) );
  inv_1 U7681 ( .ip(n7568), .op(n7570) );
  nand2_1 U7682 ( .ip1(n7570), .ip2(n7569), .op(n7571) );
  xor2_1 U7683 ( .ip1(n7572), .ip2(n7571), .op(\STAGE_1/M7/sum [11]) );
  and3_1 U7684 ( .ip1(n7578), .ip2(n7577), .ip3(n7582), .op(n7574) );
  nor3_1 U7685 ( .ip1(n7578), .ip2(n7577), .ip3(n7582), .op(n7573) );
  nor2_1 U7686 ( .ip1(n7574), .ip2(n7573), .op(n7575) );
  xor2_1 U7687 ( .ip1(n7576), .ip2(n7575), .op(\STAGE_1/M7/sum [10]) );
  inv_1 U7688 ( .ip(n7582), .op(n7583) );
  nand2_1 U7689 ( .ip1(n7578), .ip2(n7577), .op(n7580) );
  or2_1 U7690 ( .ip1(n7578), .ip2(n7577), .op(n7579) );
  nand2_1 U7691 ( .ip1(n7580), .ip2(n7579), .op(n7581) );
  mux2_1 U7692 ( .ip1(n7583), .ip2(n7582), .s(n7581), .op(\STAGE_1/M7/sum [9])
         );
  fulladder U7693 ( .a(n7586), .b(n7585), .ci(n7584), .co(n7578), .s(n7587) );
  inv_1 U7694 ( .ip(n7587), .op(\STAGE_1/M7/sum [8]) );
  fulladder U7695 ( .a(n7590), .b(n7589), .ci(n7588), .co(n7584), .s(n7591) );
  inv_1 U7696 ( .ip(n7591), .op(\STAGE_1/M7/sum [7]) );
  fulladder U7697 ( .a(n7594), .b(n7593), .ci(n7592), .co(n7588), .s(n7595) );
  inv_1 U7698 ( .ip(n7595), .op(\STAGE_1/M7/sum [6]) );
  fulladder U7699 ( .a(n7598), .b(n7597), .ci(n7596), .co(n7592), .s(n7599) );
  inv_1 U7700 ( .ip(n7599), .op(\STAGE_1/M7/sum [5]) );
  fulladder U7701 ( .a(n7602), .b(n7601), .ci(n7600), .co(n7596), .s(n7603) );
  inv_1 U7702 ( .ip(n7603), .op(\STAGE_1/M7/sum [4]) );
  or2_1 U7703 ( .ip1(n7609), .ip2(n7604), .op(n7606) );
  nand2_1 U7704 ( .ip1(n7606), .ip2(n7605), .op(n7608) );
  nand2_1 U7705 ( .ip1(n8009), .ip2(column[109]), .op(n7607) );
  nand2_1 U7706 ( .ip1(n8009), .ip2(column[110]), .op(n7613) );
  inv_1 U7707 ( .ip(n7607), .op(n7612) );
  fulladder U7708 ( .a(n7609), .b(n7608), .ci(n7607), .co(n7611), .s(
        \STAGE_1/M7/sum [13]) );
  nor2_1 U7709 ( .ip1(column[110]), .ip2(column[111]), .op(n7610) );
  not_ab_or_c_or_d U7710 ( .ip1(column[110]), .ip2(column[111]), .ip3(n7610), 
        .ip4(n8180), .op(n7615) );
  fulladder U7711 ( .a(n7613), .b(n7612), .ci(n7611), .co(n7614), .s(
        \STAGE_1/M7/sum [14]) );
  xnor2_1 U7712 ( .ip1(n7615), .ip2(n7614), .op(\STAGE_1/M7/sum [15]) );
  nand2_1 U7713 ( .ip1(n8078), .ip2(m1Inputs[119]), .op(n7724) );
  nor2_1 U7714 ( .ip1(n7617), .ip2(n7616), .op(n7618) );
  nor2_1 U7715 ( .ip1(n7619), .ip2(n7618), .op(n7723) );
  fulladder U7716 ( .a(n7622), .b(n7621), .ci(n7620), .co(n7722), .s(n6151) );
  inv_1 U7717 ( .ip(n7623), .op(n7733) );
  nand2_1 U7718 ( .ip1(n8037), .ip2(m1Inputs[118]), .op(n7677) );
  nor3_1 U7719 ( .ip1(n7624), .ip2(n7677), .ip3(n7684), .op(n7706) );
  or2_1 U7720 ( .ip1(n7675), .ip2(n7706), .op(n7627) );
  nand2_1 U7721 ( .ip1(n8037), .ip2(m1Inputs[117]), .op(n7625) );
  or2_1 U7722 ( .ip1(n7625), .ip2(n7706), .op(n7626) );
  nand2_1 U7723 ( .ip1(n7627), .ip2(n7626), .op(n7704) );
  nand2_1 U7724 ( .ip1(n8009), .ip2(column[115]), .op(n7705) );
  xor2_1 U7725 ( .ip1(n7704), .ip2(n7705), .op(n7737) );
  nand2_1 U7726 ( .ip1(n7882), .ip2(m1Inputs[116]), .op(n7712) );
  nor2_1 U7727 ( .ip1(n7629), .ip2(n7628), .op(n7711) );
  nand2_1 U7728 ( .ip1(n8001), .ip2(m1Inputs[120]), .op(n7710) );
  fulladder U7729 ( .a(n7632), .b(n7631), .ci(n7630), .co(n7735), .s(n6157) );
  inv_1 U7730 ( .ip(n7633), .op(n7732) );
  fulladder U7731 ( .a(n7636), .b(n7635), .ci(n7634), .co(n7731), .s(n6144) );
  inv_1 U7732 ( .ip(n7637), .op(n7747) );
  fulladder U7733 ( .a(n7640), .b(n7639), .ci(n7638), .co(n7641), .s(n7647) );
  inv_1 U7734 ( .ip(n7641), .op(n7746) );
  fulladder U7735 ( .a(n7644), .b(n7643), .ci(n7642), .co(n7745), .s(n6149) );
  inv_1 U7736 ( .ip(n7645), .op(n7743) );
  fulladder U7737 ( .a(n7648), .b(n7647), .ci(n7646), .co(n7742), .s(n7651) );
  fulladder U7738 ( .a(n7651), .b(n7650), .ci(n7649), .co(n7741), .s(
        \STAGE_1/M8/sum [2]) );
  inv_1 U7739 ( .ip(column[125]), .op(n7794) );
  nor2_1 U7740 ( .ip1(n8180), .ip2(n7794), .op(n7800) );
  nor2_1 U7741 ( .ip1(n7683), .ip2(n8029), .op(n7750) );
  nand2_1 U7742 ( .ip1(n7882), .ip2(m1Inputs[120]), .op(n7655) );
  nor2_1 U7743 ( .ip1(n7652), .ip2(n8029), .op(n7654) );
  nand2_1 U7744 ( .ip1(n8175), .ip2(column[119]), .op(n7653) );
  nand2_1 U7745 ( .ip1(n8175), .ip2(column[120]), .op(n7748) );
  fulladder U7746 ( .a(n7655), .b(n7654), .ci(n7653), .co(n7749), .s(n7671) );
  nand2_1 U7747 ( .ip1(n8037), .ip2(m1Inputs[119]), .op(n7676) );
  nor2_1 U7748 ( .ip1(n7655), .ip2(n7676), .op(n7660) );
  nand2_1 U7749 ( .ip1(n8037), .ip2(m1Inputs[120]), .op(n7656) );
  or2_1 U7750 ( .ip1(n7656), .ip2(n7660), .op(n7658) );
  nand2_1 U7751 ( .ip1(n7882), .ip2(m1Inputs[119]), .op(n7664) );
  or2_1 U7752 ( .ip1(n7664), .ip2(n7660), .op(n7657) );
  nand2_1 U7753 ( .ip1(n7658), .ip2(n7657), .op(n7662) );
  and3_1 U7754 ( .ip1(n8051), .ip2(column[118]), .ip3(n7662), .op(n7659) );
  nor2_1 U7755 ( .ip1(n7660), .ip2(n7659), .op(n7670) );
  nand2_1 U7756 ( .ip1(n8175), .ip2(column[118]), .op(n7661) );
  xor2_1 U7757 ( .ip1(n7662), .ip2(n7661), .op(n7674) );
  nor2_1 U7758 ( .ip1(n7663), .ip2(n8029), .op(n7673) );
  nor2_1 U7759 ( .ip1(n7664), .ip2(n7677), .op(n7668) );
  or2_1 U7760 ( .ip1(n7676), .ip2(n7668), .op(n7667) );
  nand2_1 U7761 ( .ip1(n7882), .ip2(m1Inputs[118]), .op(n7665) );
  or2_1 U7762 ( .ip1(n7665), .ip2(n7668), .op(n7666) );
  nand2_1 U7763 ( .ip1(n7667), .ip2(n7666), .op(n7690) );
  and3_1 U7764 ( .ip1(n8051), .ip2(column[117]), .ip3(n7690), .op(n7692) );
  nor2_1 U7765 ( .ip1(n7668), .ip2(n7692), .op(n7672) );
  fulladder U7766 ( .a(n7671), .b(n7670), .ci(n7669), .co(n7775), .s(n7780) );
  fulladder U7767 ( .a(n7674), .b(n7673), .ci(n7672), .co(n7669), .s(n7699) );
  nand2_1 U7768 ( .ip1(\STAGE_1/weightReg [5]), .ip2(m1Inputs[120]), .op(n7688) );
  nor2_1 U7769 ( .ip1(n7684), .ip2(n8029), .op(n7687) );
  nor2_1 U7770 ( .ip1(n7676), .ip2(n7675), .op(n7682) );
  or2_1 U7771 ( .ip1(n7677), .ip2(n7682), .op(n7680) );
  or2_1 U7772 ( .ip1(n7678), .ip2(n7682), .op(n7679) );
  nand2_1 U7773 ( .ip1(n7680), .ip2(n7679), .op(n7714) );
  and3_1 U7774 ( .ip1(n8051), .ip2(column[116]), .ip3(n7714), .op(n7681) );
  nor2_1 U7775 ( .ip1(n7682), .ip2(n7681), .op(n7686) );
  nor2_1 U7776 ( .ip1(n5060), .ip2(n7683), .op(n7717) );
  nor2_1 U7777 ( .ip1(n7685), .ip2(n7684), .op(n7716) );
  nand2_1 U7778 ( .ip1(m1Inputs[116]), .ip2(\STAGE_1/weightReg [15]), .op(
        n7715) );
  fulladder U7779 ( .a(n7688), .b(n7687), .ci(n7686), .co(n7698), .s(n7689) );
  inv_1 U7780 ( .ip(n7689), .op(n7701) );
  inv_1 U7781 ( .ip(n7690), .op(n7691) );
  or2_1 U7782 ( .ip1(n7691), .ip2(n7692), .op(n7695) );
  nand2_1 U7783 ( .ip1(n8009), .ip2(column[117]), .op(n7693) );
  or2_1 U7784 ( .ip1(n7693), .ip2(n7692), .op(n7694) );
  nand2_1 U7785 ( .ip1(n7695), .ip2(n7694), .op(n7700) );
  inv_1 U7786 ( .ip(n7696), .op(n7697) );
  fulladder U7787 ( .a(n7699), .b(n7698), .ci(n7697), .co(n7779), .s(n7784) );
  fulladder U7788 ( .a(n7702), .b(n7701), .ci(n7700), .co(n7696), .s(n7703) );
  inv_1 U7789 ( .ip(n7703), .op(n7727) );
  or2_1 U7790 ( .ip1(n7704), .ip2(n7706), .op(n7709) );
  inv_1 U7791 ( .ip(n7705), .op(n7707) );
  or2_1 U7792 ( .ip1(n7707), .ip2(n7706), .op(n7708) );
  nand2_1 U7793 ( .ip1(n7709), .ip2(n7708), .op(n7721) );
  fulladder U7794 ( .a(n7712), .b(n7711), .ci(n7710), .co(n7720), .s(n7736) );
  nand2_1 U7795 ( .ip1(n8175), .ip2(column[116]), .op(n7713) );
  xor2_1 U7796 ( .ip1(n7714), .ip2(n7713), .op(n7719) );
  fulladder U7797 ( .a(n7717), .b(n7716), .ci(n7715), .co(n7702), .s(n7718) );
  inv_1 U7798 ( .ip(n7718), .op(n7730) );
  fulladder U7799 ( .a(n7721), .b(n7720), .ci(n7719), .co(n7726), .s(n7729) );
  fulladder U7800 ( .a(n7724), .b(n7723), .ci(n7722), .co(n7728), .s(n7623) );
  fulladder U7801 ( .a(n7727), .b(n7726), .ci(n7725), .co(n7783), .s(n7788) );
  fulladder U7802 ( .a(n7730), .b(n7729), .ci(n7728), .co(n7725), .s(n7740) );
  fulladder U7803 ( .a(n7733), .b(n7732), .ci(n7731), .co(n7734), .s(n7637) );
  inv_1 U7804 ( .ip(n7734), .op(n7739) );
  fulladder U7805 ( .a(n7737), .b(n7736), .ci(n7735), .co(n7738), .s(n7633) );
  fulladder U7806 ( .a(n7740), .b(n7739), .ci(n7738), .co(n7787), .s(n7792) );
  fulladder U7807 ( .a(n7743), .b(n7742), .ci(n7741), .co(n7744), .s(
        \STAGE_1/M8/sum [3]) );
  inv_1 U7808 ( .ip(n7744), .op(n7791) );
  fulladder U7809 ( .a(n7747), .b(n7746), .ci(n7745), .co(n7790), .s(n7645) );
  fulladder U7810 ( .a(n7750), .b(n7749), .ci(n7748), .co(n7767), .s(n7776) );
  nand2_1 U7811 ( .ip1(n8175), .ip2(column[121]), .op(n7772) );
  nor3_1 U7812 ( .ip1(n7768), .ip2(n7767), .ip3(n7772), .op(n7762) );
  and2_1 U7813 ( .ip1(column[122]), .ip2(n7762), .op(n7758) );
  nand2_1 U7814 ( .ip1(column[123]), .ip2(n7758), .op(n7755) );
  inv_1 U7815 ( .ip(n7755), .op(n7751) );
  nand2_1 U7816 ( .ip1(column[124]), .ip2(n7751), .op(n7753) );
  and2_1 U7817 ( .ip1(n8175), .ip2(column[124]), .op(n7757) );
  and2_1 U7818 ( .ip1(n8175), .ip2(column[122]), .op(n7766) );
  nand3_1 U7819 ( .ip1(n7768), .ip2(n7767), .ip3(n7772), .op(n7763) );
  nor2_1 U7820 ( .ip1(n7766), .ip2(n7763), .op(n7759) );
  nand2_1 U7821 ( .ip1(n8175), .ip2(column[123]), .op(n7761) );
  nand2_1 U7822 ( .ip1(n7759), .ip2(n7761), .op(n7754) );
  nor2_1 U7823 ( .ip1(n7757), .ip2(n7754), .op(n7797) );
  inv_1 U7824 ( .ip(n7797), .op(n7752) );
  nand2_1 U7825 ( .ip1(n7753), .ip2(n7752), .op(n7795) );
  xor2_1 U7826 ( .ip1(n7800), .ip2(n7795), .op(\STAGE_1/M8/sum [13]) );
  nand2_1 U7827 ( .ip1(n7755), .ip2(n7754), .op(n7756) );
  xor2_1 U7828 ( .ip1(n7757), .ip2(n7756), .op(\STAGE_1/M8/sum [12]) );
  nor2_1 U7829 ( .ip1(n7759), .ip2(n7758), .op(n7760) );
  xor2_1 U7830 ( .ip1(n7761), .ip2(n7760), .op(\STAGE_1/M8/sum [11]) );
  inv_1 U7831 ( .ip(n7762), .op(n7764) );
  nand2_1 U7832 ( .ip1(n7764), .ip2(n7763), .op(n7765) );
  xor2_1 U7833 ( .ip1(n7766), .ip2(n7765), .op(\STAGE_1/M8/sum [10]) );
  inv_1 U7834 ( .ip(n7772), .op(n7773) );
  nand2_1 U7835 ( .ip1(n7768), .ip2(n7767), .op(n7770) );
  or2_1 U7836 ( .ip1(n7768), .ip2(n7767), .op(n7769) );
  nand2_1 U7837 ( .ip1(n7770), .ip2(n7769), .op(n7771) );
  mux2_1 U7838 ( .ip1(n7773), .ip2(n7772), .s(n7771), .op(\STAGE_1/M8/sum [9])
         );
  fulladder U7839 ( .a(n7776), .b(n7775), .ci(n7774), .co(n7768), .s(n7777) );
  inv_1 U7840 ( .ip(n7777), .op(\STAGE_1/M8/sum [8]) );
  fulladder U7841 ( .a(n7780), .b(n7779), .ci(n7778), .co(n7774), .s(n7781) );
  inv_1 U7842 ( .ip(n7781), .op(\STAGE_1/M8/sum [7]) );
  fulladder U7843 ( .a(n7784), .b(n7783), .ci(n7782), .co(n7778), .s(n7785) );
  inv_1 U7844 ( .ip(n7785), .op(\STAGE_1/M8/sum [6]) );
  fulladder U7845 ( .a(n7788), .b(n7787), .ci(n7786), .co(n7782), .s(n7789) );
  inv_1 U7846 ( .ip(n7789), .op(\STAGE_1/M8/sum [5]) );
  fulladder U7847 ( .a(n7792), .b(n7791), .ci(n7790), .co(n7786), .s(n7793) );
  inv_1 U7848 ( .ip(n7793), .op(\STAGE_1/M8/sum [4]) );
  nand2_1 U7849 ( .ip1(n8175), .ip2(column[126]), .op(n7801) );
  nor3_1 U7850 ( .ip1(n8180), .ip2(n7795), .ip3(n7794), .op(n7796) );
  nor2_1 U7851 ( .ip1(n7797), .ip2(n7796), .op(n7799) );
  nor2_1 U7852 ( .ip1(column[126]), .ip2(column[127]), .op(n7798) );
  not_ab_or_c_or_d U7853 ( .ip1(column[126]), .ip2(column[127]), .ip3(n7798), 
        .ip4(n8180), .op(n7803) );
  fulladder U7854 ( .a(n7801), .b(n7800), .ci(n7799), .co(n7802), .s(
        \STAGE_1/M8/sum [14]) );
  xnor2_1 U7855 ( .ip1(n7803), .ip2(n7802), .op(\STAGE_1/M8/sum [15]) );
  nand2_1 U7856 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[135]), .op(n7908) );
  inv_1 U7857 ( .ip(n7804), .op(n7808) );
  nor2_1 U7858 ( .ip1(n7806), .ip2(n7805), .op(n7807) );
  nor2_1 U7859 ( .ip1(n7808), .ip2(n7807), .op(n7907) );
  fulladder U7860 ( .a(n7811), .b(n7810), .ci(n7809), .co(n7906), .s(n6222) );
  inv_1 U7861 ( .ip(n7812), .op(n7922) );
  nand2_1 U7862 ( .ip1(\STAGE_1/weightReg [5]), .ip2(m1Inputs[134]), .op(n7866) );
  nand2_1 U7863 ( .ip1(n8037), .ip2(m1Inputs[134]), .op(n7868) );
  nor3_1 U7864 ( .ip1(n7813), .ip2(n7868), .ip3(n7865), .op(n7891) );
  or2_1 U7865 ( .ip1(n7866), .ip2(n7891), .op(n7816) );
  nand2_1 U7866 ( .ip1(n8037), .ip2(m1Inputs[133]), .op(n7814) );
  or2_1 U7867 ( .ip1(n7814), .ip2(n7891), .op(n7815) );
  nand2_1 U7868 ( .ip1(n7816), .ip2(n7815), .op(n7889) );
  nand2_1 U7869 ( .ip1(n8175), .ip2(column[131]), .op(n7890) );
  xor2_1 U7870 ( .ip1(n7889), .ip2(n7890), .op(n7918) );
  fulladder U7871 ( .a(n7819), .b(n7818), .ci(n7817), .co(n7917), .s(n6228) );
  nand2_1 U7872 ( .ip1(n7882), .ip2(m1Inputs[132]), .op(n7897) );
  nor2_1 U7873 ( .ip1(n7820), .ip2(n8029), .op(n7896) );
  nand2_1 U7874 ( .ip1(n8001), .ip2(m1Inputs[136]), .op(n7895) );
  inv_1 U7875 ( .ip(n7821), .op(n7921) );
  fulladder U7876 ( .a(n7824), .b(n7823), .ci(n7822), .co(n7920), .s(n6215) );
  inv_1 U7877 ( .ip(n7825), .op(n7934) );
  fulladder U7878 ( .a(n7828), .b(n7827), .ci(n7826), .co(n7829), .s(n7835) );
  inv_1 U7879 ( .ip(n7829), .op(n7933) );
  fulladder U7880 ( .a(n7832), .b(n7831), .ci(n7830), .co(n7932), .s(n6220) );
  inv_1 U7881 ( .ip(n7833), .op(n7930) );
  fulladder U7882 ( .a(n7836), .b(n7835), .ci(n7834), .co(n7929), .s(n7839) );
  fulladder U7883 ( .a(n7839), .b(n7838), .ci(n7837), .co(n7928), .s(
        \STAGE_1/M9/sum [2]) );
  and2_1 U7884 ( .ip1(n8051), .ip2(column[141]), .op(n7987) );
  nor2_1 U7885 ( .ip1(n7840), .ip2(n8029), .op(n7937) );
  nand2_1 U7886 ( .ip1(n7882), .ip2(m1Inputs[136]), .op(n7858) );
  nor2_1 U7887 ( .ip1(n7841), .ip2(n8029), .op(n7857) );
  nand2_1 U7888 ( .ip1(n8175), .ip2(column[135]), .op(n7856) );
  nand2_1 U7889 ( .ip1(n8175), .ip2(column[136]), .op(n7935) );
  nand2_1 U7890 ( .ip1(n8037), .ip2(m1Inputs[135]), .op(n7867) );
  nor2_1 U7891 ( .ip1(n7858), .ip2(n7867), .op(n7846) );
  nand2_1 U7892 ( .ip1(n7882), .ip2(m1Inputs[135]), .op(n7850) );
  or2_1 U7893 ( .ip1(n7850), .ip2(n7846), .op(n7844) );
  nand2_1 U7894 ( .ip1(n8037), .ip2(m1Inputs[136]), .op(n7842) );
  or2_1 U7895 ( .ip1(n7842), .ip2(n7846), .op(n7843) );
  nand2_1 U7896 ( .ip1(n7844), .ip2(n7843), .op(n7848) );
  and3_1 U7897 ( .ip1(n8051), .ip2(column[134]), .ip3(n7848), .op(n7845) );
  nor2_1 U7898 ( .ip1(n7846), .ip2(n7845), .op(n7861) );
  nand2_1 U7899 ( .ip1(n8175), .ip2(column[134]), .op(n7847) );
  xor2_1 U7900 ( .ip1(n7848), .ip2(n7847), .op(n7864) );
  nor2_1 U7901 ( .ip1(n7849), .ip2(n8029), .op(n7863) );
  nor2_1 U7902 ( .ip1(n7850), .ip2(n7868), .op(n7855) );
  or2_1 U7903 ( .ip1(n7867), .ip2(n7855), .op(n7853) );
  nand2_1 U7904 ( .ip1(n7882), .ip2(m1Inputs[134]), .op(n7851) );
  or2_1 U7905 ( .ip1(n7851), .ip2(n7855), .op(n7852) );
  nand2_1 U7906 ( .ip1(n7853), .ip2(n7852), .op(n7877) );
  and3_1 U7907 ( .ip1(n8051), .ip2(column[133]), .ip3(n7877), .op(n7854) );
  nor2_1 U7908 ( .ip1(n7855), .ip2(n7854), .op(n7862) );
  fulladder U7909 ( .a(n7858), .b(n7857), .ci(n7856), .co(n7936), .s(n7859) );
  fulladder U7910 ( .a(n7861), .b(n7860), .ci(n7859), .co(n7963), .s(n7968) );
  fulladder U7911 ( .a(n7864), .b(n7863), .ci(n7862), .co(n7860), .s(n7885) );
  nand2_1 U7912 ( .ip1(\STAGE_1/weightReg [5]), .ip2(m1Inputs[136]), .op(n7880) );
  nor2_1 U7913 ( .ip1(n7865), .ip2(n8029), .op(n7879) );
  nor2_1 U7914 ( .ip1(n7867), .ip2(n7866), .op(n7872) );
  or2_1 U7915 ( .ip1(n7868), .ip2(n7872), .op(n7871) );
  nand2_1 U7916 ( .ip1(n8064), .ip2(m1Inputs[135]), .op(n7869) );
  or2_1 U7917 ( .ip1(n7869), .ip2(n7872), .op(n7870) );
  nand2_1 U7918 ( .ip1(n7871), .ip2(n7870), .op(n7899) );
  or2_1 U7919 ( .ip1(n7899), .ip2(n7872), .op(n7875) );
  nand2_1 U7920 ( .ip1(n8175), .ip2(column[132]), .op(n7898) );
  inv_1 U7921 ( .ip(n7898), .op(n7873) );
  or2_1 U7922 ( .ip1(n7873), .ip2(n7872), .op(n7874) );
  nand2_1 U7923 ( .ip1(n7875), .ip2(n7874), .op(n7878) );
  nand2_1 U7924 ( .ip1(n8175), .ip2(column[133]), .op(n7876) );
  xor2_1 U7925 ( .ip1(n7877), .ip2(n7876), .op(n7888) );
  fulladder U7926 ( .a(n7880), .b(n7879), .ci(n7878), .co(n7884), .s(n7887) );
  nor2_1 U7927 ( .ip1(n7881), .ip2(n8029), .op(n7902) );
  nand2_1 U7928 ( .ip1(n7882), .ip2(m1Inputs[133]), .op(n7901) );
  nand2_1 U7929 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[136]), .op(n7900) );
  fulladder U7930 ( .a(n7885), .b(n7884), .ci(n7883), .co(n7967), .s(n7972) );
  fulladder U7931 ( .a(n7888), .b(n7887), .ci(n7886), .co(n7883), .s(n7911) );
  or2_1 U7932 ( .ip1(n7889), .ip2(n7891), .op(n7894) );
  inv_1 U7933 ( .ip(n7890), .op(n7892) );
  or2_1 U7934 ( .ip1(n7892), .ip2(n7891), .op(n7893) );
  nand2_1 U7935 ( .ip1(n7894), .ip2(n7893), .op(n7905) );
  fulladder U7936 ( .a(n7897), .b(n7896), .ci(n7895), .co(n7904), .s(n7916) );
  xor2_1 U7937 ( .ip1(n7899), .ip2(n7898), .op(n7903) );
  fulladder U7938 ( .a(n7902), .b(n7901), .ci(n7900), .co(n7886), .s(n7914) );
  fulladder U7939 ( .a(n7905), .b(n7904), .ci(n7903), .co(n7910), .s(n7913) );
  fulladder U7940 ( .a(n7908), .b(n7907), .ci(n7906), .co(n7912), .s(n7812) );
  fulladder U7941 ( .a(n7911), .b(n7910), .ci(n7909), .co(n7971), .s(n7976) );
  fulladder U7942 ( .a(n7914), .b(n7913), .ci(n7912), .co(n7909), .s(n7915) );
  inv_1 U7943 ( .ip(n7915), .op(n7926) );
  fulladder U7944 ( .a(n7918), .b(n7917), .ci(n7916), .co(n7919), .s(n7821) );
  inv_1 U7945 ( .ip(n7919), .op(n7925) );
  fulladder U7946 ( .a(n7922), .b(n7921), .ci(n7920), .co(n7924), .s(n7825) );
  inv_1 U7947 ( .ip(n7923), .op(n7975) );
  fulladder U7948 ( .a(n7926), .b(n7925), .ci(n7924), .co(n7923), .s(n7927) );
  inv_1 U7949 ( .ip(n7927), .op(n7980) );
  fulladder U7950 ( .a(n7930), .b(n7929), .ci(n7928), .co(n7931), .s(
        \STAGE_1/M9/sum [3]) );
  inv_1 U7951 ( .ip(n7931), .op(n7979) );
  fulladder U7952 ( .a(n7934), .b(n7933), .ci(n7932), .co(n7978), .s(n7833) );
  fulladder U7953 ( .a(n7937), .b(n7936), .ci(n7935), .co(n7955), .s(n7964) );
  nand2_1 U7954 ( .ip1(n8175), .ip2(column[137]), .op(n7960) );
  nor3_1 U7955 ( .ip1(n7956), .ip2(n7955), .ip3(n7960), .op(n7951) );
  nand2_1 U7956 ( .ip1(n8175), .ip2(column[139]), .op(n7950) );
  inv_1 U7957 ( .ip(n7950), .op(n7949) );
  nand3_1 U7958 ( .ip1(column[138]), .ip2(n7951), .ip3(n7949), .op(n7942) );
  inv_1 U7959 ( .ip(n7942), .op(n7938) );
  nand2_1 U7960 ( .ip1(column[140]), .ip2(n7938), .op(n7983) );
  and2_1 U7961 ( .ip1(n8051), .ip2(column[140]), .op(n7944) );
  nand2_1 U7962 ( .ip1(n8175), .ip2(column[138]), .op(n7954) );
  and4_1 U7963 ( .ip1(n7956), .ip2(n7955), .ip3(n7954), .ip4(n7960), .op(n7945) );
  nand2_1 U7964 ( .ip1(n7945), .ip2(n7950), .op(n7941) );
  nor2_1 U7965 ( .ip1(n7944), .ip2(n7941), .op(n7982) );
  inv_1 U7966 ( .ip(n7982), .op(n7939) );
  nand2_1 U7967 ( .ip1(n7983), .ip2(n7939), .op(n7940) );
  xor2_1 U7968 ( .ip1(n7987), .ip2(n7940), .op(\STAGE_1/M9/sum [13]) );
  nand2_1 U7969 ( .ip1(n7942), .ip2(n7941), .op(n7943) );
  xor2_1 U7970 ( .ip1(n7944), .ip2(n7943), .op(\STAGE_1/M9/sum [12]) );
  or2_1 U7971 ( .ip1(column[138]), .ip2(n7945), .op(n7947) );
  or2_1 U7972 ( .ip1(n7951), .ip2(n7945), .op(n7946) );
  nand2_1 U7973 ( .ip1(n7947), .ip2(n7946), .op(n7948) );
  mux2_1 U7974 ( .ip1(n7950), .ip2(n7949), .s(n7948), .op(\STAGE_1/M9/sum [11]) );
  and3_1 U7975 ( .ip1(n7956), .ip2(n7955), .ip3(n7960), .op(n7952) );
  nor2_1 U7976 ( .ip1(n7952), .ip2(n7951), .op(n7953) );
  xor2_1 U7977 ( .ip1(n7954), .ip2(n7953), .op(\STAGE_1/M9/sum [10]) );
  inv_1 U7978 ( .ip(n7960), .op(n7961) );
  nand2_1 U7979 ( .ip1(n7956), .ip2(n7955), .op(n7958) );
  or2_1 U7980 ( .ip1(n7956), .ip2(n7955), .op(n7957) );
  nand2_1 U7981 ( .ip1(n7958), .ip2(n7957), .op(n7959) );
  mux2_1 U7982 ( .ip1(n7961), .ip2(n7960), .s(n7959), .op(\STAGE_1/M9/sum [9])
         );
  fulladder U7983 ( .a(n7964), .b(n7963), .ci(n7962), .co(n7956), .s(n7965) );
  inv_1 U7984 ( .ip(n7965), .op(\STAGE_1/M9/sum [8]) );
  fulladder U7985 ( .a(n7968), .b(n7967), .ci(n7966), .co(n7962), .s(n7969) );
  inv_1 U7986 ( .ip(n7969), .op(\STAGE_1/M9/sum [7]) );
  fulladder U7987 ( .a(n7972), .b(n7971), .ci(n7970), .co(n7966), .s(n7973) );
  inv_1 U7988 ( .ip(n7973), .op(\STAGE_1/M9/sum [6]) );
  fulladder U7989 ( .a(n7976), .b(n7975), .ci(n7974), .co(n7970), .s(n7977) );
  inv_1 U7990 ( .ip(n7977), .op(\STAGE_1/M9/sum [5]) );
  fulladder U7991 ( .a(n7980), .b(n7979), .ci(n7978), .co(n7974), .s(n7981) );
  inv_1 U7992 ( .ip(n7981), .op(\STAGE_1/M9/sum [4]) );
  nand2_1 U7993 ( .ip1(n8175), .ip2(column[142]), .op(n7988) );
  or2_1 U7994 ( .ip1(n7987), .ip2(n7982), .op(n7984) );
  nand2_1 U7995 ( .ip1(n7984), .ip2(n7983), .op(n7986) );
  nor2_1 U7996 ( .ip1(column[142]), .ip2(column[143]), .op(n7985) );
  not_ab_or_c_or_d U7997 ( .ip1(column[142]), .ip2(column[143]), .ip3(n7985), 
        .ip4(n8180), .op(n7990) );
  fulladder U7998 ( .a(n7988), .b(n7987), .ci(n7986), .co(n7989), .s(
        \STAGE_1/M9/sum [14]) );
  xnor2_1 U7999 ( .ip1(n7990), .ip2(n7989), .op(\STAGE_1/M9/sum [15]) );
  nand2_1 U8000 ( .ip1(n8078), .ip2(m1Inputs[151]), .op(n8104) );
  inv_1 U8001 ( .ip(n7991), .op(n7995) );
  nor2_1 U8002 ( .ip1(n7993), .ip2(n7992), .op(n7994) );
  nor2_1 U8003 ( .ip1(n7995), .ip2(n7994), .op(n8103) );
  fulladder U8004 ( .a(n7998), .b(n7997), .ci(n7996), .co(n8102), .s(n6281) );
  inv_1 U8005 ( .ip(n7999), .op(n8118) );
  nand2_1 U8006 ( .ip1(n7882), .ip2(m1Inputs[148]), .op(n8093) );
  nor2_1 U8007 ( .ip1(n8000), .ip2(n8029), .op(n8092) );
  nand2_1 U8008 ( .ip1(n8001), .ip2(m1Inputs[152]), .op(n8091) );
  fulladder U8009 ( .a(n8004), .b(n8003), .ci(n8002), .co(n8113), .s(n6287) );
  nand2_1 U8010 ( .ip1(\STAGE_1/weightReg [5]), .ip2(m1Inputs[150]), .op(n8061) );
  nand2_1 U8011 ( .ip1(n8037), .ip2(m1Inputs[150]), .op(n8063) );
  nor2_1 U8012 ( .ip1(n8063), .ip2(n8005), .op(n8087) );
  or2_1 U8013 ( .ip1(n8061), .ip2(n8087), .op(n8008) );
  nand2_1 U8014 ( .ip1(n8037), .ip2(m1Inputs[149]), .op(n8006) );
  or2_1 U8015 ( .ip1(n8006), .ip2(n8087), .op(n8007) );
  nand2_1 U8016 ( .ip1(n8008), .ip2(n8007), .op(n8085) );
  nand2_1 U8017 ( .ip1(n8009), .ip2(column[147]), .op(n8086) );
  xor2_1 U8018 ( .ip1(n8085), .ip2(n8086), .op(n8112) );
  inv_1 U8019 ( .ip(n8010), .op(n8117) );
  fulladder U8020 ( .a(n8013), .b(n8012), .ci(n8011), .co(n8116), .s(n6300) );
  inv_1 U8021 ( .ip(n8014), .op(n8130) );
  fulladder U8022 ( .a(n8017), .b(n8016), .ci(n8015), .co(n8018), .s(n8025) );
  inv_1 U8023 ( .ip(n8018), .op(n8129) );
  fulladder U8024 ( .a(n8021), .b(n8020), .ci(n8019), .co(n8128), .s(n6305) );
  inv_1 U8025 ( .ip(n8022), .op(n8126) );
  fulladder U8026 ( .a(n8025), .b(n8024), .ci(n8023), .co(n8125), .s(n8028) );
  fulladder U8027 ( .a(n8028), .b(n8027), .ci(n8026), .co(n8124), .s(
        \STAGE_1/M10/sum [2]) );
  inv_1 U8028 ( .ip(column[157]), .op(n8176) );
  nor2_1 U8029 ( .ip1(n8180), .ip2(n8176), .op(n8183) );
  and2_1 U8030 ( .ip1(n8051), .ip2(column[156]), .op(n8137) );
  nand2_1 U8031 ( .ip1(n8175), .ip2(column[155]), .op(n8142) );
  and2_1 U8032 ( .ip1(n8051), .ip2(column[154]), .op(n8147) );
  nor2_1 U8033 ( .ip1(n8030), .ip2(n8029), .op(n8034) );
  nand2_1 U8034 ( .ip1(\STAGE_1/weightReg [7]), .ip2(m1Inputs[152]), .op(n8038) );
  nor2_1 U8035 ( .ip1(n8031), .ip2(n8029), .op(n8036) );
  nand2_1 U8036 ( .ip1(n8175), .ip2(column[151]), .op(n8035) );
  nand2_1 U8037 ( .ip1(n8175), .ip2(column[152]), .op(n8032) );
  fulladder U8038 ( .a(n8034), .b(n8033), .ci(n8032), .co(n8149), .s(n8157) );
  fulladder U8039 ( .a(n8038), .b(n8036), .ci(n8035), .co(n8033), .s(n8056) );
  nand2_1 U8040 ( .ip1(n8037), .ip2(m1Inputs[151]), .op(n8062) );
  nor2_1 U8041 ( .ip1(n8038), .ip2(n8062), .op(n8043) );
  nand2_1 U8042 ( .ip1(\STAGE_1/weightReg [7]), .ip2(m1Inputs[151]), .op(n8047) );
  or2_1 U8043 ( .ip1(n8047), .ip2(n8043), .op(n8041) );
  or2_1 U8044 ( .ip1(n8039), .ip2(n8043), .op(n8040) );
  nand2_1 U8045 ( .ip1(n8041), .ip2(n8040), .op(n8045) );
  and3_1 U8046 ( .ip1(n8051), .ip2(column[150]), .ip3(n8045), .op(n8042) );
  nor2_1 U8047 ( .ip1(n8043), .ip2(n8042), .op(n8055) );
  nand2_1 U8048 ( .ip1(n8175), .ip2(column[150]), .op(n8044) );
  xor2_1 U8049 ( .ip1(n8045), .ip2(n8044), .op(n8059) );
  nor2_1 U8050 ( .ip1(n8046), .ip2(n8029), .op(n8058) );
  nor2_1 U8051 ( .ip1(n8047), .ip2(n8063), .op(n8053) );
  or2_1 U8052 ( .ip1(n8062), .ip2(n8053), .op(n8050) );
  nand2_1 U8053 ( .ip1(\STAGE_1/weightReg [7]), .ip2(m1Inputs[150]), .op(n8048) );
  or2_1 U8054 ( .ip1(n8048), .ip2(n8053), .op(n8049) );
  nand2_1 U8055 ( .ip1(n8050), .ip2(n8049), .op(n8073) );
  and3_1 U8056 ( .ip1(n8051), .ip2(column[149]), .ip3(n8073), .op(n8052) );
  nor2_1 U8057 ( .ip1(n8053), .ip2(n8052), .op(n8057) );
  fulladder U8058 ( .a(n8056), .b(n8055), .ci(n8054), .co(n8156), .s(n8161) );
  fulladder U8059 ( .a(n8059), .b(n8058), .ci(n8057), .co(n8054), .s(n8081) );
  nand2_1 U8060 ( .ip1(\STAGE_1/weightReg [5]), .ip2(m1Inputs[152]), .op(n8076) );
  nor2_1 U8061 ( .ip1(n8060), .ip2(n8029), .op(n8075) );
  nor2_1 U8062 ( .ip1(n8062), .ip2(n8061), .op(n8068) );
  or2_1 U8063 ( .ip1(n8063), .ip2(n8068), .op(n8067) );
  nand2_1 U8064 ( .ip1(n8064), .ip2(m1Inputs[151]), .op(n8065) );
  or2_1 U8065 ( .ip1(n8065), .ip2(n8068), .op(n8066) );
  nand2_1 U8066 ( .ip1(n8067), .ip2(n8066), .op(n8095) );
  or2_1 U8067 ( .ip1(n8095), .ip2(n8068), .op(n8071) );
  nand2_1 U8068 ( .ip1(n8175), .ip2(column[148]), .op(n8094) );
  inv_1 U8069 ( .ip(n8094), .op(n8069) );
  or2_1 U8070 ( .ip1(n8069), .ip2(n8068), .op(n8070) );
  nand2_1 U8071 ( .ip1(n8071), .ip2(n8070), .op(n8074) );
  nand2_1 U8072 ( .ip1(n8175), .ip2(column[149]), .op(n8072) );
  xor2_1 U8073 ( .ip1(n8073), .ip2(n8072), .op(n8084) );
  fulladder U8074 ( .a(n8076), .b(n8075), .ci(n8074), .co(n8080), .s(n8083) );
  nor2_1 U8075 ( .ip1(n8077), .ip2(n8029), .op(n8098) );
  nand2_1 U8076 ( .ip1(\STAGE_1/weightReg [7]), .ip2(m1Inputs[149]), .op(n8097) );
  nand2_1 U8077 ( .ip1(n8078), .ip2(m1Inputs[152]), .op(n8096) );
  fulladder U8078 ( .a(n8081), .b(n8080), .ci(n8079), .co(n8160), .s(n8165) );
  fulladder U8079 ( .a(n8084), .b(n8083), .ci(n8082), .co(n8079), .s(n8107) );
  or2_1 U8080 ( .ip1(n8085), .ip2(n8087), .op(n8090) );
  inv_1 U8081 ( .ip(n8086), .op(n8088) );
  or2_1 U8082 ( .ip1(n8088), .ip2(n8087), .op(n8089) );
  nand2_1 U8083 ( .ip1(n8090), .ip2(n8089), .op(n8101) );
  fulladder U8084 ( .a(n8093), .b(n8092), .ci(n8091), .co(n8100), .s(n8114) );
  xor2_1 U8085 ( .ip1(n8095), .ip2(n8094), .op(n8099) );
  fulladder U8086 ( .a(n8098), .b(n8097), .ci(n8096), .co(n8082), .s(n8110) );
  fulladder U8087 ( .a(n8101), .b(n8100), .ci(n8099), .co(n8106), .s(n8109) );
  fulladder U8088 ( .a(n8104), .b(n8103), .ci(n8102), .co(n8108), .s(n7999) );
  fulladder U8089 ( .a(n8107), .b(n8106), .ci(n8105), .co(n8164), .s(n8169) );
  fulladder U8090 ( .a(n8110), .b(n8109), .ci(n8108), .co(n8105), .s(n8111) );
  inv_1 U8091 ( .ip(n8111), .op(n8122) );
  fulladder U8092 ( .a(n8114), .b(n8113), .ci(n8112), .co(n8115), .s(n8010) );
  inv_1 U8093 ( .ip(n8115), .op(n8121) );
  fulladder U8094 ( .a(n8118), .b(n8117), .ci(n8116), .co(n8120), .s(n8014) );
  inv_1 U8095 ( .ip(n8119), .op(n8168) );
  fulladder U8096 ( .a(n8122), .b(n8121), .ci(n8120), .co(n8119), .s(n8123) );
  inv_1 U8097 ( .ip(n8123), .op(n8173) );
  fulladder U8098 ( .a(n8126), .b(n8125), .ci(n8124), .co(n8127), .s(
        \STAGE_1/M10/sum [3]) );
  inv_1 U8099 ( .ip(n8127), .op(n8172) );
  fulladder U8100 ( .a(n8130), .b(n8129), .ci(n8128), .co(n8171), .s(n8022) );
  nand2_1 U8101 ( .ip1(n8175), .ip2(column[153]), .op(n8153) );
  nand3_1 U8102 ( .ip1(n8149), .ip2(n8148), .ip3(n8153), .op(n8145) );
  nor2_1 U8103 ( .ip1(n8147), .ip2(n8145), .op(n8139) );
  nand2_1 U8104 ( .ip1(n8142), .ip2(n8139), .op(n8134) );
  nor2_1 U8105 ( .ip1(n8137), .ip2(n8134), .op(n8179) );
  inv_1 U8106 ( .ip(n8179), .op(n8132) );
  nor3_1 U8107 ( .ip1(n8149), .ip2(n8148), .ip3(n8153), .op(n8143) );
  nand2_1 U8108 ( .ip1(column[154]), .ip2(n8143), .op(n8138) );
  nor2_1 U8109 ( .ip1(n8142), .ip2(n8138), .op(n8133) );
  nand2_1 U8110 ( .ip1(column[156]), .ip2(n8133), .op(n8131) );
  nand2_1 U8111 ( .ip1(n8132), .ip2(n8131), .op(n8177) );
  xor2_1 U8112 ( .ip1(n8183), .ip2(n8177), .op(\STAGE_1/M10/sum [13]) );
  inv_1 U8113 ( .ip(n8133), .op(n8135) );
  nand2_1 U8114 ( .ip1(n8135), .ip2(n8134), .op(n8136) );
  xor2_1 U8115 ( .ip1(n8137), .ip2(n8136), .op(\STAGE_1/M10/sum [12]) );
  inv_1 U8116 ( .ip(n8138), .op(n8140) );
  nor2_1 U8117 ( .ip1(n8140), .ip2(n8139), .op(n8141) );
  xor2_1 U8118 ( .ip1(n8142), .ip2(n8141), .op(\STAGE_1/M10/sum [11]) );
  inv_1 U8119 ( .ip(n8143), .op(n8144) );
  nand2_1 U8120 ( .ip1(n8145), .ip2(n8144), .op(n8146) );
  xor2_1 U8121 ( .ip1(n8147), .ip2(n8146), .op(\STAGE_1/M10/sum [10]) );
  inv_1 U8122 ( .ip(n8153), .op(n8154) );
  or2_1 U8123 ( .ip1(n8149), .ip2(n8148), .op(n8151) );
  nand2_1 U8124 ( .ip1(n8149), .ip2(n8148), .op(n8150) );
  nand2_1 U8125 ( .ip1(n8151), .ip2(n8150), .op(n8152) );
  mux2_1 U8126 ( .ip1(n8154), .ip2(n8153), .s(n8152), .op(\STAGE_1/M10/sum [9]) );
  fulladder U8127 ( .a(n8157), .b(n8156), .ci(n8155), .co(n8148), .s(n8158) );
  inv_1 U8128 ( .ip(n8158), .op(\STAGE_1/M10/sum [8]) );
  fulladder U8129 ( .a(n8161), .b(n8160), .ci(n8159), .co(n8155), .s(n8162) );
  inv_1 U8130 ( .ip(n8162), .op(\STAGE_1/M10/sum [7]) );
  fulladder U8131 ( .a(n8165), .b(n8164), .ci(n8163), .co(n8159), .s(n8166) );
  inv_1 U8132 ( .ip(n8166), .op(\STAGE_1/M10/sum [6]) );
  fulladder U8133 ( .a(n8169), .b(n8168), .ci(n8167), .co(n8163), .s(n8170) );
  inv_1 U8134 ( .ip(n8170), .op(\STAGE_1/M10/sum [5]) );
  fulladder U8135 ( .a(n8173), .b(n8172), .ci(n8171), .co(n8167), .s(n8174) );
  inv_1 U8136 ( .ip(n8174), .op(\STAGE_1/M10/sum [4]) );
  nand2_1 U8137 ( .ip1(n8175), .ip2(column[158]), .op(n8184) );
  nor3_1 U8138 ( .ip1(n8180), .ip2(n8177), .ip3(n8176), .op(n8178) );
  nor2_1 U8139 ( .ip1(n8179), .ip2(n8178), .op(n8182) );
  nor2_1 U8140 ( .ip1(column[158]), .ip2(column[159]), .op(n8181) );
  not_ab_or_c_or_d U8141 ( .ip1(column[158]), .ip2(column[159]), .ip3(n8181), 
        .ip4(n8180), .op(n8186) );
  fulladder U8142 ( .a(n8184), .b(n8183), .ci(n8182), .co(n8185), .s(
        \STAGE_1/M10/sum [14]) );
  xnor2_1 U8143 ( .ip1(n8186), .ip2(n8185), .op(\STAGE_1/M10/sum [15]) );
  inv_1 U8144 ( .ip(\CNTRL/count_layer1_784Q [3]), .op(n8203) );
  nand3_1 U8145 ( .ip1(\CNTRL/count_layer1_784Q [0]), .ip2(
        \CNTRL/count_layer1_784Q [1]), .ip3(\CNTRL/count_layer1_784Q [2]), 
        .op(n8202) );
  nor2_1 U8146 ( .ip1(n8203), .ip2(n8202), .op(n8207) );
  nand4_1 U8147 ( .ip1(n8187), .ip2(\CNTRL/count_layer1_784Q [8]), .ip3(
        \CNTRL/count_layer1_784Q [9]), .ip4(n8207), .op(n8295) );
  inv_1 U8148 ( .ip(n8295), .op(n8298) );
  inv_1 U8149 ( .ip(\CNTRL/count_10_2Q [2]), .op(n8256) );
  inv_1 U8150 ( .ip(\CNTRL/count_10_2Q [1]), .op(n8255) );
  and4_1 U8151 ( .ip1(n8256), .ip2(n8255), .ip3(\CNTRL/count_10_2Q [0]), .ip4(
        \CNTRL/count_10_2Q [3]), .op(n8253) );
  or2_1 U8152 ( .ip1(n8253), .ip2(n9445), .op(n8190) );
  nand4_1 U8153 ( .ip1(\CNTRL/count_10Q [0]), .ip2(\CNTRL/count_10Q [3]), 
        .ip3(n8282), .ip4(n8280), .op(n8268) );
  inv_1 U8154 ( .ip(n8268), .op(n8188) );
  or2_1 U8155 ( .ip1(n8188), .ip2(n9445), .op(n8189) );
  nand2_1 U8156 ( .ip1(n8190), .ip2(n8189), .op(n8194) );
  nor2_1 U8157 ( .ip1(\CNTRL/count_layer1_200Q [0]), .ip2(
        \CNTRL/count_layer1_200Q [1]), .op(n8192) );
  inv_1 U8158 ( .ip(\CNTRL/count_layer1_200Q [3]), .op(n8303) );
  inv_1 U8159 ( .ip(\CNTRL/count_layer1_200Q [6]), .op(n8310) );
  nor4_1 U8160 ( .ip1(\CNTRL/count_layer1_200Q [5]), .ip2(
        \CNTRL/count_layer1_200Q [4]), .ip3(n8303), .ip4(n8310), .op(n8191) );
  inv_1 U8161 ( .ip(\CNTRL/count_layer1_200Q [2]), .op(n8299) );
  nand4_1 U8162 ( .ip1(\CNTRL/count_layer1_200Q [7]), .ip2(n8192), .ip3(n8191), 
        .ip4(n8299), .op(n8197) );
  nand2_1 U8163 ( .ip1(\CNTRL/count_20Q [0]), .ip2(\CNTRL/count_20Q [1]), .op(
        n8240) );
  inv_1 U8164 ( .ip(n8240), .op(n8234) );
  nand3_1 U8165 ( .ip1(\CNTRL/count_20Q [4]), .ip2(n8336), .ip3(n8234), .op(
        n8265) );
  nor4_1 U8166 ( .ip1(n8802), .ip2(n8268), .ip3(n8197), .ip4(n8265), .op(n8193) );
  or2_1 U8167 ( .ip1(n8194), .ip2(n8193), .op(n8229) );
  not_ab_or_c_or_d U8168 ( .ip1(\CNTRL/currentState [1]), .ip2(n8195), .ip3(
        n8298), .ip4(n8229), .op(n8196) );
  nor2_1 U8169 ( .ip1(reset), .ip2(n8196), .op(n4039) );
  nor2_1 U8170 ( .ip1(reset), .ip2(n8298), .op(n8296) );
  nand2_1 U8171 ( .ip1(n8296), .ip2(n8197), .op(n8217) );
  nor2_1 U8172 ( .ip1(\CNTRL/count_layer1_784Q [0]), .ip2(n8217), .op(
        \CNTRL/N233 ) );
  and2_1 U8173 ( .ip1(\CNTRL/count_layer1_784Q [0]), .ip2(
        \CNTRL/count_layer1_784Q [1]), .op(n8199) );
  nor3_1 U8174 ( .ip1(n8198), .ip2(n8199), .ip3(n8217), .op(\CNTRL/N234 ) );
  nor2_1 U8175 ( .ip1(\CNTRL/count_layer1_784Q [2]), .ip2(n8199), .op(n8201)
         );
  inv_1 U8176 ( .ip(n8202), .op(n8200) );
  nor3_1 U8177 ( .ip1(n8201), .ip2(n8200), .ip3(n8217), .op(\CNTRL/N235 ) );
  not_ab_or_c_or_d U8178 ( .ip1(n8203), .ip2(n8202), .ip3(n8207), .ip4(n8217), 
        .op(\CNTRL/N236 ) );
  inv_1 U8179 ( .ip(\CNTRL/count_layer1_784Q [4]), .op(n8205) );
  inv_1 U8180 ( .ip(n8207), .op(n8204) );
  nor2_1 U8181 ( .ip1(n8205), .ip2(n8204), .op(n8206) );
  not_ab_or_c_or_d U8182 ( .ip1(n8205), .ip2(n8204), .ip3(n8206), .ip4(n8217), 
        .op(\CNTRL/N237 ) );
  nor2_1 U8183 ( .ip1(\CNTRL/count_layer1_784Q [5]), .ip2(n8206), .op(n8209)
         );
  nand3_1 U8184 ( .ip1(\CNTRL/count_layer1_784Q [4]), .ip2(
        \CNTRL/count_layer1_784Q [5]), .ip3(n8207), .op(n8210) );
  inv_1 U8185 ( .ip(n8210), .op(n8208) );
  nor3_1 U8186 ( .ip1(n8209), .ip2(n8208), .ip3(n8217), .op(\CNTRL/N238 ) );
  inv_1 U8187 ( .ip(\CNTRL/count_layer1_784Q [6]), .op(n8211) );
  nor2_1 U8188 ( .ip1(n8211), .ip2(n8210), .op(n8212) );
  not_ab_or_c_or_d U8189 ( .ip1(n8211), .ip2(n8210), .ip3(n8212), .ip4(n8217), 
        .op(\CNTRL/N239 ) );
  nor2_1 U8190 ( .ip1(\CNTRL/count_layer1_784Q [7]), .ip2(n8212), .op(n8213)
         );
  nand2_1 U8191 ( .ip1(\CNTRL/count_layer1_784Q [7]), .ip2(n8212), .op(n8214)
         );
  inv_1 U8192 ( .ip(n8214), .op(n8220) );
  nor3_1 U8193 ( .ip1(n8213), .ip2(n8220), .ip3(n8217), .op(\CNTRL/N240 ) );
  inv_1 U8194 ( .ip(\CNTRL/count_layer1_784Q [8]), .op(n8215) );
  nor2_1 U8195 ( .ip1(n8215), .ip2(n8214), .op(n8216) );
  not_ab_or_c_or_d U8196 ( .ip1(n8215), .ip2(n8214), .ip3(n8216), .ip4(n8217), 
        .op(\CNTRL/N241 ) );
  and2_1 U8197 ( .ip1(\CNTRL/count_layer1_784Q [8]), .ip2(
        \CNTRL/count_layer1_784Q [9]), .op(n8219) );
  nor2_1 U8198 ( .ip1(\CNTRL/count_layer1_784Q [9]), .ip2(n8216), .op(n8218)
         );
  not_ab_or_c_or_d U8199 ( .ip1(n8220), .ip2(n8219), .ip3(n8218), .ip4(n8217), 
        .op(\CNTRL/N242 ) );
  inv_1 U8200 ( .ip(\CNTRL/count_20Q [2]), .op(n8789) );
  inv_1 U8201 ( .ip(\CNTRL/count_20Q [3]), .op(n8795) );
  inv_1 U8202 ( .ip(reset), .op(n8267) );
  nand2_1 U8203 ( .ip1(\CNTRL/currentState [1]), .ip2(n8223), .op(n8221) );
  nand2_1 U8204 ( .ip1(n8802), .ip2(n8221), .op(n8222) );
  nand2_1 U8205 ( .ip1(n8267), .ip2(n8222), .op(n8233) );
  nor4_1 U8206 ( .ip1(n8789), .ip2(n8795), .ip3(n8240), .ip4(n8233), .op(n8226) );
  nor3_1 U8207 ( .ip1(n8223), .ip2(reset), .ip3(n8793), .op(n8270) );
  inv_1 U8208 ( .ip(n8270), .op(n8238) );
  inv_1 U8209 ( .ip(n8233), .op(n8232) );
  nand2_1 U8210 ( .ip1(n8265), .ip2(n8232), .op(n8239) );
  inv_1 U8211 ( .ip(n8239), .op(n8271) );
  nor2_1 U8212 ( .ip1(n8789), .ip2(n8240), .op(n8244) );
  nand2_1 U8213 ( .ip1(\CNTRL/count_20Q [3]), .ip2(n8244), .op(n8224) );
  nand2_1 U8214 ( .ip1(n8271), .ip2(n8224), .op(n8225) );
  nand2_1 U8215 ( .ip1(n8238), .ip2(n8225), .op(n8243) );
  mux2_1 U8216 ( .ip1(n8226), .ip2(n8243), .s(\CNTRL/count_20Q [4]), .op(n4043) );
  nor2_1 U8217 ( .ip1(n8268), .ip2(n8265), .op(n8228) );
  nand2_1 U8218 ( .ip1(\CNTRL/currentState [0]), .ip2(\CNTRL/currentState [1]), 
        .op(n8272) );
  inv_1 U8219 ( .ip(n8272), .op(n8227) );
  not_ab_or_c_or_d U8220 ( .ip1(n8810), .ip2(n8228), .ip3(n8227), .ip4(n8807), 
        .op(n8230) );
  nor3_1 U8221 ( .ip1(n8230), .ip2(n8229), .ip3(weight2_loadNextRow), .op(
        n8231) );
  nor2_1 U8222 ( .ip1(reset), .ip2(n8231), .op(n4041) );
  mux2_1 U8223 ( .ip1(n8232), .ip2(n8270), .s(\CNTRL/count_20Q [0]), .op(n4038) );
  nor2_1 U8224 ( .ip1(n8801), .ip2(n8238), .op(n8237) );
  inv_1 U8225 ( .ip(\CNTRL/count_20Q [0]), .op(n8235) );
  not_ab_or_c_or_d U8226 ( .ip1(n8235), .ip2(n8801), .ip3(n8234), .ip4(n8233), 
        .op(n8236) );
  or2_1 U8227 ( .ip1(n8237), .ip2(n8236), .op(n4037) );
  nor2_1 U8228 ( .ip1(n8789), .ip2(n8238), .op(n8242) );
  not_ab_or_c_or_d U8229 ( .ip1(n8789), .ip2(n8240), .ip3(n8244), .ip4(n8239), 
        .op(n8241) );
  or2_1 U8230 ( .ip1(n8242), .ip2(n8241), .op(n4036) );
  inv_1 U8231 ( .ip(n8243), .op(n8248) );
  or2_1 U8232 ( .ip1(n8271), .ip2(\CNTRL/count_20Q [3]), .op(n8246) );
  or2_1 U8233 ( .ip1(n8244), .ip2(\CNTRL/count_20Q [3]), .op(n8245) );
  nand2_1 U8234 ( .ip1(n8246), .ip2(n8245), .op(n8247) );
  nor2_1 U8235 ( .ip1(n8248), .ip2(n8247), .op(n4035) );
  nor2_1 U8236 ( .ip1(n9445), .ip2(n8268), .op(n8250) );
  nor2_1 U8237 ( .ip1(\CNTRL/count_10_2Q [0]), .ip2(n8250), .op(n8249) );
  not_ab_or_c_or_d U8238 ( .ip1(\CNTRL/count_10_2Q [0]), .ip2(n8250), .ip3(
        reset), .ip4(n8249), .op(n4034) );
  or2_1 U8239 ( .ip1(\CNTRL/count_10_2Q [0]), .ip2(reset), .op(n8252) );
  or2_1 U8240 ( .ip1(n8250), .ip2(reset), .op(n8251) );
  nand2_1 U8241 ( .ip1(n8252), .ip2(n8251), .op(n8254) );
  nor2_1 U8242 ( .ip1(n8255), .ip2(n8254), .op(n8258) );
  nor2_1 U8243 ( .ip1(reset), .ip2(n8253), .op(n8260) );
  nor2_1 U8244 ( .ip1(n8260), .ip2(n8254), .op(n8263) );
  not_ab_or_c_or_d U8245 ( .ip1(n8255), .ip2(n8254), .ip3(n8258), .ip4(n8263), 
        .op(n4033) );
  inv_1 U8246 ( .ip(n8258), .op(n8257) );
  nor2_1 U8247 ( .ip1(n8257), .ip2(n8256), .op(n8264) );
  or2_1 U8248 ( .ip1(n8258), .ip2(\CNTRL/count_10_2Q [2]), .op(n8259) );
  nand2_1 U8249 ( .ip1(n8260), .ip2(n8259), .op(n8261) );
  nor2_1 U8250 ( .ip1(n8264), .ip2(n8261), .op(n4032) );
  nor2_1 U8251 ( .ip1(\CNTRL/count_10_2Q [3]), .ip2(n8264), .op(n8262) );
  not_ab_or_c_or_d U8252 ( .ip1(\CNTRL/count_10_2Q [3]), .ip2(n8264), .ip3(
        n8263), .ip4(n8262), .op(n4031) );
  or2_1 U8253 ( .ip1(n8802), .ip2(n8265), .op(n8266) );
  nand2_1 U8254 ( .ip1(n9445), .ip2(n8266), .op(n8269) );
  nand3_1 U8255 ( .ip1(n8269), .ip2(n8268), .ip3(n8267), .op(n8287) );
  or2_1 U8256 ( .ip1(n8270), .ip2(n8271), .op(n8274) );
  or2_1 U8257 ( .ip1(n8272), .ip2(n8271), .op(n8273) );
  nand2_1 U8258 ( .ip1(n8274), .ip2(n8273), .op(n8286) );
  mux2_1 U8259 ( .ip1(n8287), .ip2(n8286), .s(\CNTRL/count_10Q [0]), .op(n8275) );
  inv_1 U8260 ( .ip(n8275), .op(n4030) );
  or2_1 U8261 ( .ip1(n8287), .ip2(\CNTRL/count_10Q [0]), .op(n8276) );
  nand2_1 U8262 ( .ip1(n8286), .ip2(n8276), .op(n8278) );
  inv_1 U8263 ( .ip(\CNTRL/count_10Q [0]), .op(n8279) );
  nor2_1 U8264 ( .ip1(n8279), .ip2(n8287), .op(n8277) );
  mux2_1 U8265 ( .ip1(n8278), .ip2(n8277), .s(n8280), .op(n4029) );
  nor2_1 U8266 ( .ip1(n8286), .ip2(n8282), .op(n8284) );
  nand2_1 U8267 ( .ip1(\CNTRL/count_10Q [1]), .ip2(\CNTRL/count_10Q [0]), .op(
        n8281) );
  nor3_1 U8268 ( .ip1(n8282), .ip2(n8280), .ip3(n8279), .op(n8289) );
  not_ab_or_c_or_d U8269 ( .ip1(n8282), .ip2(n8281), .ip3(n8289), .ip4(n8287), 
        .op(n8283) );
  or2_1 U8270 ( .ip1(n8284), .ip2(n8283), .op(n4028) );
  nor2_1 U8271 ( .ip1(n8286), .ip2(n8285), .op(n8291) );
  nor2_1 U8272 ( .ip1(\CNTRL/count_10Q [3]), .ip2(n8289), .op(n8288) );
  not_ab_or_c_or_d U8273 ( .ip1(\CNTRL/count_10Q [3]), .ip2(n8289), .ip3(n8288), .ip4(n8287), .op(n8290) );
  or2_1 U8274 ( .ip1(n8291), .ip2(n8290), .op(n4027) );
  inv_1 U8275 ( .ip(\CNTRL/count_layer1_200Q [1]), .op(n8294) );
  nand2_1 U8276 ( .ip1(n8298), .ip2(\CNTRL/count_layer1_200Q [0]), .op(n8293)
         );
  nor2_1 U8277 ( .ip1(n8294), .ip2(n8293), .op(n8292) );
  not_ab_or_c_or_d U8278 ( .ip1(n8294), .ip2(n8293), .ip3(reset), .ip4(n8292), 
        .op(n4026) );
  nor2_1 U8279 ( .ip1(reset), .ip2(n8295), .op(n8297) );
  mux2_1 U8280 ( .ip1(n8297), .ip2(n8296), .s(\CNTRL/count_layer1_200Q [0]), 
        .op(n4025) );
  nand3_1 U8281 ( .ip1(\CNTRL/count_layer1_200Q [0]), .ip2(
        \CNTRL/count_layer1_200Q [1]), .ip3(n8298), .op(n8300) );
  nor2_1 U8282 ( .ip1(n8300), .ip2(n8299), .op(n8301) );
  not_ab_or_c_or_d U8283 ( .ip1(n8300), .ip2(n8299), .ip3(reset), .ip4(n8301), 
        .op(n4024) );
  inv_1 U8284 ( .ip(n8301), .op(n8304) );
  nand2_1 U8285 ( .ip1(n8301), .ip2(\CNTRL/count_layer1_200Q [3]), .op(n8306)
         );
  inv_1 U8286 ( .ip(n8306), .op(n8302) );
  not_ab_or_c_or_d U8287 ( .ip1(n8304), .ip2(n8303), .ip3(reset), .ip4(n8302), 
        .op(n4023) );
  inv_1 U8288 ( .ip(\CNTRL/count_layer1_200Q [4]), .op(n8305) );
  nor2_1 U8289 ( .ip1(n8306), .ip2(n8305), .op(n8307) );
  not_ab_or_c_or_d U8290 ( .ip1(n8306), .ip2(n8305), .ip3(reset), .ip4(n8307), 
        .op(n4022) );
  nor2_1 U8291 ( .ip1(n8307), .ip2(\CNTRL/count_layer1_200Q [5]), .op(n8309)
         );
  nand2_1 U8292 ( .ip1(n8307), .ip2(\CNTRL/count_layer1_200Q [5]), .op(n8311)
         );
  inv_1 U8293 ( .ip(n8311), .op(n8308) );
  nor3_1 U8294 ( .ip1(n8309), .ip2(reset), .ip3(n8308), .op(n4021) );
  nor2_1 U8295 ( .ip1(n8311), .ip2(n8310), .op(n8313) );
  not_ab_or_c_or_d U8296 ( .ip1(n8311), .ip2(n8310), .ip3(reset), .ip4(n8313), 
        .op(n4020) );
  nor2_1 U8297 ( .ip1(\CNTRL/count_layer1_200Q [7]), .ip2(n8313), .op(n8312)
         );
  not_ab_or_c_or_d U8298 ( .ip1(\CNTRL/count_layer1_200Q [7]), .ip2(n8313), 
        .ip3(reset), .ip4(n8312), .op(n4019) );
  nor2_1 U8299 ( .ip1(\CNTRL/count_20Q [1]), .ip2(n8314), .op(n10052) );
  inv_1 U8300 ( .ip(\CNTRL/count_20Q [4]), .op(n8809) );
  nand2_1 U8301 ( .ip1(n8801), .ip2(n8809), .op(n8330) );
  nand3_1 U8302 ( .ip1(\CNTRL/count_20Q [2]), .ip2(\CNTRL/count_20Q [3]), 
        .ip3(n8328), .op(n8318) );
  nor2_1 U8303 ( .ip1(n8330), .ip2(n8318), .op(n10044) );
  nand2_1 U8304 ( .ip1(\ROUTEDATA/regData [96]), .ip2(n10044), .op(n8316) );
  nand2_1 U8305 ( .ip1(\ROUTEDATA/regData [144]), .ip2(n8523), .op(n8315) );
  nand2_1 U8306 ( .ip1(n8316), .ip2(n8315), .op(n8324) );
  nand3_1 U8307 ( .ip1(\CNTRL/count_20Q [3]), .ip2(n8328), .ip3(n8789), .op(
        n8317) );
  nor2_1 U8308 ( .ip1(n8330), .ip2(n8317), .op(n10036) );
  nand2_1 U8309 ( .ip1(n10036), .ip2(\ROUTEDATA/regData [64]), .op(n8322) );
  nand2_1 U8310 ( .ip1(\CNTRL/count_20Q [1]), .ip2(n8809), .op(n8325) );
  nor2_1 U8311 ( .ip1(n8317), .ip2(n8325), .op(n10040) );
  nand2_1 U8312 ( .ip1(n10040), .ip2(\ROUTEDATA/regData [80]), .op(n8321) );
  nor2_1 U8313 ( .ip1(n8325), .ip2(n8318), .op(n10048) );
  nand2_1 U8314 ( .ip1(n10048), .ip2(\ROUTEDATA/regData [112]), .op(n8320) );
  nand3_1 U8315 ( .ip1(\CNTRL/count_20Q [2]), .ip2(n8328), .ip3(n8795), .op(
        n8329) );
  nor2_1 U8316 ( .ip1(n8325), .ip2(n8329), .op(n10032) );
  nand2_1 U8317 ( .ip1(n10032), .ip2(\ROUTEDATA/regData [48]), .op(n8319) );
  nand4_1 U8318 ( .ip1(n8322), .ip2(n8321), .ip3(n8320), .ip4(n8319), .op(
        n8323) );
  not_ab_or_c_or_d U8319 ( .ip1(n10052), .ip2(\ROUTEDATA/regData [128]), .ip3(
        n8324), .ip4(n8323), .op(n8334) );
  inv_1 U8320 ( .ip(n8328), .op(n8335) );
  inv_1 U8321 ( .ip(n8336), .op(n8326) );
  nor3_1 U8322 ( .ip1(n8335), .ip2(n8326), .ip3(n8325), .op(n10023) );
  nand2_1 U8323 ( .ip1(n10023), .ip2(\ROUTEDATA/regData [16]), .op(n8333) );
  or3_1 U8324 ( .ip1(\CNTRL/count_20Q [2]), .ip2(n8330), .ip3(
        \CNTRL/count_20Q [3]), .op(n8327) );
  nand2_1 U8325 ( .ip1(n8328), .ip2(n8327), .op(n10435) );
  nand2_1 U8326 ( .ip1(\ROUTEDATA/regData [0]), .ip2(n10435), .op(n8332) );
  nor2_1 U8327 ( .ip1(n8330), .ip2(n8329), .op(n10028) );
  nand2_1 U8328 ( .ip1(n10028), .ip2(\ROUTEDATA/regData [32]), .op(n8331) );
  nand4_1 U8329 ( .ip1(n8334), .ip2(n8333), .ip3(n8332), .ip4(n8331), .op(
        n8338) );
  nor3_1 U8330 ( .ip1(n8336), .ip2(n8809), .ip3(n8335), .op(n8337) );
  nor2_1 U8331 ( .ip1(n8337), .ip2(n10053), .op(n8534) );
  mux2_1 U8332 ( .ip1(m2DataIn[0]), .ip2(n8338), .s(n8534), .op(n4018) );
  nand2_1 U8333 ( .ip1(\ROUTEDATA/regData [33]), .ip2(n10028), .op(n8340) );
  nand2_1 U8334 ( .ip1(\ROUTEDATA/regData [81]), .ip2(n10040), .op(n8339) );
  nand2_1 U8335 ( .ip1(n8340), .ip2(n8339), .op(n8346) );
  nand2_1 U8336 ( .ip1(n10052), .ip2(\ROUTEDATA/regData [129]), .op(n8344) );
  nand2_1 U8337 ( .ip1(n8523), .ip2(\ROUTEDATA/regData [145]), .op(n8343) );
  nand2_1 U8338 ( .ip1(n10032), .ip2(\ROUTEDATA/regData [49]), .op(n8342) );
  nand2_1 U8339 ( .ip1(n10048), .ip2(\ROUTEDATA/regData [113]), .op(n8341) );
  nand4_1 U8340 ( .ip1(n8344), .ip2(n8343), .ip3(n8342), .ip4(n8341), .op(
        n8345) );
  not_ab_or_c_or_d U8341 ( .ip1(n10036), .ip2(\ROUTEDATA/regData [65]), .ip3(
        n8346), .ip4(n8345), .op(n8350) );
  nand2_1 U8342 ( .ip1(n10023), .ip2(\ROUTEDATA/regData [17]), .op(n8349) );
  nand2_1 U8343 ( .ip1(n10044), .ip2(\ROUTEDATA/regData [97]), .op(n8348) );
  nand2_1 U8344 ( .ip1(\ROUTEDATA/regData [1]), .ip2(n10435), .op(n8347) );
  nand4_1 U8345 ( .ip1(n8350), .ip2(n8349), .ip3(n8348), .ip4(n8347), .op(
        n8351) );
  mux2_1 U8346 ( .ip1(m2DataIn[1]), .ip2(n8351), .s(n8534), .op(n4017) );
  nand2_1 U8347 ( .ip1(\ROUTEDATA/regData [98]), .ip2(n10044), .op(n8353) );
  nand2_1 U8348 ( .ip1(\ROUTEDATA/regData [146]), .ip2(n8523), .op(n8352) );
  nand2_1 U8349 ( .ip1(n8353), .ip2(n8352), .op(n8359) );
  nand2_1 U8350 ( .ip1(n10036), .ip2(\ROUTEDATA/regData [66]), .op(n8357) );
  nand2_1 U8351 ( .ip1(n10040), .ip2(\ROUTEDATA/regData [82]), .op(n8356) );
  nand2_1 U8352 ( .ip1(n10032), .ip2(\ROUTEDATA/regData [50]), .op(n8355) );
  nand2_1 U8353 ( .ip1(n10048), .ip2(\ROUTEDATA/regData [114]), .op(n8354) );
  nand4_1 U8354 ( .ip1(n8357), .ip2(n8356), .ip3(n8355), .ip4(n8354), .op(
        n8358) );
  not_ab_or_c_or_d U8355 ( .ip1(n10052), .ip2(\ROUTEDATA/regData [130]), .ip3(
        n8359), .ip4(n8358), .op(n8363) );
  nand2_1 U8356 ( .ip1(\ROUTEDATA/regData [2]), .ip2(n10435), .op(n8362) );
  nand2_1 U8357 ( .ip1(n10028), .ip2(\ROUTEDATA/regData [34]), .op(n8361) );
  nand2_1 U8358 ( .ip1(n10023), .ip2(\ROUTEDATA/regData [18]), .op(n8360) );
  nand4_1 U8359 ( .ip1(n8363), .ip2(n8362), .ip3(n8361), .ip4(n8360), .op(
        n8364) );
  mux2_1 U8360 ( .ip1(m2DataIn[2]), .ip2(n8364), .s(n8534), .op(n4016) );
  nand2_1 U8361 ( .ip1(\ROUTEDATA/regData [51]), .ip2(n10032), .op(n8366) );
  nand2_1 U8362 ( .ip1(\ROUTEDATA/regData [83]), .ip2(n10040), .op(n8365) );
  nand2_1 U8363 ( .ip1(n8366), .ip2(n8365), .op(n8372) );
  nand2_1 U8364 ( .ip1(n8523), .ip2(\ROUTEDATA/regData [147]), .op(n8370) );
  nand2_1 U8365 ( .ip1(n10052), .ip2(\ROUTEDATA/regData [131]), .op(n8369) );
  nand2_1 U8366 ( .ip1(n10044), .ip2(\ROUTEDATA/regData [99]), .op(n8368) );
  nand2_1 U8367 ( .ip1(n10028), .ip2(\ROUTEDATA/regData [35]), .op(n8367) );
  nand4_1 U8368 ( .ip1(n8370), .ip2(n8369), .ip3(n8368), .ip4(n8367), .op(
        n8371) );
  not_ab_or_c_or_d U8369 ( .ip1(n10036), .ip2(\ROUTEDATA/regData [67]), .ip3(
        n8372), .ip4(n8371), .op(n8376) );
  nand2_1 U8370 ( .ip1(n10048), .ip2(\ROUTEDATA/regData [115]), .op(n8375) );
  nand2_1 U8371 ( .ip1(\ROUTEDATA/regData [3]), .ip2(n10435), .op(n8374) );
  nand2_1 U8372 ( .ip1(n10023), .ip2(\ROUTEDATA/regData [19]), .op(n8373) );
  nand4_1 U8373 ( .ip1(n8376), .ip2(n8375), .ip3(n8374), .ip4(n8373), .op(
        n8377) );
  mux2_1 U8374 ( .ip1(m2DataIn[3]), .ip2(n8377), .s(n8534), .op(n4015) );
  nand2_1 U8375 ( .ip1(\ROUTEDATA/regData [100]), .ip2(n10044), .op(n8379) );
  nand2_1 U8376 ( .ip1(\ROUTEDATA/regData [148]), .ip2(n8523), .op(n8378) );
  nand2_1 U8377 ( .ip1(n8379), .ip2(n8378), .op(n8385) );
  nand2_1 U8378 ( .ip1(n10040), .ip2(\ROUTEDATA/regData [84]), .op(n8383) );
  nand2_1 U8379 ( .ip1(n10052), .ip2(\ROUTEDATA/regData [132]), .op(n8382) );
  nand2_1 U8380 ( .ip1(n10028), .ip2(\ROUTEDATA/regData [36]), .op(n8381) );
  nand2_1 U8381 ( .ip1(n10048), .ip2(\ROUTEDATA/regData [116]), .op(n8380) );
  nand4_1 U8382 ( .ip1(n8383), .ip2(n8382), .ip3(n8381), .ip4(n8380), .op(
        n8384) );
  not_ab_or_c_or_d U8383 ( .ip1(n10036), .ip2(\ROUTEDATA/regData [68]), .ip3(
        n8385), .ip4(n8384), .op(n8389) );
  nand2_1 U8384 ( .ip1(\ROUTEDATA/regData [4]), .ip2(n10435), .op(n8388) );
  nand2_1 U8385 ( .ip1(n10032), .ip2(\ROUTEDATA/regData [52]), .op(n8387) );
  nand2_1 U8386 ( .ip1(n10023), .ip2(\ROUTEDATA/regData [20]), .op(n8386) );
  nand4_1 U8387 ( .ip1(n8389), .ip2(n8388), .ip3(n8387), .ip4(n8386), .op(
        n8390) );
  mux2_1 U8388 ( .ip1(m2DataIn[4]), .ip2(n8390), .s(n8534), .op(n4014) );
  nand2_1 U8389 ( .ip1(\ROUTEDATA/regData [101]), .ip2(n10044), .op(n8392) );
  nand2_1 U8390 ( .ip1(\ROUTEDATA/regData [85]), .ip2(n10040), .op(n8391) );
  nand2_1 U8391 ( .ip1(n8392), .ip2(n8391), .op(n8398) );
  nand2_1 U8392 ( .ip1(n8523), .ip2(\ROUTEDATA/regData [149]), .op(n8396) );
  nand2_1 U8393 ( .ip1(n10052), .ip2(\ROUTEDATA/regData [133]), .op(n8395) );
  nand2_1 U8394 ( .ip1(n10028), .ip2(\ROUTEDATA/regData [37]), .op(n8394) );
  nand2_1 U8395 ( .ip1(n10048), .ip2(\ROUTEDATA/regData [117]), .op(n8393) );
  nand4_1 U8396 ( .ip1(n8396), .ip2(n8395), .ip3(n8394), .ip4(n8393), .op(
        n8397) );
  not_ab_or_c_or_d U8397 ( .ip1(n10036), .ip2(\ROUTEDATA/regData [69]), .ip3(
        n8398), .ip4(n8397), .op(n8402) );
  nand2_1 U8398 ( .ip1(n10023), .ip2(\ROUTEDATA/regData [21]), .op(n8401) );
  nand2_1 U8399 ( .ip1(\ROUTEDATA/regData [5]), .ip2(n10435), .op(n8400) );
  nand2_1 U8400 ( .ip1(n10032), .ip2(\ROUTEDATA/regData [53]), .op(n8399) );
  nand4_1 U8401 ( .ip1(n8402), .ip2(n8401), .ip3(n8400), .ip4(n8399), .op(
        n8403) );
  mux2_1 U8402 ( .ip1(m2DataIn[5]), .ip2(n8403), .s(n8534), .op(n4013) );
  nand2_1 U8403 ( .ip1(\ROUTEDATA/regData [150]), .ip2(n8523), .op(n8405) );
  nand2_1 U8404 ( .ip1(\ROUTEDATA/regData [118]), .ip2(n10048), .op(n8404) );
  nand2_1 U8405 ( .ip1(n8405), .ip2(n8404), .op(n8411) );
  nand2_1 U8406 ( .ip1(n10052), .ip2(\ROUTEDATA/regData [134]), .op(n8409) );
  nand2_1 U8407 ( .ip1(n10040), .ip2(\ROUTEDATA/regData [86]), .op(n8408) );
  nand2_1 U8408 ( .ip1(n10044), .ip2(\ROUTEDATA/regData [102]), .op(n8407) );
  nand2_1 U8409 ( .ip1(n10028), .ip2(\ROUTEDATA/regData [38]), .op(n8406) );
  nand4_1 U8410 ( .ip1(n8409), .ip2(n8408), .ip3(n8407), .ip4(n8406), .op(
        n8410) );
  not_ab_or_c_or_d U8411 ( .ip1(n10036), .ip2(\ROUTEDATA/regData [70]), .ip3(
        n8411), .ip4(n8410), .op(n8415) );
  nand2_1 U8412 ( .ip1(\ROUTEDATA/regData [6]), .ip2(n10435), .op(n8414) );
  nand2_1 U8413 ( .ip1(n10032), .ip2(\ROUTEDATA/regData [54]), .op(n8413) );
  nand2_1 U8414 ( .ip1(n10023), .ip2(\ROUTEDATA/regData [22]), .op(n8412) );
  nand4_1 U8415 ( .ip1(n8415), .ip2(n8414), .ip3(n8413), .ip4(n8412), .op(
        n8416) );
  mux2_1 U8416 ( .ip1(m2DataIn[6]), .ip2(n8416), .s(n8534), .op(n4012) );
  nand2_1 U8417 ( .ip1(\ROUTEDATA/regData [103]), .ip2(n10044), .op(n8418) );
  nand2_1 U8418 ( .ip1(\ROUTEDATA/regData [151]), .ip2(n8523), .op(n8417) );
  nand2_1 U8419 ( .ip1(n8418), .ip2(n8417), .op(n8424) );
  nand2_1 U8420 ( .ip1(n10052), .ip2(\ROUTEDATA/regData [135]), .op(n8422) );
  nand2_1 U8421 ( .ip1(n10040), .ip2(\ROUTEDATA/regData [87]), .op(n8421) );
  nand2_1 U8422 ( .ip1(n10048), .ip2(\ROUTEDATA/regData [119]), .op(n8420) );
  nand2_1 U8423 ( .ip1(n10028), .ip2(\ROUTEDATA/regData [39]), .op(n8419) );
  nand4_1 U8424 ( .ip1(n8422), .ip2(n8421), .ip3(n8420), .ip4(n8419), .op(
        n8423) );
  not_ab_or_c_or_d U8425 ( .ip1(n10036), .ip2(\ROUTEDATA/regData [71]), .ip3(
        n8424), .ip4(n8423), .op(n8428) );
  nand2_1 U8426 ( .ip1(\ROUTEDATA/regData [7]), .ip2(n10435), .op(n8427) );
  nand2_1 U8427 ( .ip1(n10032), .ip2(\ROUTEDATA/regData [55]), .op(n8426) );
  nand2_1 U8428 ( .ip1(n10023), .ip2(\ROUTEDATA/regData [23]), .op(n8425) );
  nand4_1 U8429 ( .ip1(n8428), .ip2(n8427), .ip3(n8426), .ip4(n8425), .op(
        n8429) );
  mux2_1 U8430 ( .ip1(m2DataIn[7]), .ip2(n8429), .s(n8534), .op(n4011) );
  nand2_1 U8431 ( .ip1(\ROUTEDATA/regData [152]), .ip2(n8523), .op(n8431) );
  nand2_1 U8432 ( .ip1(\ROUTEDATA/regData [120]), .ip2(n10048), .op(n8430) );
  nand2_1 U8433 ( .ip1(n8431), .ip2(n8430), .op(n8437) );
  nand2_1 U8434 ( .ip1(n10052), .ip2(\ROUTEDATA/regData [136]), .op(n8435) );
  nand2_1 U8435 ( .ip1(n10036), .ip2(\ROUTEDATA/regData [72]), .op(n8434) );
  nand2_1 U8436 ( .ip1(n10028), .ip2(\ROUTEDATA/regData [40]), .op(n8433) );
  nand2_1 U8437 ( .ip1(n10044), .ip2(\ROUTEDATA/regData [104]), .op(n8432) );
  nand4_1 U8438 ( .ip1(n8435), .ip2(n8434), .ip3(n8433), .ip4(n8432), .op(
        n8436) );
  not_ab_or_c_or_d U8439 ( .ip1(n10040), .ip2(\ROUTEDATA/regData [88]), .ip3(
        n8437), .ip4(n8436), .op(n8441) );
  nand2_1 U8440 ( .ip1(\ROUTEDATA/regData [8]), .ip2(n10435), .op(n8440) );
  nand2_1 U8441 ( .ip1(n10032), .ip2(\ROUTEDATA/regData [56]), .op(n8439) );
  nand2_1 U8442 ( .ip1(n10023), .ip2(\ROUTEDATA/regData [24]), .op(n8438) );
  nand4_1 U8443 ( .ip1(n8441), .ip2(n8440), .ip3(n8439), .ip4(n8438), .op(
        n8442) );
  mux2_1 U8444 ( .ip1(m2DataIn[8]), .ip2(n8442), .s(n8534), .op(n4010) );
  nand2_1 U8445 ( .ip1(\ROUTEDATA/regData [137]), .ip2(n10052), .op(n8444) );
  nand2_1 U8446 ( .ip1(\ROUTEDATA/regData [41]), .ip2(n10028), .op(n8443) );
  nand2_1 U8447 ( .ip1(n8444), .ip2(n8443), .op(n8450) );
  nand2_1 U8448 ( .ip1(n10036), .ip2(\ROUTEDATA/regData [73]), .op(n8448) );
  nand2_1 U8449 ( .ip1(n8523), .ip2(\ROUTEDATA/regData [153]), .op(n8447) );
  nand2_1 U8450 ( .ip1(n10044), .ip2(\ROUTEDATA/regData [105]), .op(n8446) );
  nand2_1 U8451 ( .ip1(n10048), .ip2(\ROUTEDATA/regData [121]), .op(n8445) );
  nand4_1 U8452 ( .ip1(n8448), .ip2(n8447), .ip3(n8446), .ip4(n8445), .op(
        n8449) );
  not_ab_or_c_or_d U8453 ( .ip1(n10040), .ip2(\ROUTEDATA/regData [89]), .ip3(
        n8450), .ip4(n8449), .op(n8454) );
  nand2_1 U8454 ( .ip1(\ROUTEDATA/regData [9]), .ip2(n10435), .op(n8453) );
  nand2_1 U8455 ( .ip1(n10023), .ip2(\ROUTEDATA/regData [25]), .op(n8452) );
  nand2_1 U8456 ( .ip1(n10032), .ip2(\ROUTEDATA/regData [57]), .op(n8451) );
  nand4_1 U8457 ( .ip1(n8454), .ip2(n8453), .ip3(n8452), .ip4(n8451), .op(
        n8455) );
  mux2_1 U8458 ( .ip1(m2DataIn[9]), .ip2(n8455), .s(n8534), .op(n4009) );
  nand2_1 U8459 ( .ip1(\ROUTEDATA/regData [106]), .ip2(n10044), .op(n8457) );
  nand2_1 U8460 ( .ip1(\ROUTEDATA/regData [154]), .ip2(n8523), .op(n8456) );
  nand2_1 U8461 ( .ip1(n8457), .ip2(n8456), .op(n8463) );
  nand2_1 U8462 ( .ip1(n10040), .ip2(\ROUTEDATA/regData [90]), .op(n8461) );
  nand2_1 U8463 ( .ip1(n10052), .ip2(\ROUTEDATA/regData [138]), .op(n8460) );
  nand2_1 U8464 ( .ip1(n10048), .ip2(\ROUTEDATA/regData [122]), .op(n8459) );
  nand2_1 U8465 ( .ip1(n10032), .ip2(\ROUTEDATA/regData [58]), .op(n8458) );
  nand4_1 U8466 ( .ip1(n8461), .ip2(n8460), .ip3(n8459), .ip4(n8458), .op(
        n8462) );
  not_ab_or_c_or_d U8467 ( .ip1(n10036), .ip2(\ROUTEDATA/regData [74]), .ip3(
        n8463), .ip4(n8462), .op(n8467) );
  nand2_1 U8468 ( .ip1(n10023), .ip2(\ROUTEDATA/regData [26]), .op(n8466) );
  nand2_1 U8469 ( .ip1(\ROUTEDATA/regData [10]), .ip2(n10435), .op(n8465) );
  nand2_1 U8470 ( .ip1(n10028), .ip2(\ROUTEDATA/regData [42]), .op(n8464) );
  nand4_1 U8471 ( .ip1(n8467), .ip2(n8466), .ip3(n8465), .ip4(n8464), .op(
        n8468) );
  mux2_1 U8472 ( .ip1(m2DataIn[10]), .ip2(n8468), .s(n8534), .op(n4008) );
  nand2_1 U8473 ( .ip1(\ROUTEDATA/regData [155]), .ip2(n8523), .op(n8470) );
  nand2_1 U8474 ( .ip1(\ROUTEDATA/regData [139]), .ip2(n10052), .op(n8469) );
  nand2_1 U8475 ( .ip1(n8470), .ip2(n8469), .op(n8476) );
  nand2_1 U8476 ( .ip1(n10036), .ip2(\ROUTEDATA/regData [75]), .op(n8474) );
  nand2_1 U8477 ( .ip1(n10040), .ip2(\ROUTEDATA/regData [91]), .op(n8473) );
  nand2_1 U8478 ( .ip1(n10044), .ip2(\ROUTEDATA/regData [107]), .op(n8472) );
  nand2_1 U8479 ( .ip1(n10028), .ip2(\ROUTEDATA/regData [43]), .op(n8471) );
  nand4_1 U8480 ( .ip1(n8474), .ip2(n8473), .ip3(n8472), .ip4(n8471), .op(
        n8475) );
  not_ab_or_c_or_d U8481 ( .ip1(n10032), .ip2(\ROUTEDATA/regData [59]), .ip3(
        n8476), .ip4(n8475), .op(n8480) );
  nand2_1 U8482 ( .ip1(n10048), .ip2(\ROUTEDATA/regData [123]), .op(n8479) );
  nand2_1 U8483 ( .ip1(\ROUTEDATA/regData [11]), .ip2(n10435), .op(n8478) );
  nand2_1 U8484 ( .ip1(n10023), .ip2(\ROUTEDATA/regData [27]), .op(n8477) );
  nand4_1 U8485 ( .ip1(n8480), .ip2(n8479), .ip3(n8478), .ip4(n8477), .op(
        n8481) );
  mux2_1 U8486 ( .ip1(m2DataIn[11]), .ip2(n8481), .s(n8534), .op(n4007) );
  nand2_1 U8487 ( .ip1(\ROUTEDATA/regData [124]), .ip2(n10048), .op(n8483) );
  nand2_1 U8488 ( .ip1(\ROUTEDATA/regData [92]), .ip2(n10040), .op(n8482) );
  nand2_1 U8489 ( .ip1(n8483), .ip2(n8482), .op(n8489) );
  nand2_1 U8490 ( .ip1(n8523), .ip2(\ROUTEDATA/regData [156]), .op(n8487) );
  nand2_1 U8491 ( .ip1(n10052), .ip2(\ROUTEDATA/regData [140]), .op(n8486) );
  nand2_1 U8492 ( .ip1(n10044), .ip2(\ROUTEDATA/regData [108]), .op(n8485) );
  nand2_1 U8493 ( .ip1(n10028), .ip2(\ROUTEDATA/regData [44]), .op(n8484) );
  nand4_1 U8494 ( .ip1(n8487), .ip2(n8486), .ip3(n8485), .ip4(n8484), .op(
        n8488) );
  not_ab_or_c_or_d U8495 ( .ip1(n10036), .ip2(\ROUTEDATA/regData [76]), .ip3(
        n8489), .ip4(n8488), .op(n8493) );
  nand2_1 U8496 ( .ip1(n10023), .ip2(\ROUTEDATA/regData [28]), .op(n8492) );
  nand2_1 U8497 ( .ip1(n10032), .ip2(\ROUTEDATA/regData [60]), .op(n8491) );
  nand2_1 U8498 ( .ip1(\ROUTEDATA/regData [12]), .ip2(n10435), .op(n8490) );
  nand4_1 U8499 ( .ip1(n8493), .ip2(n8492), .ip3(n8491), .ip4(n8490), .op(
        n8494) );
  mux2_1 U8500 ( .ip1(m2DataIn[12]), .ip2(n8494), .s(n8534), .op(n4006) );
  nand2_1 U8501 ( .ip1(\ROUTEDATA/regData [141]), .ip2(n10052), .op(n8496) );
  nand2_1 U8502 ( .ip1(\ROUTEDATA/regData [45]), .ip2(n10028), .op(n8495) );
  nand2_1 U8503 ( .ip1(n8496), .ip2(n8495), .op(n8502) );
  nand2_1 U8504 ( .ip1(n10040), .ip2(\ROUTEDATA/regData [93]), .op(n8500) );
  nand2_1 U8505 ( .ip1(n8523), .ip2(\ROUTEDATA/regData [157]), .op(n8499) );
  nand2_1 U8506 ( .ip1(n10048), .ip2(\ROUTEDATA/regData [125]), .op(n8498) );
  nand2_1 U8507 ( .ip1(n10044), .ip2(\ROUTEDATA/regData [109]), .op(n8497) );
  nand4_1 U8508 ( .ip1(n8500), .ip2(n8499), .ip3(n8498), .ip4(n8497), .op(
        n8501) );
  not_ab_or_c_or_d U8509 ( .ip1(n10036), .ip2(\ROUTEDATA/regData [77]), .ip3(
        n8502), .ip4(n8501), .op(n8506) );
  nand2_1 U8510 ( .ip1(n10023), .ip2(\ROUTEDATA/regData [29]), .op(n8505) );
  nand2_1 U8511 ( .ip1(n10032), .ip2(\ROUTEDATA/regData [61]), .op(n8504) );
  nand2_1 U8512 ( .ip1(\ROUTEDATA/regData [13]), .ip2(n10435), .op(n8503) );
  nand4_1 U8513 ( .ip1(n8506), .ip2(n8505), .ip3(n8504), .ip4(n8503), .op(
        n8507) );
  mux2_1 U8514 ( .ip1(m2DataIn[13]), .ip2(n8507), .s(n8534), .op(n4005) );
  nand2_1 U8515 ( .ip1(\ROUTEDATA/regData [110]), .ip2(n10044), .op(n8509) );
  nand2_1 U8516 ( .ip1(\ROUTEDATA/regData [142]), .ip2(n10052), .op(n8508) );
  nand2_1 U8517 ( .ip1(n8509), .ip2(n8508), .op(n8515) );
  nand2_1 U8518 ( .ip1(n10036), .ip2(\ROUTEDATA/regData [78]), .op(n8513) );
  nand2_1 U8519 ( .ip1(n8523), .ip2(\ROUTEDATA/regData [158]), .op(n8512) );
  nand2_1 U8520 ( .ip1(n10032), .ip2(\ROUTEDATA/regData [62]), .op(n8511) );
  nand2_1 U8521 ( .ip1(n10028), .ip2(\ROUTEDATA/regData [46]), .op(n8510) );
  nand4_1 U8522 ( .ip1(n8513), .ip2(n8512), .ip3(n8511), .ip4(n8510), .op(
        n8514) );
  not_ab_or_c_or_d U8523 ( .ip1(n10040), .ip2(\ROUTEDATA/regData [94]), .ip3(
        n8515), .ip4(n8514), .op(n8519) );
  nand2_1 U8524 ( .ip1(n10048), .ip2(\ROUTEDATA/regData [126]), .op(n8518) );
  nand2_1 U8525 ( .ip1(n10023), .ip2(\ROUTEDATA/regData [30]), .op(n8517) );
  nand2_1 U8526 ( .ip1(\ROUTEDATA/regData [14]), .ip2(n10435), .op(n8516) );
  nand4_1 U8527 ( .ip1(n8519), .ip2(n8518), .ip3(n8517), .ip4(n8516), .op(
        n8520) );
  mux2_1 U8528 ( .ip1(m2DataIn[14]), .ip2(n8520), .s(n8534), .op(n4004) );
  nand2_1 U8529 ( .ip1(\ROUTEDATA/regData [143]), .ip2(n10052), .op(n8522) );
  nand2_1 U8530 ( .ip1(\ROUTEDATA/regData [127]), .ip2(n10048), .op(n8521) );
  nand2_1 U8531 ( .ip1(n8522), .ip2(n8521), .op(n8529) );
  nand2_1 U8532 ( .ip1(n10036), .ip2(\ROUTEDATA/regData [79]), .op(n8527) );
  nand2_1 U8533 ( .ip1(n8523), .ip2(\ROUTEDATA/regData [159]), .op(n8526) );
  nand2_1 U8534 ( .ip1(n10028), .ip2(\ROUTEDATA/regData [47]), .op(n8525) );
  nand2_1 U8535 ( .ip1(n10044), .ip2(\ROUTEDATA/regData [111]), .op(n8524) );
  nand4_1 U8536 ( .ip1(n8527), .ip2(n8526), .ip3(n8525), .ip4(n8524), .op(
        n8528) );
  not_ab_or_c_or_d U8537 ( .ip1(n10040), .ip2(\ROUTEDATA/regData [95]), .ip3(
        n8529), .ip4(n8528), .op(n8533) );
  nand2_1 U8538 ( .ip1(n10032), .ip2(\ROUTEDATA/regData [63]), .op(n8532) );
  nand2_1 U8539 ( .ip1(n10023), .ip2(\ROUTEDATA/regData [31]), .op(n8531) );
  nand2_1 U8540 ( .ip1(\ROUTEDATA/regData [15]), .ip2(n10435), .op(n8530) );
  nand4_1 U8541 ( .ip1(n8533), .ip2(n8532), .ip3(n8531), .ip4(n8530), .op(
        n8535) );
  mux2_1 U8542 ( .ip1(m2DataIn[15]), .ip2(n8535), .s(n8534), .op(n4003) );
  inv_1 U8543 ( .ip(weight2AddrOffChip[3]), .op(n8536) );
  nand2_1 U8544 ( .ip1(n8536), .ip2(w2SramWeOffChip), .op(n8557) );
  nor2_1 U8545 ( .ip1(n8537), .ip2(n8557), .op(n8538) );
  mux2_1 U8546 ( .ip1(\WEIGHT_2/mem_w2[0][0] ), .ip2(weight2[0]), .s(n8538), 
        .op(n4002) );
  mux2_1 U8547 ( .ip1(\WEIGHT_2/mem_w2[0][1] ), .ip2(weight2[1]), .s(n8538), 
        .op(n4001) );
  mux2_1 U8548 ( .ip1(\WEIGHT_2/mem_w2[0][2] ), .ip2(weight2[2]), .s(n8538), 
        .op(n4000) );
  mux2_1 U8549 ( .ip1(\WEIGHT_2/mem_w2[0][3] ), .ip2(weight2[3]), .s(n8538), 
        .op(n3999) );
  mux2_1 U8550 ( .ip1(\WEIGHT_2/mem_w2[0][4] ), .ip2(weight2[4]), .s(n8538), 
        .op(n3998) );
  mux2_1 U8551 ( .ip1(\WEIGHT_2/mem_w2[0][5] ), .ip2(weight2[5]), .s(n8538), 
        .op(n3997) );
  mux2_1 U8552 ( .ip1(\WEIGHT_2/mem_w2[0][6] ), .ip2(weight2[6]), .s(n8538), 
        .op(n3996) );
  mux2_1 U8553 ( .ip1(\WEIGHT_2/mem_w2[0][7] ), .ip2(weight2[7]), .s(n8538), 
        .op(n3995) );
  mux2_1 U8554 ( .ip1(\WEIGHT_2/mem_w2[0][8] ), .ip2(weight2[8]), .s(n8538), 
        .op(n3994) );
  mux2_1 U8555 ( .ip1(\WEIGHT_2/mem_w2[0][9] ), .ip2(weight2[9]), .s(n8538), 
        .op(n3993) );
  mux2_1 U8556 ( .ip1(\WEIGHT_2/mem_w2[0][10] ), .ip2(weight2[10]), .s(n8538), 
        .op(n3992) );
  mux2_1 U8557 ( .ip1(\WEIGHT_2/mem_w2[0][11] ), .ip2(weight2[11]), .s(n8538), 
        .op(n3991) );
  mux2_1 U8558 ( .ip1(\WEIGHT_2/mem_w2[0][12] ), .ip2(weight2[12]), .s(n8538), 
        .op(n3990) );
  mux2_1 U8559 ( .ip1(\WEIGHT_2/mem_w2[0][13] ), .ip2(weight2[13]), .s(n8538), 
        .op(n3989) );
  mux2_1 U8560 ( .ip1(\WEIGHT_2/mem_w2[0][14] ), .ip2(weight2[14]), .s(n8538), 
        .op(n3988) );
  mux2_1 U8561 ( .ip1(\WEIGHT_2/mem_w2[0][15] ), .ip2(weight2[15]), .s(n8538), 
        .op(n3987) );
  nor2_1 U8562 ( .ip1(n8539), .ip2(n8557), .op(n8540) );
  mux2_1 U8563 ( .ip1(\WEIGHT_2/mem_w2[1][0] ), .ip2(weight2[0]), .s(n8540), 
        .op(n3986) );
  mux2_1 U8564 ( .ip1(\WEIGHT_2/mem_w2[1][1] ), .ip2(weight2[1]), .s(n8540), 
        .op(n3985) );
  mux2_1 U8565 ( .ip1(\WEIGHT_2/mem_w2[1][2] ), .ip2(weight2[2]), .s(n8540), 
        .op(n3984) );
  mux2_1 U8566 ( .ip1(\WEIGHT_2/mem_w2[1][3] ), .ip2(weight2[3]), .s(n8540), 
        .op(n3983) );
  mux2_1 U8567 ( .ip1(\WEIGHT_2/mem_w2[1][4] ), .ip2(weight2[4]), .s(n8540), 
        .op(n3982) );
  mux2_1 U8568 ( .ip1(\WEIGHT_2/mem_w2[1][5] ), .ip2(weight2[5]), .s(n8540), 
        .op(n3981) );
  mux2_1 U8569 ( .ip1(\WEIGHT_2/mem_w2[1][6] ), .ip2(weight2[6]), .s(n8540), 
        .op(n3980) );
  mux2_1 U8570 ( .ip1(\WEIGHT_2/mem_w2[1][7] ), .ip2(weight2[7]), .s(n8540), 
        .op(n3979) );
  mux2_1 U8571 ( .ip1(\WEIGHT_2/mem_w2[1][8] ), .ip2(weight2[8]), .s(n8540), 
        .op(n3978) );
  mux2_1 U8572 ( .ip1(\WEIGHT_2/mem_w2[1][9] ), .ip2(weight2[9]), .s(n8540), 
        .op(n3977) );
  mux2_1 U8573 ( .ip1(\WEIGHT_2/mem_w2[1][10] ), .ip2(weight2[10]), .s(n8540), 
        .op(n3976) );
  mux2_1 U8574 ( .ip1(\WEIGHT_2/mem_w2[1][11] ), .ip2(weight2[11]), .s(n8540), 
        .op(n3975) );
  mux2_1 U8575 ( .ip1(\WEIGHT_2/mem_w2[1][12] ), .ip2(weight2[12]), .s(n8540), 
        .op(n3974) );
  mux2_1 U8576 ( .ip1(\WEIGHT_2/mem_w2[1][13] ), .ip2(weight2[13]), .s(n8540), 
        .op(n3973) );
  mux2_1 U8577 ( .ip1(\WEIGHT_2/mem_w2[1][14] ), .ip2(weight2[14]), .s(n8540), 
        .op(n3972) );
  mux2_1 U8578 ( .ip1(\WEIGHT_2/mem_w2[1][15] ), .ip2(weight2[15]), .s(n8540), 
        .op(n3971) );
  inv_1 U8579 ( .ip(n8541), .op(n8542) );
  nor2_1 U8580 ( .ip1(n8542), .ip2(n8557), .op(n8543) );
  mux2_1 U8581 ( .ip1(\WEIGHT_2/mem_w2[2][0] ), .ip2(weight2[0]), .s(n8543), 
        .op(n3970) );
  mux2_1 U8582 ( .ip1(\WEIGHT_2/mem_w2[2][1] ), .ip2(weight2[1]), .s(n8543), 
        .op(n3969) );
  mux2_1 U8583 ( .ip1(\WEIGHT_2/mem_w2[2][2] ), .ip2(weight2[2]), .s(n8543), 
        .op(n3968) );
  mux2_1 U8584 ( .ip1(\WEIGHT_2/mem_w2[2][3] ), .ip2(weight2[3]), .s(n8543), 
        .op(n3967) );
  mux2_1 U8585 ( .ip1(\WEIGHT_2/mem_w2[2][4] ), .ip2(weight2[4]), .s(n8543), 
        .op(n3966) );
  mux2_1 U8586 ( .ip1(\WEIGHT_2/mem_w2[2][5] ), .ip2(weight2[5]), .s(n8543), 
        .op(n3965) );
  mux2_1 U8587 ( .ip1(\WEIGHT_2/mem_w2[2][6] ), .ip2(weight2[6]), .s(n8543), 
        .op(n3964) );
  mux2_1 U8588 ( .ip1(\WEIGHT_2/mem_w2[2][7] ), .ip2(weight2[7]), .s(n8543), 
        .op(n3963) );
  mux2_1 U8589 ( .ip1(\WEIGHT_2/mem_w2[2][8] ), .ip2(weight2[8]), .s(n8543), 
        .op(n3962) );
  mux2_1 U8590 ( .ip1(\WEIGHT_2/mem_w2[2][9] ), .ip2(weight2[9]), .s(n8543), 
        .op(n3961) );
  mux2_1 U8591 ( .ip1(\WEIGHT_2/mem_w2[2][10] ), .ip2(weight2[10]), .s(n8543), 
        .op(n3960) );
  mux2_1 U8592 ( .ip1(\WEIGHT_2/mem_w2[2][11] ), .ip2(weight2[11]), .s(n8543), 
        .op(n3959) );
  mux2_1 U8593 ( .ip1(\WEIGHT_2/mem_w2[2][12] ), .ip2(weight2[12]), .s(n8543), 
        .op(n3958) );
  mux2_1 U8594 ( .ip1(\WEIGHT_2/mem_w2[2][13] ), .ip2(weight2[13]), .s(n8543), 
        .op(n3957) );
  mux2_1 U8595 ( .ip1(\WEIGHT_2/mem_w2[2][14] ), .ip2(weight2[14]), .s(n8543), 
        .op(n3956) );
  mux2_1 U8596 ( .ip1(\WEIGHT_2/mem_w2[2][15] ), .ip2(weight2[15]), .s(n8543), 
        .op(n3955) );
  inv_1 U8597 ( .ip(n8544), .op(n8545) );
  nor2_1 U8598 ( .ip1(n8545), .ip2(n8557), .op(n8546) );
  mux2_1 U8599 ( .ip1(\WEIGHT_2/mem_w2[3][0] ), .ip2(weight2[0]), .s(n8546), 
        .op(n3954) );
  mux2_1 U8600 ( .ip1(\WEIGHT_2/mem_w2[3][1] ), .ip2(weight2[1]), .s(n8546), 
        .op(n3953) );
  mux2_1 U8601 ( .ip1(\WEIGHT_2/mem_w2[3][2] ), .ip2(weight2[2]), .s(n8546), 
        .op(n3952) );
  mux2_1 U8602 ( .ip1(\WEIGHT_2/mem_w2[3][3] ), .ip2(weight2[3]), .s(n8546), 
        .op(n3951) );
  mux2_1 U8603 ( .ip1(\WEIGHT_2/mem_w2[3][4] ), .ip2(weight2[4]), .s(n8546), 
        .op(n3950) );
  mux2_1 U8604 ( .ip1(\WEIGHT_2/mem_w2[3][5] ), .ip2(weight2[5]), .s(n8546), 
        .op(n3949) );
  mux2_1 U8605 ( .ip1(\WEIGHT_2/mem_w2[3][6] ), .ip2(weight2[6]), .s(n8546), 
        .op(n3948) );
  mux2_1 U8606 ( .ip1(\WEIGHT_2/mem_w2[3][7] ), .ip2(weight2[7]), .s(n8546), 
        .op(n3947) );
  mux2_1 U8607 ( .ip1(\WEIGHT_2/mem_w2[3][8] ), .ip2(weight2[8]), .s(n8546), 
        .op(n3946) );
  mux2_1 U8608 ( .ip1(\WEIGHT_2/mem_w2[3][9] ), .ip2(weight2[9]), .s(n8546), 
        .op(n3945) );
  mux2_1 U8609 ( .ip1(\WEIGHT_2/mem_w2[3][10] ), .ip2(weight2[10]), .s(n8546), 
        .op(n3944) );
  mux2_1 U8610 ( .ip1(\WEIGHT_2/mem_w2[3][11] ), .ip2(weight2[11]), .s(n8546), 
        .op(n3943) );
  mux2_1 U8611 ( .ip1(\WEIGHT_2/mem_w2[3][12] ), .ip2(weight2[12]), .s(n8546), 
        .op(n3942) );
  mux2_1 U8612 ( .ip1(\WEIGHT_2/mem_w2[3][13] ), .ip2(weight2[13]), .s(n8546), 
        .op(n3941) );
  mux2_1 U8613 ( .ip1(\WEIGHT_2/mem_w2[3][14] ), .ip2(weight2[14]), .s(n8546), 
        .op(n3940) );
  mux2_1 U8614 ( .ip1(\WEIGHT_2/mem_w2[3][15] ), .ip2(weight2[15]), .s(n8546), 
        .op(n3939) );
  inv_1 U8615 ( .ip(n8547), .op(n8548) );
  nor2_1 U8616 ( .ip1(n8548), .ip2(n8557), .op(n8549) );
  mux2_1 U8617 ( .ip1(\WEIGHT_2/mem_w2[4][0] ), .ip2(weight2[0]), .s(n8549), 
        .op(n3938) );
  mux2_1 U8618 ( .ip1(\WEIGHT_2/mem_w2[4][1] ), .ip2(weight2[1]), .s(n8549), 
        .op(n3937) );
  mux2_1 U8619 ( .ip1(\WEIGHT_2/mem_w2[4][2] ), .ip2(weight2[2]), .s(n8549), 
        .op(n3936) );
  mux2_1 U8620 ( .ip1(\WEIGHT_2/mem_w2[4][3] ), .ip2(weight2[3]), .s(n8549), 
        .op(n3935) );
  mux2_1 U8621 ( .ip1(\WEIGHT_2/mem_w2[4][4] ), .ip2(weight2[4]), .s(n8549), 
        .op(n3934) );
  mux2_1 U8622 ( .ip1(\WEIGHT_2/mem_w2[4][5] ), .ip2(weight2[5]), .s(n8549), 
        .op(n3933) );
  mux2_1 U8623 ( .ip1(\WEIGHT_2/mem_w2[4][6] ), .ip2(weight2[6]), .s(n8549), 
        .op(n3932) );
  mux2_1 U8624 ( .ip1(\WEIGHT_2/mem_w2[4][7] ), .ip2(weight2[7]), .s(n8549), 
        .op(n3931) );
  mux2_1 U8625 ( .ip1(\WEIGHT_2/mem_w2[4][8] ), .ip2(weight2[8]), .s(n8549), 
        .op(n3930) );
  mux2_1 U8626 ( .ip1(\WEIGHT_2/mem_w2[4][9] ), .ip2(weight2[9]), .s(n8549), 
        .op(n3929) );
  mux2_1 U8627 ( .ip1(\WEIGHT_2/mem_w2[4][10] ), .ip2(weight2[10]), .s(n8549), 
        .op(n3928) );
  mux2_1 U8628 ( .ip1(\WEIGHT_2/mem_w2[4][11] ), .ip2(weight2[11]), .s(n8549), 
        .op(n3927) );
  mux2_1 U8629 ( .ip1(\WEIGHT_2/mem_w2[4][12] ), .ip2(weight2[12]), .s(n8549), 
        .op(n3926) );
  mux2_1 U8630 ( .ip1(\WEIGHT_2/mem_w2[4][13] ), .ip2(weight2[13]), .s(n8549), 
        .op(n3925) );
  mux2_1 U8631 ( .ip1(\WEIGHT_2/mem_w2[4][14] ), .ip2(weight2[14]), .s(n8549), 
        .op(n3924) );
  mux2_1 U8632 ( .ip1(\WEIGHT_2/mem_w2[4][15] ), .ip2(weight2[15]), .s(n8549), 
        .op(n3923) );
  inv_1 U8633 ( .ip(n8550), .op(n8551) );
  nor2_1 U8634 ( .ip1(n8551), .ip2(n8557), .op(n8552) );
  mux2_1 U8635 ( .ip1(\WEIGHT_2/mem_w2[5][0] ), .ip2(weight2[0]), .s(n8552), 
        .op(n3922) );
  mux2_1 U8636 ( .ip1(\WEIGHT_2/mem_w2[5][1] ), .ip2(weight2[1]), .s(n8552), 
        .op(n3921) );
  mux2_1 U8637 ( .ip1(\WEIGHT_2/mem_w2[5][2] ), .ip2(weight2[2]), .s(n8552), 
        .op(n3920) );
  mux2_1 U8638 ( .ip1(\WEIGHT_2/mem_w2[5][3] ), .ip2(weight2[3]), .s(n8552), 
        .op(n3919) );
  mux2_1 U8639 ( .ip1(\WEIGHT_2/mem_w2[5][4] ), .ip2(weight2[4]), .s(n8552), 
        .op(n3918) );
  mux2_1 U8640 ( .ip1(\WEIGHT_2/mem_w2[5][5] ), .ip2(weight2[5]), .s(n8552), 
        .op(n3917) );
  mux2_1 U8641 ( .ip1(\WEIGHT_2/mem_w2[5][6] ), .ip2(weight2[6]), .s(n8552), 
        .op(n3916) );
  mux2_1 U8642 ( .ip1(\WEIGHT_2/mem_w2[5][7] ), .ip2(weight2[7]), .s(n8552), 
        .op(n3915) );
  mux2_1 U8643 ( .ip1(\WEIGHT_2/mem_w2[5][8] ), .ip2(weight2[8]), .s(n8552), 
        .op(n3914) );
  mux2_1 U8644 ( .ip1(\WEIGHT_2/mem_w2[5][9] ), .ip2(weight2[9]), .s(n8552), 
        .op(n3913) );
  mux2_1 U8645 ( .ip1(\WEIGHT_2/mem_w2[5][10] ), .ip2(weight2[10]), .s(n8552), 
        .op(n3912) );
  mux2_1 U8646 ( .ip1(\WEIGHT_2/mem_w2[5][11] ), .ip2(weight2[11]), .s(n8552), 
        .op(n3911) );
  mux2_1 U8647 ( .ip1(\WEIGHT_2/mem_w2[5][12] ), .ip2(weight2[12]), .s(n8552), 
        .op(n3910) );
  mux2_1 U8648 ( .ip1(\WEIGHT_2/mem_w2[5][13] ), .ip2(weight2[13]), .s(n8552), 
        .op(n3909) );
  mux2_1 U8649 ( .ip1(\WEIGHT_2/mem_w2[5][14] ), .ip2(weight2[14]), .s(n8552), 
        .op(n3908) );
  mux2_1 U8650 ( .ip1(\WEIGHT_2/mem_w2[5][15] ), .ip2(weight2[15]), .s(n8552), 
        .op(n3907) );
  inv_1 U8651 ( .ip(n8553), .op(n8554) );
  nor2_1 U8652 ( .ip1(n8554), .ip2(n8557), .op(n8555) );
  mux2_1 U8653 ( .ip1(\WEIGHT_2/mem_w2[6][0] ), .ip2(weight2[0]), .s(n8555), 
        .op(n3906) );
  mux2_1 U8654 ( .ip1(\WEIGHT_2/mem_w2[6][1] ), .ip2(weight2[1]), .s(n8555), 
        .op(n3905) );
  mux2_1 U8655 ( .ip1(\WEIGHT_2/mem_w2[6][2] ), .ip2(weight2[2]), .s(n8555), 
        .op(n3904) );
  mux2_1 U8656 ( .ip1(\WEIGHT_2/mem_w2[6][3] ), .ip2(weight2[3]), .s(n8555), 
        .op(n3903) );
  mux2_1 U8657 ( .ip1(\WEIGHT_2/mem_w2[6][4] ), .ip2(weight2[4]), .s(n8555), 
        .op(n3902) );
  mux2_1 U8658 ( .ip1(\WEIGHT_2/mem_w2[6][5] ), .ip2(weight2[5]), .s(n8555), 
        .op(n3901) );
  mux2_1 U8659 ( .ip1(\WEIGHT_2/mem_w2[6][6] ), .ip2(weight2[6]), .s(n8555), 
        .op(n3900) );
  mux2_1 U8660 ( .ip1(\WEIGHT_2/mem_w2[6][7] ), .ip2(weight2[7]), .s(n8555), 
        .op(n3899) );
  mux2_1 U8661 ( .ip1(\WEIGHT_2/mem_w2[6][8] ), .ip2(weight2[8]), .s(n8555), 
        .op(n3898) );
  mux2_1 U8662 ( .ip1(\WEIGHT_2/mem_w2[6][9] ), .ip2(weight2[9]), .s(n8555), 
        .op(n3897) );
  mux2_1 U8663 ( .ip1(\WEIGHT_2/mem_w2[6][10] ), .ip2(weight2[10]), .s(n8555), 
        .op(n3896) );
  mux2_1 U8664 ( .ip1(\WEIGHT_2/mem_w2[6][11] ), .ip2(weight2[11]), .s(n8555), 
        .op(n3895) );
  mux2_1 U8665 ( .ip1(\WEIGHT_2/mem_w2[6][12] ), .ip2(weight2[12]), .s(n8555), 
        .op(n3894) );
  mux2_1 U8666 ( .ip1(\WEIGHT_2/mem_w2[6][13] ), .ip2(weight2[13]), .s(n8555), 
        .op(n3893) );
  mux2_1 U8667 ( .ip1(\WEIGHT_2/mem_w2[6][14] ), .ip2(weight2[14]), .s(n8555), 
        .op(n3892) );
  mux2_1 U8668 ( .ip1(\WEIGHT_2/mem_w2[6][15] ), .ip2(weight2[15]), .s(n8555), 
        .op(n3891) );
  inv_1 U8669 ( .ip(n8556), .op(n8558) );
  nor2_1 U8670 ( .ip1(n8558), .ip2(n8557), .op(n8559) );
  mux2_1 U8671 ( .ip1(\WEIGHT_2/mem_w2[7][0] ), .ip2(weight2[0]), .s(n8559), 
        .op(n3890) );
  mux2_1 U8672 ( .ip1(\WEIGHT_2/mem_w2[7][1] ), .ip2(weight2[1]), .s(n8559), 
        .op(n3889) );
  mux2_1 U8673 ( .ip1(\WEIGHT_2/mem_w2[7][2] ), .ip2(weight2[2]), .s(n8559), 
        .op(n3888) );
  mux2_1 U8674 ( .ip1(\WEIGHT_2/mem_w2[7][3] ), .ip2(weight2[3]), .s(n8559), 
        .op(n3887) );
  mux2_1 U8675 ( .ip1(\WEIGHT_2/mem_w2[7][4] ), .ip2(weight2[4]), .s(n8559), 
        .op(n3886) );
  mux2_1 U8676 ( .ip1(\WEIGHT_2/mem_w2[7][5] ), .ip2(weight2[5]), .s(n8559), 
        .op(n3885) );
  mux2_1 U8677 ( .ip1(\WEIGHT_2/mem_w2[7][6] ), .ip2(weight2[6]), .s(n8559), 
        .op(n3884) );
  mux2_1 U8678 ( .ip1(\WEIGHT_2/mem_w2[7][7] ), .ip2(weight2[7]), .s(n8559), 
        .op(n3883) );
  mux2_1 U8679 ( .ip1(\WEIGHT_2/mem_w2[7][8] ), .ip2(weight2[8]), .s(n8559), 
        .op(n3882) );
  mux2_1 U8680 ( .ip1(\WEIGHT_2/mem_w2[7][9] ), .ip2(weight2[9]), .s(n8559), 
        .op(n3881) );
  mux2_1 U8681 ( .ip1(\WEIGHT_2/mem_w2[7][10] ), .ip2(weight2[10]), .s(n8559), 
        .op(n3880) );
  mux2_1 U8682 ( .ip1(\WEIGHT_2/mem_w2[7][11] ), .ip2(weight2[11]), .s(n8559), 
        .op(n3879) );
  mux2_1 U8683 ( .ip1(\WEIGHT_2/mem_w2[7][12] ), .ip2(weight2[12]), .s(n8559), 
        .op(n3878) );
  mux2_1 U8684 ( .ip1(\WEIGHT_2/mem_w2[7][13] ), .ip2(weight2[13]), .s(n8559), 
        .op(n3877) );
  mux2_1 U8685 ( .ip1(\WEIGHT_2/mem_w2[7][14] ), .ip2(weight2[14]), .s(n8559), 
        .op(n3876) );
  mux2_1 U8686 ( .ip1(\WEIGHT_2/mem_w2[7][15] ), .ip2(weight2[15]), .s(n8559), 
        .op(n3875) );
  nand3_1 U8687 ( .ip1(w2SramWeOffChip), .ip2(n8560), .ip3(
        weight2AddrOffChip[3]), .op(n8561) );
  mux2_1 U8688 ( .ip1(weight2[0]), .ip2(\WEIGHT_2/mem_w2[8][0] ), .s(n8561), 
        .op(n3874) );
  mux2_1 U8689 ( .ip1(weight2[1]), .ip2(\WEIGHT_2/mem_w2[8][1] ), .s(n8561), 
        .op(n3873) );
  mux2_1 U8690 ( .ip1(weight2[2]), .ip2(\WEIGHT_2/mem_w2[8][2] ), .s(n8561), 
        .op(n3872) );
  mux2_1 U8691 ( .ip1(weight2[3]), .ip2(\WEIGHT_2/mem_w2[8][3] ), .s(n8561), 
        .op(n3871) );
  mux2_1 U8692 ( .ip1(weight2[4]), .ip2(\WEIGHT_2/mem_w2[8][4] ), .s(n8561), 
        .op(n3870) );
  mux2_1 U8693 ( .ip1(weight2[5]), .ip2(\WEIGHT_2/mem_w2[8][5] ), .s(n8561), 
        .op(n3869) );
  mux2_1 U8694 ( .ip1(weight2[6]), .ip2(\WEIGHT_2/mem_w2[8][6] ), .s(n8561), 
        .op(n3868) );
  mux2_1 U8695 ( .ip1(weight2[7]), .ip2(\WEIGHT_2/mem_w2[8][7] ), .s(n8561), 
        .op(n3867) );
  mux2_1 U8696 ( .ip1(weight2[8]), .ip2(\WEIGHT_2/mem_w2[8][8] ), .s(n8561), 
        .op(n3866) );
  mux2_1 U8697 ( .ip1(weight2[9]), .ip2(\WEIGHT_2/mem_w2[8][9] ), .s(n8561), 
        .op(n3865) );
  mux2_1 U8698 ( .ip1(weight2[10]), .ip2(\WEIGHT_2/mem_w2[8][10] ), .s(n8561), 
        .op(n3864) );
  mux2_1 U8699 ( .ip1(weight2[11]), .ip2(\WEIGHT_2/mem_w2[8][11] ), .s(n8561), 
        .op(n3863) );
  mux2_1 U8700 ( .ip1(weight2[12]), .ip2(\WEIGHT_2/mem_w2[8][12] ), .s(n8561), 
        .op(n3862) );
  mux2_1 U8701 ( .ip1(weight2[13]), .ip2(\WEIGHT_2/mem_w2[8][13] ), .s(n8561), 
        .op(n3861) );
  mux2_1 U8702 ( .ip1(weight2[14]), .ip2(\WEIGHT_2/mem_w2[8][14] ), .s(n8561), 
        .op(n3860) );
  mux2_1 U8703 ( .ip1(weight2[15]), .ip2(\WEIGHT_2/mem_w2[8][15] ), .s(n8561), 
        .op(n3859) );
  nand3_1 U8704 ( .ip1(w2SramWeOffChip), .ip2(n8562), .ip3(
        weight2AddrOffChip[3]), .op(n8563) );
  mux2_1 U8705 ( .ip1(weight2[0]), .ip2(\WEIGHT_2/mem_w2[9][0] ), .s(n8563), 
        .op(n3858) );
  mux2_1 U8706 ( .ip1(weight2[1]), .ip2(\WEIGHT_2/mem_w2[9][1] ), .s(n8563), 
        .op(n3857) );
  mux2_1 U8707 ( .ip1(weight2[2]), .ip2(\WEIGHT_2/mem_w2[9][2] ), .s(n8563), 
        .op(n3856) );
  mux2_1 U8708 ( .ip1(weight2[3]), .ip2(\WEIGHT_2/mem_w2[9][3] ), .s(n8563), 
        .op(n3855) );
  mux2_1 U8709 ( .ip1(weight2[4]), .ip2(\WEIGHT_2/mem_w2[9][4] ), .s(n8563), 
        .op(n3854) );
  mux2_1 U8710 ( .ip1(weight2[5]), .ip2(\WEIGHT_2/mem_w2[9][5] ), .s(n8563), 
        .op(n3853) );
  mux2_1 U8711 ( .ip1(weight2[6]), .ip2(\WEIGHT_2/mem_w2[9][6] ), .s(n8563), 
        .op(n3852) );
  mux2_1 U8712 ( .ip1(weight2[7]), .ip2(\WEIGHT_2/mem_w2[9][7] ), .s(n8563), 
        .op(n3851) );
  mux2_1 U8713 ( .ip1(weight2[8]), .ip2(\WEIGHT_2/mem_w2[9][8] ), .s(n8563), 
        .op(n3850) );
  mux2_1 U8714 ( .ip1(weight2[9]), .ip2(\WEIGHT_2/mem_w2[9][9] ), .s(n8563), 
        .op(n3849) );
  mux2_1 U8715 ( .ip1(weight2[10]), .ip2(\WEIGHT_2/mem_w2[9][10] ), .s(n8563), 
        .op(n3848) );
  mux2_1 U8716 ( .ip1(weight2[11]), .ip2(\WEIGHT_2/mem_w2[9][11] ), .s(n8563), 
        .op(n3847) );
  mux2_1 U8717 ( .ip1(weight2[12]), .ip2(\WEIGHT_2/mem_w2[9][12] ), .s(n8563), 
        .op(n3846) );
  mux2_1 U8718 ( .ip1(weight2[13]), .ip2(\WEIGHT_2/mem_w2[9][13] ), .s(n8563), 
        .op(n3845) );
  mux2_1 U8719 ( .ip1(weight2[14]), .ip2(\WEIGHT_2/mem_w2[9][14] ), .s(n8563), 
        .op(n3844) );
  mux2_1 U8720 ( .ip1(weight2[15]), .ip2(\WEIGHT_2/mem_w2[9][15] ), .s(n8563), 
        .op(n3843) );
  inv_1 U8721 ( .ip(n8564), .op(n8590) );
  nand2_1 U8722 ( .ip1(n8566), .ip2(n8565), .op(n8602) );
  nor2_1 U8723 ( .ip1(n8591), .ip2(n8567), .op(n8605) );
  or2_1 U8724 ( .ip1(n8602), .ip2(n8605), .op(n8568) );
  nand2_1 U8725 ( .ip1(n8569), .ip2(n8568), .op(n8642) );
  nand3_1 U8726 ( .ip1(n8642), .ip2(n8620), .ip3(n8570), .op(n8589) );
  nor3_1 U8727 ( .ip1(n8584), .ip2(n8581), .ip3(n8571), .op(n8573) );
  nor2_1 U8728 ( .ip1(n8573), .ip2(n8572), .op(n8630) );
  nor2_1 U8729 ( .ip1(n8630), .ip2(n8574), .op(n8611) );
  nand2_1 U8730 ( .ip1(n8585), .ip2(n8575), .op(n8626) );
  nand2_1 U8731 ( .ip1(n8576), .ip2(n8634), .op(n8577) );
  nand4_1 U8732 ( .ip1(n8626), .ip2(n8579), .ip3(n8578), .ip4(n8577), .op(
        n8580) );
  not_ab_or_c_or_d U8733 ( .ip1(n8583), .ip2(n8582), .ip3(n8581), .ip4(n8580), 
        .op(n8587) );
  nand2_1 U8734 ( .ip1(n8585), .ip2(n8584), .op(n8624) );
  nand4_1 U8735 ( .ip1(n8611), .ip2(n8587), .ip3(n8586), .ip4(n8624), .op(
        n8588) );
  not_ab_or_c_or_d U8736 ( .ip1(n8590), .ip2(n8631), .ip3(n8589), .ip4(n8588), 
        .op(n8596) );
  nor3_1 U8737 ( .ip1(n8593), .ip2(n8592), .ip3(n8591), .op(n8595) );
  not_ab_or_c_or_d U8738 ( .ip1(n8597), .ip2(n8596), .ip3(n8595), .ip4(n8594), 
        .op(n3842) );
  inv_1 U8739 ( .ip(n8598), .op(n8615) );
  ab_or_c_or_d U8740 ( .ip1(n8601), .ip2(n8600), .ip3(n8599), .ip4(n8616), 
        .op(n8619) );
  inv_1 U8741 ( .ip(n8602), .op(n8606) );
  inv_1 U8742 ( .ip(n8637), .op(n8603) );
  not_ab_or_c_or_d U8743 ( .ip1(n8606), .ip2(n8605), .ip3(n8604), .ip4(n8603), 
        .op(n8610) );
  nand2_1 U8744 ( .ip1(n8624), .ip2(n8623), .op(n8627) );
  nor3_1 U8745 ( .ip1(n8627), .ip2(n8608), .ip3(n8607), .op(n8609) );
  nand4_1 U8746 ( .ip1(n8611), .ip2(n8619), .ip3(n8610), .ip4(n8609), .op(
        n8612) );
  or4_1 U8747 ( .ip1(n8615), .ip2(n8614), .ip3(n8613), .ip4(n8612), .op(n3841)
         );
  or2_1 U8748 ( .ip1(n8617), .ip2(n8616), .op(n8618) );
  nand4_1 U8749 ( .ip1(n8621), .ip2(n8620), .ip3(n8619), .ip4(n8618), .op(
        n8644) );
  nor4_1 U8750 ( .ip1(n8633), .ip2(n8622), .ip3(n8630), .ip4(n8644), .op(n8625) );
  nand3_1 U8751 ( .ip1(n8625), .ip2(n8624), .ip3(n8623), .op(n3838) );
  inv_1 U8752 ( .ip(n8626), .op(n8629) );
  nor3_1 U8753 ( .ip1(n8629), .ip2(n8628), .ip3(n8627), .op(n8638) );
  nor2_1 U8754 ( .ip1(n8631), .ip2(n8630), .op(n8641) );
  nand2_1 U8755 ( .ip1(n8638), .ip2(n8641), .op(n3837) );
  not_ab_or_c_or_d U8756 ( .ip1(n8635), .ip2(n8634), .ip3(n8633), .ip4(n8632), 
        .op(n8636) );
  nand3_1 U8757 ( .ip1(n8638), .ip2(n8637), .ip3(n8636), .op(n3836) );
  nand4_1 U8758 ( .ip1(n8642), .ip2(n8641), .ip3(n8640), .ip4(n8639), .op(
        n8643) );
  nor3_1 U8759 ( .ip1(n3836), .ip2(n8644), .ip3(n8643), .op(n3835) );
  inv_1 U8760 ( .ip(q_w2[5]), .op(n9703) );
  nor2_1 U8761 ( .ip1(n9335), .ip2(n9703), .op(n8645) );
  or2_1 U8762 ( .ip1(q_w2[2]), .ip2(n8645), .op(n8647) );
  or2_1 U8763 ( .ip1(m2DataIn[3]), .ip2(n8645), .op(n8646) );
  nand2_1 U8764 ( .ip1(n8647), .ip2(n8646), .op(n8682) );
  inv_1 U8765 ( .ip(m2DataIn[5]), .op(n9702) );
  inv_1 U8766 ( .ip(q_w2[0]), .op(n9141) );
  nor3_1 U8767 ( .ip1(n8682), .ip2(n9702), .ip3(n9141), .op(n8648) );
  inv_1 U8768 ( .ip(q_w2[2]), .op(n9499) );
  nor4_1 U8769 ( .ip1(n9530), .ip2(n9335), .ip3(n9499), .ip4(n9703), .op(n8683) );
  or2_1 U8770 ( .ip1(n8648), .ip2(n8683), .op(n8677) );
  nand2_1 U8771 ( .ip1(m2DataIn[2]), .ip2(q_w2[4]), .op(n8649) );
  inv_1 U8772 ( .ip(m2DataIn[2]), .op(n9500) );
  inv_1 U8773 ( .ip(q_w2[4]), .op(n9638) );
  nor4_1 U8774 ( .ip1(n9500), .ip2(n9417), .ip3(n9638), .ip4(n9703), .op(n8759) );
  or2_1 U8775 ( .ip1(n8649), .ip2(n8759), .op(n8652) );
  nand2_1 U8776 ( .ip1(m2DataIn[1]), .ip2(q_w2[5]), .op(n8650) );
  or2_1 U8777 ( .ip1(n8650), .ip2(n8759), .op(n8651) );
  nand2_1 U8778 ( .ip1(n8652), .ip2(n8651), .op(n8676) );
  inv_1 U8779 ( .ip(q_w2[6]), .op(n9732) );
  nor2_1 U8780 ( .ip1(n9335), .ip2(n9732), .op(n8854) );
  inv_1 U8781 ( .ip(q_w2[1]), .op(n9334) );
  nor2_1 U8782 ( .ip1(n9702), .ip2(n9334), .op(n8669) );
  nor2_1 U8783 ( .ip1(n9467), .ip2(n9141), .op(n8668) );
  and3_1 U8784 ( .ip1(m2DataIn[1]), .ip2(q_w2[6]), .ip3(n8653), .op(n8850) );
  nor2_1 U8785 ( .ip1(n9417), .ip2(n9732), .op(n8654) );
  nor2_1 U8786 ( .ip1(n8654), .ip2(n8653), .op(n8655) );
  nor2_1 U8787 ( .ip1(n8850), .ip2(n8655), .op(n8776) );
  inv_1 U8788 ( .ip(m2DataIn[4]), .op(n9640) );
  nor2_1 U8789 ( .ip1(n9640), .ip2(n9499), .op(n8679) );
  inv_1 U8790 ( .ip(q_w2[3]), .op(n9372) );
  nor4_1 U8791 ( .ip1(n9500), .ip2(n9417), .ip3(n9372), .ip4(n9638), .op(n8674) );
  and2_1 U8792 ( .ip1(m2DataIn[3]), .ip2(n8674), .op(n8657) );
  or2_1 U8793 ( .ip1(n8679), .ip2(n8657), .op(n8659) );
  nor2_1 U8794 ( .ip1(n9530), .ip2(n9372), .op(n8656) );
  mux2_1 U8795 ( .ip1(n8656), .ip2(n9530), .s(n8674), .op(n8678) );
  or2_1 U8796 ( .ip1(n8678), .ip2(n8657), .op(n8658) );
  nand2_1 U8797 ( .ip1(n8659), .ip2(n8658), .op(n8772) );
  nand2_1 U8798 ( .ip1(m2DataIn[0]), .ip2(q_w2[7]), .op(n8948) );
  nor2_1 U8799 ( .ip1(n9335), .ip2(n9638), .op(n8689) );
  and3_1 U8800 ( .ip1(m2DataIn[3]), .ip2(q_w2[7]), .ip3(n8689), .op(n8762) );
  or2_1 U8801 ( .ip1(n8948), .ip2(n8762), .op(n8662) );
  nand2_1 U8802 ( .ip1(m2DataIn[3]), .ip2(q_w2[4]), .op(n8660) );
  or2_1 U8803 ( .ip1(n8660), .ip2(n8762), .op(n8661) );
  nand2_1 U8804 ( .ip1(n8662), .ip2(n8661), .op(n8761) );
  nor2_1 U8805 ( .ip1(n9500), .ip2(n9703), .op(n8763) );
  xnor2_1 U8806 ( .ip1(n8761), .ip2(n8763), .op(n8771) );
  and3_1 U8807 ( .ip1(m2DataIn[5]), .ip2(q_w2[3]), .ip3(n8679), .op(n8769) );
  nor2_1 U8808 ( .ip1(n9640), .ip2(n9372), .op(n8663) );
  or2_1 U8809 ( .ip1(q_w2[2]), .ip2(n8663), .op(n8665) );
  or2_1 U8810 ( .ip1(m2DataIn[5]), .ip2(n8663), .op(n8664) );
  nand2_1 U8811 ( .ip1(n8665), .ip2(n8664), .op(n8767) );
  nor2_1 U8812 ( .ip1(n8769), .ip2(n8767), .op(n8666) );
  nand2_1 U8813 ( .ip1(m2DataIn[7]), .ip2(q_w2[0]), .op(n8766) );
  xor2_1 U8814 ( .ip1(n8666), .ip2(n8766), .op(n8770) );
  inv_1 U8815 ( .ip(n8667), .op(n8775) );
  fulladder U8816 ( .a(n8854), .b(n8669), .ci(n8668), .co(n8758), .s(n8675) );
  nor2_1 U8817 ( .ip1(n9467), .ip2(n9334), .op(n8757) );
  nand2_1 U8818 ( .ip1(m2DataIn[1]), .ip2(q_w2[2]), .op(n8695) );
  nor3_1 U8819 ( .ip1(n9500), .ip2(n9372), .ip3(n8695), .op(n8691) );
  nor2_1 U8820 ( .ip1(n9500), .ip2(n9372), .op(n8670) );
  or2_1 U8821 ( .ip1(q_w2[4]), .ip2(n8670), .op(n8672) );
  or2_1 U8822 ( .ip1(m2DataIn[1]), .ip2(n8670), .op(n8671) );
  nand2_1 U8823 ( .ip1(n8672), .ip2(n8671), .op(n8673) );
  nor2_1 U8824 ( .ip1(n8674), .ip2(n8673), .op(n8681) );
  nor2_1 U8825 ( .ip1(n9640), .ip2(n9334), .op(n8680) );
  fulladder U8826 ( .a(n8677), .b(n8676), .ci(n8675), .co(n8653), .s(n8729) );
  xor2_1 U8827 ( .ip1(n8679), .ip2(n8678), .op(n8728) );
  nand2_1 U8828 ( .ip1(n8738), .ip2(n8737), .op(n8743) );
  fulladder U8829 ( .a(n8691), .b(n8681), .ci(n8680), .co(n8730), .s(n8727) );
  nor2_1 U8830 ( .ip1(n9530), .ip2(n9334), .op(n8688) );
  nor2_1 U8831 ( .ip1(n9640), .ip2(n9141), .op(n8687) );
  nor2_1 U8832 ( .ip1(n8683), .ip2(n8682), .op(n8685) );
  nor2_1 U8833 ( .ip1(n9702), .ip2(n9141), .op(n8684) );
  xor2_1 U8834 ( .ip1(n8685), .ip2(n8684), .op(n8725) );
  nand2_1 U8835 ( .ip1(m2DataIn[1]), .ip2(q_w2[1]), .op(n8703) );
  or3_1 U8836 ( .ip1(n9500), .ip2(n9141), .ip3(n8703), .op(n8700) );
  nand2_1 U8837 ( .ip1(m2DataIn[0]), .ip2(q_w2[3]), .op(n8699) );
  and2_1 U8838 ( .ip1(n8700), .ip2(n8699), .op(n8686) );
  nor3_1 U8839 ( .ip1(n8686), .ip2(n9334), .ip3(n9500), .op(n8713) );
  fulladder U8840 ( .a(n8689), .b(n8688), .ci(n8687), .co(n8726), .s(n8721) );
  nor3_1 U8841 ( .ip1(n9530), .ip2(n9141), .ip3(n8695), .op(n8720) );
  nand2_1 U8842 ( .ip1(m2DataIn[1]), .ip2(q_w2[3]), .op(n8690) );
  or2_1 U8843 ( .ip1(n8690), .ip2(n8691), .op(n8694) );
  nand2_1 U8844 ( .ip1(m2DataIn[2]), .ip2(q_w2[2]), .op(n8692) );
  or2_1 U8845 ( .ip1(n8692), .ip2(n8691), .op(n8693) );
  nand2_1 U8846 ( .ip1(n8694), .ip2(n8693), .op(n8719) );
  nand2_1 U8847 ( .ip1(n8713), .ip2(n8715), .op(n8718) );
  or2_1 U8848 ( .ip1(n8695), .ip2(n8720), .op(n8698) );
  nand2_1 U8849 ( .ip1(m2DataIn[3]), .ip2(q_w2[0]), .op(n8696) );
  or2_1 U8850 ( .ip1(n8696), .ip2(n8720), .op(n8697) );
  nand2_1 U8851 ( .ip1(n8698), .ip2(n8697), .op(n8707) );
  nor2_1 U8852 ( .ip1(n9500), .ip2(n9334), .op(n8702) );
  xor2_1 U8853 ( .ip1(n8700), .ip2(n8699), .op(n8701) );
  xor2_1 U8854 ( .ip1(n8702), .ip2(n8701), .op(n8709) );
  nand2_1 U8855 ( .ip1(n8707), .ip2(n8709), .op(n8712) );
  nor4_1 U8856 ( .ip1(m2DataIn[2]), .ip2(n9335), .ip3(n9141), .ip4(n8703), 
        .op(n8706) );
  nand2_1 U8857 ( .ip1(m2DataIn[2]), .ip2(q_w2[0]), .op(n8704) );
  not_ab_or_c_or_d U8858 ( .ip1(n8704), .ip2(n8703), .ip3(n9335), .ip4(n9499), 
        .op(n8705) );
  or2_1 U8859 ( .ip1(n8706), .ip2(n8705), .op(n8708) );
  nand2_1 U8860 ( .ip1(n8707), .ip2(n8708), .op(n8711) );
  nand2_1 U8861 ( .ip1(n8709), .ip2(n8708), .op(n8710) );
  nand3_1 U8862 ( .ip1(n8712), .ip2(n8711), .ip3(n8710), .op(n8714) );
  nand2_1 U8863 ( .ip1(n8713), .ip2(n8714), .op(n8717) );
  nand2_1 U8864 ( .ip1(n8715), .ip2(n8714), .op(n8716) );
  nand3_1 U8865 ( .ip1(n8718), .ip2(n8717), .ip3(n8716), .op(n8722) );
  nand2_1 U8866 ( .ip1(n8724), .ip2(n8722), .op(n8734) );
  fulladder U8867 ( .a(n8721), .b(n8720), .ci(n8719), .co(n8723), .s(n8715) );
  nand2_1 U8868 ( .ip1(n8722), .ip2(n8723), .op(n8733) );
  nand2_1 U8869 ( .ip1(n8724), .ip2(n8723), .op(n8732) );
  fulladder U8870 ( .a(n8727), .b(n8726), .ci(n8725), .co(n8736), .s(n8724) );
  fulladder U8871 ( .a(n8730), .b(n8729), .ci(n8728), .co(n8737), .s(n8735) );
  nand2_1 U8872 ( .ip1(n8736), .ip2(n8735), .op(n8731) );
  nand4_1 U8873 ( .ip1(n8734), .ip2(n8733), .ip3(n8732), .ip4(n8731), .op(
        n8741) );
  or2_1 U8874 ( .ip1(n8736), .ip2(n8735), .op(n8740) );
  or2_1 U8875 ( .ip1(n8738), .ip2(n8737), .op(n8739) );
  nand3_1 U8876 ( .ip1(n8741), .ip2(n8740), .ip3(n8739), .op(n8742) );
  nand2_1 U8877 ( .ip1(n8743), .ip2(n8742), .op(n8853) );
  nand2_1 U8878 ( .ip1(m2DataIn[4]), .ip2(q_w2[4]), .op(n8744) );
  nand2_1 U8879 ( .ip1(m2DataIn[5]), .ip2(q_w2[4]), .op(n8860) );
  nor3_1 U8880 ( .ip1(n9640), .ip2(n9372), .ip3(n8860), .op(n8866) );
  or2_1 U8881 ( .ip1(n8744), .ip2(n8866), .op(n8747) );
  nand2_1 U8882 ( .ip1(m2DataIn[5]), .ip2(q_w2[3]), .op(n8745) );
  or2_1 U8883 ( .ip1(n8745), .ip2(n8866), .op(n8746) );
  nand2_1 U8884 ( .ip1(n8747), .ip2(n8746), .op(n8865) );
  inv_1 U8885 ( .ip(m2DataIn[7]), .op(n9725) );
  nor2_1 U8886 ( .ip1(n9725), .ip2(n9334), .op(n8867) );
  xor2_1 U8887 ( .ip1(n8865), .ip2(n8867), .op(n8890) );
  nand2_1 U8888 ( .ip1(m2DataIn[0]), .ip2(q_w2[8]), .op(n8748) );
  nand2_1 U8889 ( .ip1(m2DataIn[3]), .ip2(q_w2[8]), .op(n8970) );
  nor3_1 U8890 ( .ip1(n9335), .ip2(n9703), .ip3(n8970), .op(n8875) );
  or2_1 U8891 ( .ip1(n8748), .ip2(n8875), .op(n8751) );
  nand2_1 U8892 ( .ip1(m2DataIn[3]), .ip2(q_w2[5]), .op(n8749) );
  or2_1 U8893 ( .ip1(n8749), .ip2(n8875), .op(n8750) );
  nand2_1 U8894 ( .ip1(n8751), .ip2(n8750), .op(n8874) );
  nor2_1 U8895 ( .ip1(n9817), .ip2(n9141), .op(n8876) );
  xor2_1 U8896 ( .ip1(n8874), .ip2(n8876), .op(n8889) );
  nand2_1 U8897 ( .ip1(m2DataIn[1]), .ip2(q_w2[7]), .op(n8870) );
  nand4_1 U8898 ( .ip1(m2DataIn[2]), .ip2(m2DataIn[1]), .ip3(q_w2[6]), .ip4(
        q_w2[7]), .op(n8887) );
  inv_1 U8899 ( .ip(n8887), .op(n8752) );
  or2_1 U8900 ( .ip1(n8870), .ip2(n8752), .op(n8755) );
  nand2_1 U8901 ( .ip1(m2DataIn[2]), .ip2(q_w2[6]), .op(n8753) );
  or2_1 U8902 ( .ip1(n8753), .ip2(n8752), .op(n8754) );
  nand2_1 U8903 ( .ip1(n8755), .ip2(n8754), .op(n8885) );
  mux2_1 U8904 ( .ip1(rdata[0]), .ip2(n8756), .s(n8885), .op(n8888) );
  fulladder U8905 ( .a(n8759), .b(n8758), .ci(n8757), .co(n8760), .s(n8774) );
  inv_1 U8906 ( .ip(n8760), .op(n8894) );
  or2_1 U8907 ( .ip1(n8761), .ip2(n8762), .op(n8765) );
  or2_1 U8908 ( .ip1(n8763), .ip2(n8762), .op(n8764) );
  nand2_1 U8909 ( .ip1(n8765), .ip2(n8764), .op(n8864) );
  nand2_1 U8910 ( .ip1(m2DataIn[6]), .ip2(q_w2[2]), .op(n8880) );
  nor2_1 U8911 ( .ip1(n8767), .ip2(n8766), .op(n8768) );
  nor2_1 U8912 ( .ip1(n8769), .ip2(n8768), .op(n8863) );
  fulladder U8913 ( .a(n8772), .b(n8771), .ci(n8770), .co(n8892), .s(n8667) );
  inv_1 U8914 ( .ip(n8773), .op(n8848) );
  fulladder U8915 ( .a(n8776), .b(n8775), .ci(n8774), .co(n8851), .s(n8738) );
  mux2_1 U8916 ( .ip1(n8777), .ip2(\SIGMOID/N64 ), .s(n9907), .op(n8831) );
  buf_1 U8917 ( .ip(n8831), .op(n8840) );
  or2_1 U8918 ( .ip1(\CNTRL/count_10_2Q [2]), .ip2(n8778), .op(n8780) );
  or2_1 U8919 ( .ip1(n8804), .ip2(n8778), .op(n8779) );
  nand2_1 U8920 ( .ip1(n8780), .ip2(n8779), .op(n8814) );
  or2_1 U8921 ( .ip1(n8804), .ip2(n8781), .op(n8783) );
  or2_1 U8922 ( .ip1(\CNTRL/count_10_2Q [1]), .ip2(n8781), .op(n8782) );
  nand2_1 U8923 ( .ip1(n8783), .ip2(n8782), .op(n8813) );
  nand2_1 U8924 ( .ip1(n8814), .ip2(n8813), .op(n8815) );
  nand2_1 U8925 ( .ip1(n8804), .ip2(\CNTRL/count_10_2Q [0]), .op(n8785) );
  nand2_1 U8926 ( .ip1(n8785), .ip2(n8784), .op(n8816) );
  nor2_1 U8927 ( .ip1(n8815), .ip2(n8816), .op(n12108) );
  or2_1 U8928 ( .ip1(n8804), .ip2(n8786), .op(n8788) );
  or2_1 U8929 ( .ip1(\CNTRL/count_10_2Q [3]), .ip2(n8786), .op(n8787) );
  nand2_1 U8930 ( .ip1(n8788), .ip2(n8787), .op(n12190) );
  nand2_1 U8931 ( .ip1(n12108), .ip2(n12190), .op(n8835) );
  nor2_1 U8932 ( .ip1(n8802), .ip2(n8789), .op(n8790) );
  or2_1 U8933 ( .ip1(\CNTRL/count_10Q [1]), .ip2(n8790), .op(n8792) );
  or2_1 U8934 ( .ip1(n8804), .ip2(n8790), .op(n8791) );
  nand2_1 U8935 ( .ip1(n8792), .ip2(n8791), .op(n12098) );
  nand2_1 U8936 ( .ip1(n8793), .ip2(\CNTRL/count_20Q [0]), .op(n8794) );
  nand2_1 U8937 ( .ip1(n9445), .ip2(n8794), .op(n8828) );
  nand2_1 U8938 ( .ip1(n12098), .ip2(n8828), .op(n8800) );
  nor2_1 U8939 ( .ip1(n8802), .ip2(n8795), .op(n8796) );
  or2_1 U8940 ( .ip1(\CNTRL/count_10Q [2]), .ip2(n8796), .op(n8798) );
  or2_1 U8941 ( .ip1(n8804), .ip2(n8796), .op(n8797) );
  nand2_1 U8942 ( .ip1(n8798), .ip2(n8797), .op(n8799) );
  inv_1 U8943 ( .ip(n8799), .op(n8821) );
  nor2_1 U8944 ( .ip1(n8800), .ip2(n8821), .op(n8834) );
  nor2_1 U8945 ( .ip1(n8802), .ip2(n8801), .op(n8803) );
  or2_1 U8946 ( .ip1(\CNTRL/count_10Q [0]), .ip2(n8803), .op(n8806) );
  or2_1 U8947 ( .ip1(n8804), .ip2(n8803), .op(n8805) );
  nand2_1 U8948 ( .ip1(n8806), .ip2(n8805), .op(n12109) );
  inv_1 U8949 ( .ip(n12109), .op(n10878) );
  nor2_1 U8950 ( .ip1(\CNTRL/count_10Q [3]), .ip2(n8810), .op(n8808) );
  not_ab_or_c_or_d U8951 ( .ip1(n8810), .ip2(n8809), .ip3(n8808), .ip4(n8807), 
        .op(n11565) );
  nand3_1 U8952 ( .ip1(n8834), .ip2(n12109), .ip3(n11996), .op(n8819) );
  nor2_1 U8953 ( .ip1(n8835), .ip2(n8819), .op(n9910) );
  mux2_1 U8954 ( .ip1(\ANSWER/mem[0][0][0] ), .ip2(n8840), .s(n9910), .op(
        n3834) );
  inv_1 U8955 ( .ip(n8816), .op(n8817) );
  nor2_1 U8956 ( .ip1(n8817), .ip2(n8815), .op(n12157) );
  nand2_1 U8957 ( .ip1(n12190), .ip2(n12157), .op(n8836) );
  nor2_1 U8958 ( .ip1(n8819), .ip2(n8836), .op(n9911) );
  mux2_1 U8959 ( .ip1(\ANSWER/mem[0][1][0] ), .ip2(n8840), .s(n9911), .op(
        n3833) );
  inv_1 U8960 ( .ip(n8814), .op(n8811) );
  nor3_1 U8961 ( .ip1(n8813), .ip2(n8811), .ip3(n8816), .op(n12147) );
  nand2_1 U8962 ( .ip1(n12190), .ip2(n12147), .op(n8837) );
  nor2_1 U8963 ( .ip1(n8819), .ip2(n8837), .op(n9912) );
  mux2_1 U8964 ( .ip1(\ANSWER/mem[0][2][0] ), .ip2(n8840), .s(n9912), .op(
        n3832) );
  nor3_1 U8965 ( .ip1(n8813), .ip2(n8817), .ip3(n8811), .op(n12137) );
  nand2_1 U8966 ( .ip1(n12190), .ip2(n12137), .op(n8838) );
  nor2_1 U8967 ( .ip1(n8819), .ip2(n8838), .op(n9913) );
  mux2_1 U8968 ( .ip1(\ANSWER/mem[0][3][0] ), .ip2(n8840), .s(n9913), .op(
        n3831) );
  inv_1 U8969 ( .ip(n8813), .op(n8812) );
  nor3_1 U8970 ( .ip1(n8814), .ip2(n8812), .ip3(n8816), .op(n12176) );
  nand2_1 U8971 ( .ip1(n12190), .ip2(n12176), .op(n8839) );
  nor2_1 U8972 ( .ip1(n8819), .ip2(n8839), .op(n9914) );
  mux2_1 U8973 ( .ip1(\ANSWER/mem[0][4][0] ), .ip2(n8840), .s(n9914), .op(
        n3830) );
  nor3_1 U8974 ( .ip1(n8814), .ip2(n8817), .ip3(n8812), .op(n12127) );
  nand2_1 U8975 ( .ip1(n12190), .ip2(n12127), .op(n8841) );
  nor2_1 U8976 ( .ip1(n8819), .ip2(n8841), .op(n9915) );
  mux2_1 U8977 ( .ip1(\ANSWER/mem[0][5][0] ), .ip2(n8840), .s(n9915), .op(
        n3829) );
  nor3_1 U8978 ( .ip1(n8814), .ip2(n8813), .ip3(n8816), .op(n12168) );
  nand2_1 U8979 ( .ip1(n12190), .ip2(n12168), .op(n8842) );
  nor2_1 U8980 ( .ip1(n8819), .ip2(n8842), .op(n9916) );
  mux2_1 U8981 ( .ip1(\ANSWER/mem[0][6][0] ), .ip2(n8840), .s(n9916), .op(
        n3828) );
  nor3_1 U8982 ( .ip1(n8814), .ip2(n8813), .ip3(n8817), .op(n12186) );
  nand2_1 U8983 ( .ip1(n12190), .ip2(n12186), .op(n8843) );
  nor2_1 U8984 ( .ip1(n8819), .ip2(n8843), .op(n9917) );
  mux2_1 U8985 ( .ip1(\ANSWER/mem[0][7][0] ), .ip2(n8840), .s(n9917), .op(
        n3827) );
  inv_1 U8986 ( .ip(n8815), .op(n8818) );
  nor2_1 U8987 ( .ip1(n12190), .ip2(n8816), .op(n12201) );
  nand2_1 U8988 ( .ip1(n8818), .ip2(n12201), .op(n8844) );
  nor2_1 U8989 ( .ip1(n8819), .ip2(n8844), .op(n9918) );
  mux2_1 U8990 ( .ip1(\ANSWER/mem[0][8][0] ), .ip2(n8840), .s(n9918), .op(
        n3826) );
  nor2_1 U8991 ( .ip1(n8817), .ip2(n12190), .op(n12215) );
  nand2_1 U8992 ( .ip1(n8818), .ip2(n12215), .op(n8846) );
  nor2_1 U8993 ( .ip1(n8819), .ip2(n8846), .op(n9919) );
  mux2_1 U8994 ( .ip1(\ANSWER/mem[0][9][0] ), .ip2(n8840), .s(n9919), .op(
        n3825) );
  inv_1 U8995 ( .ip(n12109), .op(n8833) );
  nand3_1 U8996 ( .ip1(n8834), .ip2(n11996), .ip3(n8833), .op(n8820) );
  nor2_1 U8997 ( .ip1(n8835), .ip2(n8820), .op(n9920) );
  mux2_1 U8998 ( .ip1(\ANSWER/mem[1][0][0] ), .ip2(n8840), .s(n9920), .op(
        n3824) );
  nor2_1 U8999 ( .ip1(n8836), .ip2(n8820), .op(n9921) );
  mux2_1 U9000 ( .ip1(\ANSWER/mem[1][1][0] ), .ip2(n8840), .s(n9921), .op(
        n3823) );
  nor2_1 U9001 ( .ip1(n8837), .ip2(n8820), .op(n9922) );
  mux2_1 U9002 ( .ip1(\ANSWER/mem[1][2][0] ), .ip2(n8831), .s(n9922), .op(
        n3822) );
  nor2_1 U9003 ( .ip1(n8838), .ip2(n8820), .op(n9923) );
  mux2_1 U9004 ( .ip1(\ANSWER/mem[1][3][0] ), .ip2(n8831), .s(n9923), .op(
        n3821) );
  nor2_1 U9005 ( .ip1(n8839), .ip2(n8820), .op(n9924) );
  mux2_1 U9006 ( .ip1(\ANSWER/mem[1][4][0] ), .ip2(n8831), .s(n9924), .op(
        n3820) );
  nor2_1 U9007 ( .ip1(n8841), .ip2(n8820), .op(n9925) );
  mux2_1 U9008 ( .ip1(\ANSWER/mem[1][5][0] ), .ip2(n8831), .s(n9925), .op(
        n3819) );
  nor2_1 U9009 ( .ip1(n8842), .ip2(n8820), .op(n9926) );
  mux2_1 U9010 ( .ip1(\ANSWER/mem[1][6][0] ), .ip2(n8831), .s(n9926), .op(
        n3818) );
  nor2_1 U9011 ( .ip1(n8843), .ip2(n8820), .op(n9927) );
  mux2_1 U9012 ( .ip1(\ANSWER/mem[1][7][0] ), .ip2(n8831), .s(n9927), .op(
        n3817) );
  nor2_1 U9013 ( .ip1(n8844), .ip2(n8820), .op(n9928) );
  mux2_1 U9014 ( .ip1(\ANSWER/mem[1][8][0] ), .ip2(n8831), .s(n9928), .op(
        n3816) );
  nor2_1 U9015 ( .ip1(n8846), .ip2(n8820), .op(n9929) );
  mux2_1 U9016 ( .ip1(\ANSWER/mem[1][9][0] ), .ip2(n8840), .s(n9929), .op(
        n3815) );
  inv_1 U9017 ( .ip(n11996), .op(n11336) );
  nor2_1 U9018 ( .ip1(n10878), .ip2(n11336), .op(n8826) );
  inv_1 U9019 ( .ip(n12098), .op(n11224) );
  nand4_1 U9020 ( .ip1(n8799), .ip2(n8826), .ip3(n8828), .ip4(n11224), .op(
        n8822) );
  nor2_1 U9021 ( .ip1(n8835), .ip2(n8822), .op(n9930) );
  mux2_1 U9022 ( .ip1(\ANSWER/mem[2][0][0] ), .ip2(n8840), .s(n9930), .op(
        n3814) );
  buf_1 U9023 ( .ip(n8831), .op(n8847) );
  nor2_1 U9024 ( .ip1(n8836), .ip2(n8822), .op(n9931) );
  mux2_1 U9025 ( .ip1(\ANSWER/mem[2][1][0] ), .ip2(n8847), .s(n9931), .op(
        n3813) );
  nor2_1 U9026 ( .ip1(n8837), .ip2(n8822), .op(n9932) );
  mux2_1 U9027 ( .ip1(\ANSWER/mem[2][2][0] ), .ip2(n8831), .s(n9932), .op(
        n3812) );
  nor2_1 U9028 ( .ip1(n8838), .ip2(n8822), .op(n9933) );
  mux2_1 U9029 ( .ip1(\ANSWER/mem[2][3][0] ), .ip2(n8831), .s(n9933), .op(
        n3811) );
  nor2_1 U9030 ( .ip1(n8839), .ip2(n8822), .op(n9934) );
  mux2_1 U9031 ( .ip1(\ANSWER/mem[2][4][0] ), .ip2(n8831), .s(n9934), .op(
        n3810) );
  nor2_1 U9032 ( .ip1(n8841), .ip2(n8822), .op(n9935) );
  mux2_1 U9033 ( .ip1(\ANSWER/mem[2][5][0] ), .ip2(n8831), .s(n9935), .op(
        n3809) );
  nor2_1 U9034 ( .ip1(n8842), .ip2(n8822), .op(n9936) );
  mux2_1 U9035 ( .ip1(\ANSWER/mem[2][6][0] ), .ip2(n8831), .s(n9936), .op(
        n3808) );
  nor2_1 U9036 ( .ip1(n8843), .ip2(n8822), .op(n9937) );
  mux2_1 U9037 ( .ip1(\ANSWER/mem[2][7][0] ), .ip2(n8831), .s(n9937), .op(
        n3807) );
  nor2_1 U9038 ( .ip1(n8844), .ip2(n8822), .op(n9938) );
  mux2_1 U9039 ( .ip1(\ANSWER/mem[2][8][0] ), .ip2(n8831), .s(n9938), .op(
        n3806) );
  nor2_1 U9040 ( .ip1(n8846), .ip2(n8822), .op(n9939) );
  mux2_1 U9041 ( .ip1(\ANSWER/mem[2][9][0] ), .ip2(n8831), .s(n9939), .op(
        n3805) );
  nor2_1 U9042 ( .ip1(n12109), .ip2(n11336), .op(n8829) );
  inv_1 U9043 ( .ip(n12098), .op(n11008) );
  nand4_1 U9044 ( .ip1(n8799), .ip2(n8829), .ip3(n8828), .ip4(n11008), .op(
        n8823) );
  nor2_1 U9045 ( .ip1(n8835), .ip2(n8823), .op(n9940) );
  mux2_1 U9046 ( .ip1(\ANSWER/mem[3][0][0] ), .ip2(n8831), .s(n9940), .op(
        n3804) );
  nor2_1 U9047 ( .ip1(n8836), .ip2(n8823), .op(n9941) );
  mux2_1 U9048 ( .ip1(\ANSWER/mem[3][1][0] ), .ip2(n8831), .s(n9941), .op(
        n3803) );
  nor2_1 U9049 ( .ip1(n8837), .ip2(n8823), .op(n9942) );
  mux2_1 U9050 ( .ip1(\ANSWER/mem[3][2][0] ), .ip2(n8831), .s(n9942), .op(
        n3802) );
  nor2_1 U9051 ( .ip1(n8838), .ip2(n8823), .op(n9943) );
  mux2_1 U9052 ( .ip1(\ANSWER/mem[3][3][0] ), .ip2(n8831), .s(n9943), .op(
        n3801) );
  nor2_1 U9053 ( .ip1(n8839), .ip2(n8823), .op(n9944) );
  mux2_1 U9054 ( .ip1(\ANSWER/mem[3][4][0] ), .ip2(n8831), .s(n9944), .op(
        n3800) );
  nor2_1 U9055 ( .ip1(n8841), .ip2(n8823), .op(n9945) );
  mux2_1 U9056 ( .ip1(\ANSWER/mem[3][5][0] ), .ip2(n8831), .s(n9945), .op(
        n3799) );
  nor2_1 U9057 ( .ip1(n8842), .ip2(n8823), .op(n9946) );
  mux2_1 U9058 ( .ip1(\ANSWER/mem[3][6][0] ), .ip2(n8847), .s(n9946), .op(
        n3798) );
  nor2_1 U9059 ( .ip1(n8843), .ip2(n8823), .op(n9947) );
  mux2_1 U9060 ( .ip1(\ANSWER/mem[3][7][0] ), .ip2(n8840), .s(n9947), .op(
        n3797) );
  nor2_1 U9061 ( .ip1(n8844), .ip2(n8823), .op(n9948) );
  mux2_1 U9062 ( .ip1(\ANSWER/mem[3][8][0] ), .ip2(n8831), .s(n9948), .op(
        n3796) );
  nor2_1 U9063 ( .ip1(n8846), .ip2(n8823), .op(n9949) );
  mux2_1 U9064 ( .ip1(\ANSWER/mem[3][9][0] ), .ip2(n8831), .s(n9949), .op(
        n3795) );
  inv_1 U9065 ( .ip(n8799), .op(n11979) );
  buf_1 U9066 ( .ip(n11979), .op(n11937) );
  nand4_1 U9067 ( .ip1(n12098), .ip2(n8826), .ip3(n8828), .ip4(n11937), .op(
        n8824) );
  nor2_1 U9068 ( .ip1(n8835), .ip2(n8824), .op(n9950) );
  mux2_1 U9069 ( .ip1(\ANSWER/mem[4][0][0] ), .ip2(n8831), .s(n9950), .op(
        n3794) );
  nor2_1 U9070 ( .ip1(n8836), .ip2(n8824), .op(n9951) );
  mux2_1 U9071 ( .ip1(\ANSWER/mem[4][1][0] ), .ip2(n8831), .s(n9951), .op(
        n3793) );
  nor2_1 U9072 ( .ip1(n8837), .ip2(n8824), .op(n9952) );
  mux2_1 U9073 ( .ip1(\ANSWER/mem[4][2][0] ), .ip2(n8831), .s(n9952), .op(
        n3792) );
  nor2_1 U9074 ( .ip1(n8838), .ip2(n8824), .op(n9953) );
  mux2_1 U9075 ( .ip1(\ANSWER/mem[4][3][0] ), .ip2(n8847), .s(n9953), .op(
        n3791) );
  nor2_1 U9076 ( .ip1(n8839), .ip2(n8824), .op(n9954) );
  mux2_1 U9077 ( .ip1(\ANSWER/mem[4][4][0] ), .ip2(n8840), .s(n9954), .op(
        n3790) );
  nor2_1 U9078 ( .ip1(n8841), .ip2(n8824), .op(n9955) );
  mux2_1 U9079 ( .ip1(\ANSWER/mem[4][5][0] ), .ip2(n8831), .s(n9955), .op(
        n3789) );
  nor2_1 U9080 ( .ip1(n8842), .ip2(n8824), .op(n9956) );
  mux2_1 U9081 ( .ip1(\ANSWER/mem[4][6][0] ), .ip2(n8847), .s(n9956), .op(
        n3788) );
  nor2_1 U9082 ( .ip1(n8843), .ip2(n8824), .op(n9957) );
  mux2_1 U9083 ( .ip1(\ANSWER/mem[4][7][0] ), .ip2(n8831), .s(n9957), .op(
        n3787) );
  nor2_1 U9084 ( .ip1(n8844), .ip2(n8824), .op(n9958) );
  mux2_1 U9085 ( .ip1(\ANSWER/mem[4][8][0] ), .ip2(n8840), .s(n9958), .op(
        n3786) );
  nor2_1 U9086 ( .ip1(n8846), .ip2(n8824), .op(n9959) );
  mux2_1 U9087 ( .ip1(\ANSWER/mem[4][9][0] ), .ip2(n8831), .s(n9959), .op(
        n3785) );
  buf_1 U9088 ( .ip(n11979), .op(n11454) );
  nand4_1 U9089 ( .ip1(n12098), .ip2(n8829), .ip3(n8828), .ip4(n11454), .op(
        n8825) );
  nor2_1 U9090 ( .ip1(n8835), .ip2(n8825), .op(n9960) );
  mux2_1 U9091 ( .ip1(\ANSWER/mem[5][0][0] ), .ip2(n8840), .s(n9960), .op(
        n3784) );
  nor2_1 U9092 ( .ip1(n8836), .ip2(n8825), .op(n9961) );
  mux2_1 U9093 ( .ip1(\ANSWER/mem[5][1][0] ), .ip2(n8847), .s(n9961), .op(
        n3783) );
  nor2_1 U9094 ( .ip1(n8837), .ip2(n8825), .op(n9962) );
  mux2_1 U9095 ( .ip1(\ANSWER/mem[5][2][0] ), .ip2(n8847), .s(n9962), .op(
        n3782) );
  nor2_1 U9096 ( .ip1(n8838), .ip2(n8825), .op(n9963) );
  mux2_1 U9097 ( .ip1(\ANSWER/mem[5][3][0] ), .ip2(n8847), .s(n9963), .op(
        n3781) );
  nor2_1 U9098 ( .ip1(n8839), .ip2(n8825), .op(n9964) );
  mux2_1 U9099 ( .ip1(\ANSWER/mem[5][4][0] ), .ip2(n8847), .s(n9964), .op(
        n3780) );
  nor2_1 U9100 ( .ip1(n8841), .ip2(n8825), .op(n9965) );
  mux2_1 U9101 ( .ip1(\ANSWER/mem[5][5][0] ), .ip2(n8847), .s(n9965), .op(
        n3779) );
  nor2_1 U9102 ( .ip1(n8842), .ip2(n8825), .op(n9966) );
  mux2_1 U9103 ( .ip1(\ANSWER/mem[5][6][0] ), .ip2(n8847), .s(n9966), .op(
        n3778) );
  nor2_1 U9104 ( .ip1(n8843), .ip2(n8825), .op(n9967) );
  mux2_1 U9105 ( .ip1(\ANSWER/mem[5][7][0] ), .ip2(n8847), .s(n9967), .op(
        n3777) );
  nor2_1 U9106 ( .ip1(n8844), .ip2(n8825), .op(n9968) );
  mux2_1 U9107 ( .ip1(\ANSWER/mem[5][8][0] ), .ip2(n8847), .s(n9968), .op(
        n3776) );
  nor2_1 U9108 ( .ip1(n8846), .ip2(n8825), .op(n9969) );
  mux2_1 U9109 ( .ip1(\ANSWER/mem[5][9][0] ), .ip2(n8840), .s(n9969), .op(
        n3775) );
  inv_1 U9110 ( .ip(n12098), .op(n11868) );
  buf_1 U9111 ( .ip(n11979), .op(n11656) );
  nand4_1 U9112 ( .ip1(n8826), .ip2(n8828), .ip3(n11868), .ip4(n11656), .op(
        n8827) );
  nor2_1 U9113 ( .ip1(n8835), .ip2(n8827), .op(n9970) );
  mux2_1 U9114 ( .ip1(\ANSWER/mem[6][0][0] ), .ip2(n8831), .s(n9970), .op(
        n3774) );
  nor2_1 U9115 ( .ip1(n8836), .ip2(n8827), .op(n9971) );
  mux2_1 U9116 ( .ip1(\ANSWER/mem[6][1][0] ), .ip2(n8847), .s(n9971), .op(
        n3773) );
  nor2_1 U9117 ( .ip1(n8837), .ip2(n8827), .op(n9972) );
  mux2_1 U9118 ( .ip1(\ANSWER/mem[6][2][0] ), .ip2(n8847), .s(n9972), .op(
        n3772) );
  nor2_1 U9119 ( .ip1(n8838), .ip2(n8827), .op(n9973) );
  mux2_1 U9120 ( .ip1(\ANSWER/mem[6][3][0] ), .ip2(n8847), .s(n9973), .op(
        n3771) );
  nor2_1 U9121 ( .ip1(n8839), .ip2(n8827), .op(n9974) );
  mux2_1 U9122 ( .ip1(\ANSWER/mem[6][4][0] ), .ip2(n8831), .s(n9974), .op(
        n3770) );
  nor2_1 U9123 ( .ip1(n8841), .ip2(n8827), .op(n9975) );
  mux2_1 U9124 ( .ip1(\ANSWER/mem[6][5][0] ), .ip2(n8840), .s(n9975), .op(
        n3769) );
  nor2_1 U9125 ( .ip1(n8842), .ip2(n8827), .op(n9976) );
  mux2_1 U9126 ( .ip1(\ANSWER/mem[6][6][0] ), .ip2(n8847), .s(n9976), .op(
        n3768) );
  nor2_1 U9127 ( .ip1(n8843), .ip2(n8827), .op(n9977) );
  mux2_1 U9128 ( .ip1(\ANSWER/mem[6][7][0] ), .ip2(n8831), .s(n9977), .op(
        n3767) );
  nor2_1 U9129 ( .ip1(n8844), .ip2(n8827), .op(n9978) );
  mux2_1 U9130 ( .ip1(\ANSWER/mem[6][8][0] ), .ip2(n8831), .s(n9978), .op(
        n3766) );
  nor2_1 U9131 ( .ip1(n8846), .ip2(n8827), .op(n9979) );
  mux2_1 U9132 ( .ip1(\ANSWER/mem[6][9][0] ), .ip2(n8831), .s(n9979), .op(
        n3765) );
  inv_1 U9133 ( .ip(n12098), .op(n11976) );
  buf_1 U9134 ( .ip(n11979), .op(n11440) );
  nand4_1 U9135 ( .ip1(n8829), .ip2(n8828), .ip3(n11976), .ip4(n11440), .op(
        n8830) );
  nor2_1 U9136 ( .ip1(n8835), .ip2(n8830), .op(n9980) );
  mux2_1 U9137 ( .ip1(\ANSWER/mem[7][0][0] ), .ip2(n8847), .s(n9980), .op(
        n3764) );
  nor2_1 U9138 ( .ip1(n8836), .ip2(n8830), .op(n9981) );
  mux2_1 U9139 ( .ip1(\ANSWER/mem[7][1][0] ), .ip2(n8831), .s(n9981), .op(
        n3763) );
  nor2_1 U9140 ( .ip1(n8837), .ip2(n8830), .op(n9983) );
  mux2_1 U9141 ( .ip1(\ANSWER/mem[7][2][0] ), .ip2(n8831), .s(n9983), .op(
        n3762) );
  nor2_1 U9142 ( .ip1(n8838), .ip2(n8830), .op(n9984) );
  mux2_1 U9143 ( .ip1(\ANSWER/mem[7][3][0] ), .ip2(n8840), .s(n9984), .op(
        n3761) );
  nor2_1 U9144 ( .ip1(n8839), .ip2(n8830), .op(n9985) );
  mux2_1 U9145 ( .ip1(\ANSWER/mem[7][4][0] ), .ip2(n8847), .s(n9985), .op(
        n3760) );
  nor2_1 U9146 ( .ip1(n8841), .ip2(n8830), .op(n9986) );
  mux2_1 U9147 ( .ip1(\ANSWER/mem[7][5][0] ), .ip2(n8840), .s(n9986), .op(
        n3759) );
  nor2_1 U9148 ( .ip1(n8842), .ip2(n8830), .op(n9987) );
  mux2_1 U9149 ( .ip1(\ANSWER/mem[7][6][0] ), .ip2(n8847), .s(n9987), .op(
        n3758) );
  nor2_1 U9150 ( .ip1(n8843), .ip2(n8830), .op(n9988) );
  mux2_1 U9151 ( .ip1(\ANSWER/mem[7][7][0] ), .ip2(n8847), .s(n9988), .op(
        n3757) );
  nor2_1 U9152 ( .ip1(n8844), .ip2(n8830), .op(n9989) );
  mux2_1 U9153 ( .ip1(\ANSWER/mem[7][8][0] ), .ip2(n8847), .s(n9989), .op(
        n3756) );
  nor2_1 U9154 ( .ip1(n8846), .ip2(n8830), .op(n9990) );
  mux2_1 U9155 ( .ip1(\ANSWER/mem[7][9][0] ), .ip2(n8831), .s(n9990), .op(
        n3755) );
  nand3_1 U9156 ( .ip1(n12109), .ip2(n8834), .ip3(n11336), .op(n8832) );
  nor2_1 U9157 ( .ip1(n8835), .ip2(n8832), .op(n9991) );
  mux2_1 U9158 ( .ip1(\ANSWER/mem[8][0][0] ), .ip2(n8831), .s(n9991), .op(
        n3754) );
  nor2_1 U9159 ( .ip1(n8836), .ip2(n8832), .op(n9992) );
  mux2_1 U9160 ( .ip1(\ANSWER/mem[8][1][0] ), .ip2(n8831), .s(n9992), .op(
        n3753) );
  nor2_1 U9161 ( .ip1(n8837), .ip2(n8832), .op(n9993) );
  mux2_1 U9162 ( .ip1(\ANSWER/mem[8][2][0] ), .ip2(n8840), .s(n9993), .op(
        n3752) );
  nor2_1 U9163 ( .ip1(n8838), .ip2(n8832), .op(n9994) );
  mux2_1 U9164 ( .ip1(\ANSWER/mem[8][3][0] ), .ip2(n8847), .s(n9994), .op(
        n3751) );
  nor2_1 U9165 ( .ip1(n8839), .ip2(n8832), .op(n9996) );
  mux2_1 U9166 ( .ip1(\ANSWER/mem[8][4][0] ), .ip2(n8847), .s(n9996), .op(
        n3750) );
  nor2_1 U9167 ( .ip1(n8841), .ip2(n8832), .op(n9997) );
  mux2_1 U9168 ( .ip1(\ANSWER/mem[8][5][0] ), .ip2(n8840), .s(n9997), .op(
        n3749) );
  nor2_1 U9169 ( .ip1(n8842), .ip2(n8832), .op(n9998) );
  mux2_1 U9170 ( .ip1(\ANSWER/mem[8][6][0] ), .ip2(n8847), .s(n9998), .op(
        n3748) );
  nor2_1 U9171 ( .ip1(n8843), .ip2(n8832), .op(n9999) );
  mux2_1 U9172 ( .ip1(\ANSWER/mem[8][7][0] ), .ip2(n8840), .s(n9999), .op(
        n3747) );
  nor2_1 U9173 ( .ip1(n8844), .ip2(n8832), .op(n10000) );
  mux2_1 U9174 ( .ip1(\ANSWER/mem[8][8][0] ), .ip2(n8847), .s(n10000), .op(
        n3746) );
  nor2_1 U9175 ( .ip1(n8846), .ip2(n8832), .op(n10001) );
  mux2_1 U9176 ( .ip1(\ANSWER/mem[8][9][0] ), .ip2(n8840), .s(n10001), .op(
        n3745) );
  nand3_1 U9177 ( .ip1(n8834), .ip2(n8833), .ip3(n11336), .op(n8845) );
  nor2_1 U9178 ( .ip1(n8835), .ip2(n8845), .op(n10002) );
  mux2_1 U9179 ( .ip1(\ANSWER/mem[9][0][0] ), .ip2(n8847), .s(n10002), .op(
        n3744) );
  nor2_1 U9180 ( .ip1(n8836), .ip2(n8845), .op(n10003) );
  mux2_1 U9181 ( .ip1(\ANSWER/mem[9][1][0] ), .ip2(n8840), .s(n10003), .op(
        n3743) );
  nor2_1 U9182 ( .ip1(n8837), .ip2(n8845), .op(n10004) );
  mux2_1 U9183 ( .ip1(\ANSWER/mem[9][2][0] ), .ip2(n8840), .s(n10004), .op(
        n3742) );
  nor2_1 U9184 ( .ip1(n8838), .ip2(n8845), .op(n10005) );
  mux2_1 U9185 ( .ip1(\ANSWER/mem[9][3][0] ), .ip2(n8847), .s(n10005), .op(
        n3741) );
  nor2_1 U9186 ( .ip1(n8839), .ip2(n8845), .op(n10006) );
  mux2_1 U9187 ( .ip1(\ANSWER/mem[9][4][0] ), .ip2(n8840), .s(n10006), .op(
        n3740) );
  nor2_1 U9188 ( .ip1(n8841), .ip2(n8845), .op(n10007) );
  mux2_1 U9189 ( .ip1(\ANSWER/mem[9][5][0] ), .ip2(n8847), .s(n10007), .op(
        n3739) );
  nor2_1 U9190 ( .ip1(n8842), .ip2(n8845), .op(n10008) );
  mux2_1 U9191 ( .ip1(\ANSWER/mem[9][6][0] ), .ip2(n8847), .s(n10008), .op(
        n3738) );
  nor2_1 U9192 ( .ip1(n8843), .ip2(n8845), .op(n10009) );
  mux2_1 U9193 ( .ip1(\ANSWER/mem[9][7][0] ), .ip2(n8847), .s(n10009), .op(
        n3737) );
  nor2_1 U9194 ( .ip1(n8844), .ip2(n8845), .op(n10010) );
  mux2_1 U9195 ( .ip1(\ANSWER/mem[9][8][0] ), .ip2(n8847), .s(n10010), .op(
        n3736) );
  nor2_1 U9196 ( .ip1(n8846), .ip2(n8845), .op(n10011) );
  mux2_1 U9197 ( .ip1(\ANSWER/mem[9][9][0] ), .ip2(n8847), .s(n10011), .op(
        n3735) );
  fulladder U9198 ( .a(n8850), .b(n8849), .ci(n8848), .co(n8896), .s(n8852) );
  inv_1 U9199 ( .ip(n8896), .op(n8906) );
  fulladder U9200 ( .a(n8853), .b(n8852), .ci(n8851), .co(n8908), .s(n8777) );
  inv_1 U9201 ( .ip(q_w2[9]), .op(n9864) );
  nor2_1 U9202 ( .ip1(n9530), .ip2(n9864), .op(n9056) );
  and2_1 U9203 ( .ip1(n9056), .ip2(n8854), .op(n8921) );
  nor2_1 U9204 ( .ip1(n9335), .ip2(n9864), .op(n8855) );
  or2_1 U9205 ( .ip1(q_w2[6]), .ip2(n8855), .op(n8857) );
  or2_1 U9206 ( .ip1(m2DataIn[3]), .ip2(n8855), .op(n8856) );
  nand2_1 U9207 ( .ip1(n8857), .ip2(n8856), .op(n8920) );
  nor2_1 U9208 ( .ip1(n8921), .ip2(n8920), .op(n8859) );
  nand2_1 U9209 ( .ip1(m2DataIn[9]), .ip2(q_w2[0]), .op(n8858) );
  xor2_1 U9210 ( .ip1(n8859), .ip2(n8858), .op(n8941) );
  nand2_1 U9211 ( .ip1(m2DataIn[4]), .ip2(q_w2[5]), .op(n8915) );
  nor4_1 U9212 ( .ip1(n9702), .ip2(n9640), .ip3(n9638), .ip4(n9703), .op(n8935) );
  or2_1 U9213 ( .ip1(n8915), .ip2(n8935), .op(n8862) );
  or2_1 U9214 ( .ip1(n8860), .ip2(n8935), .op(n8861) );
  nand2_1 U9215 ( .ip1(n8862), .ip2(n8861), .op(n8934) );
  nor2_1 U9216 ( .ip1(n9817), .ip2(n9334), .op(n8936) );
  xnor2_1 U9217 ( .ip1(n8934), .ip2(n8936), .op(n8940) );
  fulladder U9218 ( .a(n8864), .b(n8880), .ci(n8863), .co(n8939), .s(n8893) );
  or2_1 U9219 ( .ip1(n8865), .ip2(n8866), .op(n8869) );
  or2_1 U9220 ( .ip1(n8867), .ip2(n8866), .op(n8868) );
  nand2_1 U9221 ( .ip1(n8869), .ip2(n8868), .op(n8954) );
  nand2_1 U9222 ( .ip1(m2DataIn[2]), .ip2(q_w2[7]), .op(n9386) );
  inv_1 U9223 ( .ip(q_w2[8]), .op(n9788) );
  nor3_1 U9224 ( .ip1(n9500), .ip2(n9788), .ip3(n8870), .op(n8924) );
  or2_1 U9225 ( .ip1(n9386), .ip2(n8924), .op(n8872) );
  nand2_1 U9226 ( .ip1(m2DataIn[1]), .ip2(q_w2[8]), .op(n8928) );
  or2_1 U9227 ( .ip1(n8928), .ip2(n8924), .op(n8871) );
  nand2_1 U9228 ( .ip1(n8872), .ip2(n8871), .op(n8925) );
  mux2_1 U9229 ( .ip1(n8873), .ip2(rdata[1]), .s(n8925), .op(n8953) );
  or2_1 U9230 ( .ip1(n8874), .ip2(n8875), .op(n8878) );
  or2_1 U9231 ( .ip1(n8876), .ip2(n8875), .op(n8877) );
  nand2_1 U9232 ( .ip1(n8878), .ip2(n8877), .op(n8952) );
  inv_1 U9233 ( .ip(n8879), .op(n8958) );
  nor3_1 U9234 ( .ip1(n9725), .ip2(n9372), .ip3(n8880), .op(n8944) );
  nor2_1 U9235 ( .ip1(n9467), .ip2(n9372), .op(n8881) );
  or2_1 U9236 ( .ip1(q_w2[2]), .ip2(n8881), .op(n8883) );
  or2_1 U9237 ( .ip1(m2DataIn[7]), .ip2(n8881), .op(n8882) );
  nand2_1 U9238 ( .ip1(n8883), .ip2(n8882), .op(n8884) );
  nor2_1 U9239 ( .ip1(n8944), .ip2(n8884), .op(n8943) );
  nand2_1 U9240 ( .ip1(rdata[0]), .ip2(n8885), .op(n8886) );
  nand2_1 U9241 ( .ip1(n8887), .ip2(n8886), .op(n8945) );
  xor2_1 U9242 ( .ip1(n8943), .ip2(n8945), .op(n8957) );
  fulladder U9243 ( .a(n8890), .b(n8889), .ci(n8888), .co(n8956), .s(n8849) );
  inv_1 U9244 ( .ip(n8891), .op(n8963) );
  fulladder U9245 ( .a(n8894), .b(n8893), .ci(n8892), .co(n8962), .s(n8773) );
  xor2_1 U9246 ( .ip1(n8908), .ip2(n8904), .op(n8895) );
  mux2_1 U9247 ( .ip1(n8906), .ip2(n8896), .s(n8895), .op(n8898) );
  inv_1 U9248 ( .ip(\SIGMOID/sign_bit ), .op(n9187) );
  and2_1 U9249 ( .ip1(n9187), .ip2(\SIGMOID/N64 ), .op(n8897) );
  xor2_1 U9250 ( .ip1(\SIGMOID/lut_out [1]), .ip2(n8897), .op(n10232) );
  mux2_1 U9251 ( .ip1(n8898), .ip2(n10232), .s(n9907), .op(n8900) );
  buf_1 U9252 ( .ip(n8900), .op(n8899) );
  mux2_1 U9253 ( .ip1(\ANSWER/mem[0][0][1] ), .ip2(n8899), .s(n9910), .op(
        n3734) );
  mux2_1 U9254 ( .ip1(\ANSWER/mem[0][1][1] ), .ip2(n8899), .s(n9911), .op(
        n3733) );
  mux2_1 U9255 ( .ip1(\ANSWER/mem[0][2][1] ), .ip2(n8899), .s(n9912), .op(
        n3732) );
  mux2_1 U9256 ( .ip1(\ANSWER/mem[0][3][1] ), .ip2(n8899), .s(n9913), .op(
        n3731) );
  mux2_1 U9257 ( .ip1(\ANSWER/mem[0][4][1] ), .ip2(n8899), .s(n9914), .op(
        n3730) );
  mux2_1 U9258 ( .ip1(\ANSWER/mem[0][5][1] ), .ip2(n8899), .s(n9915), .op(
        n3729) );
  mux2_1 U9259 ( .ip1(\ANSWER/mem[0][6][1] ), .ip2(n8899), .s(n9916), .op(
        n3728) );
  mux2_1 U9260 ( .ip1(\ANSWER/mem[0][7][1] ), .ip2(n8899), .s(n9917), .op(
        n3727) );
  mux2_1 U9261 ( .ip1(\ANSWER/mem[0][8][1] ), .ip2(n8899), .s(n9918), .op(
        n3726) );
  mux2_1 U9262 ( .ip1(\ANSWER/mem[0][9][1] ), .ip2(n8899), .s(n9919), .op(
        n3725) );
  mux2_1 U9263 ( .ip1(\ANSWER/mem[1][0][1] ), .ip2(n8899), .s(n9920), .op(
        n3724) );
  mux2_1 U9264 ( .ip1(\ANSWER/mem[1][1][1] ), .ip2(n8899), .s(n9921), .op(
        n3723) );
  mux2_1 U9265 ( .ip1(\ANSWER/mem[1][2][1] ), .ip2(n8899), .s(n9922), .op(
        n3722) );
  mux2_1 U9266 ( .ip1(\ANSWER/mem[1][3][1] ), .ip2(n8899), .s(n9923), .op(
        n3721) );
  mux2_1 U9267 ( .ip1(\ANSWER/mem[1][4][1] ), .ip2(n8899), .s(n9924), .op(
        n3720) );
  mux2_1 U9268 ( .ip1(\ANSWER/mem[1][5][1] ), .ip2(n8899), .s(n9925), .op(
        n3719) );
  mux2_1 U9269 ( .ip1(\ANSWER/mem[1][6][1] ), .ip2(n8899), .s(n9926), .op(
        n3718) );
  mux2_1 U9270 ( .ip1(\ANSWER/mem[1][7][1] ), .ip2(n8899), .s(n9927), .op(
        n3717) );
  mux2_1 U9271 ( .ip1(\ANSWER/mem[1][8][1] ), .ip2(n8899), .s(n9928), .op(
        n3716) );
  mux2_1 U9272 ( .ip1(\ANSWER/mem[1][9][1] ), .ip2(n8899), .s(n9929), .op(
        n3715) );
  mux2_1 U9273 ( .ip1(\ANSWER/mem[2][0][1] ), .ip2(n8899), .s(n9930), .op(
        n3714) );
  mux2_1 U9274 ( .ip1(\ANSWER/mem[2][1][1] ), .ip2(n8899), .s(n9931), .op(
        n3713) );
  mux2_1 U9275 ( .ip1(\ANSWER/mem[2][2][1] ), .ip2(n8899), .s(n9932), .op(
        n3712) );
  mux2_1 U9276 ( .ip1(\ANSWER/mem[2][3][1] ), .ip2(n8899), .s(n9933), .op(
        n3711) );
  mux2_1 U9277 ( .ip1(\ANSWER/mem[2][4][1] ), .ip2(n8899), .s(n9934), .op(
        n3710) );
  mux2_1 U9278 ( .ip1(\ANSWER/mem[2][5][1] ), .ip2(n8899), .s(n9935), .op(
        n3709) );
  mux2_1 U9279 ( .ip1(\ANSWER/mem[2][6][1] ), .ip2(n8899), .s(n9936), .op(
        n3708) );
  mux2_1 U9280 ( .ip1(\ANSWER/mem[2][7][1] ), .ip2(n8899), .s(n9937), .op(
        n3707) );
  mux2_1 U9281 ( .ip1(\ANSWER/mem[2][8][1] ), .ip2(n8899), .s(n9938), .op(
        n3706) );
  mux2_1 U9282 ( .ip1(\ANSWER/mem[2][9][1] ), .ip2(n8899), .s(n9939), .op(
        n3705) );
  mux2_1 U9283 ( .ip1(\ANSWER/mem[3][0][1] ), .ip2(n8899), .s(n9940), .op(
        n3704) );
  mux2_1 U9284 ( .ip1(\ANSWER/mem[3][1][1] ), .ip2(n8899), .s(n9941), .op(
        n3703) );
  mux2_1 U9285 ( .ip1(\ANSWER/mem[3][2][1] ), .ip2(n8899), .s(n9942), .op(
        n3702) );
  mux2_1 U9286 ( .ip1(\ANSWER/mem[3][3][1] ), .ip2(n8899), .s(n9943), .op(
        n3701) );
  mux2_1 U9287 ( .ip1(\ANSWER/mem[3][4][1] ), .ip2(n8899), .s(n9944), .op(
        n3700) );
  mux2_1 U9288 ( .ip1(\ANSWER/mem[3][5][1] ), .ip2(n8899), .s(n9945), .op(
        n3699) );
  mux2_1 U9289 ( .ip1(\ANSWER/mem[3][6][1] ), .ip2(n8901), .s(n9946), .op(
        n3698) );
  mux2_1 U9290 ( .ip1(\ANSWER/mem[3][7][1] ), .ip2(n8900), .s(n9947), .op(
        n3697) );
  mux2_1 U9291 ( .ip1(\ANSWER/mem[3][8][1] ), .ip2(n8900), .s(n9948), .op(
        n3696) );
  mux2_1 U9292 ( .ip1(\ANSWER/mem[3][9][1] ), .ip2(n8900), .s(n9949), .op(
        n3695) );
  mux2_1 U9293 ( .ip1(\ANSWER/mem[4][0][1] ), .ip2(n8900), .s(n9950), .op(
        n3694) );
  mux2_1 U9294 ( .ip1(\ANSWER/mem[4][1][1] ), .ip2(n8900), .s(n9951), .op(
        n3693) );
  mux2_1 U9295 ( .ip1(\ANSWER/mem[4][2][1] ), .ip2(n8901), .s(n9952), .op(
        n3692) );
  mux2_1 U9296 ( .ip1(\ANSWER/mem[4][3][1] ), .ip2(n8901), .s(n9953), .op(
        n3691) );
  mux2_1 U9297 ( .ip1(\ANSWER/mem[4][4][1] ), .ip2(n8901), .s(n9954), .op(
        n3690) );
  mux2_1 U9298 ( .ip1(\ANSWER/mem[4][5][1] ), .ip2(n8901), .s(n9955), .op(
        n3689) );
  mux2_1 U9299 ( .ip1(\ANSWER/mem[4][6][1] ), .ip2(n8901), .s(n9956), .op(
        n3688) );
  mux2_1 U9300 ( .ip1(\ANSWER/mem[4][7][1] ), .ip2(n8901), .s(n9957), .op(
        n3687) );
  mux2_1 U9301 ( .ip1(\ANSWER/mem[4][8][1] ), .ip2(n8901), .s(n9958), .op(
        n3686) );
  mux2_1 U9302 ( .ip1(\ANSWER/mem[4][9][1] ), .ip2(n8901), .s(n9959), .op(
        n3685) );
  mux2_1 U9303 ( .ip1(\ANSWER/mem[5][0][1] ), .ip2(n8901), .s(n9960), .op(
        n3684) );
  mux2_1 U9304 ( .ip1(\ANSWER/mem[5][1][1] ), .ip2(n8900), .s(n9961), .op(
        n3683) );
  mux2_1 U9305 ( .ip1(\ANSWER/mem[5][2][1] ), .ip2(n8901), .s(n9962), .op(
        n3682) );
  mux2_1 U9306 ( .ip1(\ANSWER/mem[5][3][1] ), .ip2(n8900), .s(n9963), .op(
        n3681) );
  mux2_1 U9307 ( .ip1(\ANSWER/mem[5][4][1] ), .ip2(n8900), .s(n9964), .op(
        n3680) );
  mux2_1 U9308 ( .ip1(\ANSWER/mem[5][5][1] ), .ip2(n8900), .s(n9965), .op(
        n3679) );
  mux2_1 U9309 ( .ip1(\ANSWER/mem[5][6][1] ), .ip2(n8900), .s(n9966), .op(
        n3678) );
  mux2_1 U9310 ( .ip1(\ANSWER/mem[5][7][1] ), .ip2(n8900), .s(n9967), .op(
        n3677) );
  mux2_1 U9311 ( .ip1(\ANSWER/mem[5][8][1] ), .ip2(n8900), .s(n9968), .op(
        n3676) );
  mux2_1 U9312 ( .ip1(\ANSWER/mem[5][9][1] ), .ip2(n8900), .s(n9969), .op(
        n3675) );
  mux2_1 U9313 ( .ip1(\ANSWER/mem[6][0][1] ), .ip2(n8900), .s(n9970), .op(
        n3674) );
  mux2_1 U9314 ( .ip1(\ANSWER/mem[6][1][1] ), .ip2(n8900), .s(n9971), .op(
        n3673) );
  mux2_1 U9315 ( .ip1(\ANSWER/mem[6][2][1] ), .ip2(n8900), .s(n9972), .op(
        n3672) );
  mux2_1 U9316 ( .ip1(\ANSWER/mem[6][3][1] ), .ip2(n8900), .s(n9973), .op(
        n3671) );
  mux2_1 U9317 ( .ip1(\ANSWER/mem[6][4][1] ), .ip2(n8900), .s(n9974), .op(
        n3670) );
  mux2_1 U9318 ( .ip1(\ANSWER/mem[6][5][1] ), .ip2(n8900), .s(n9975), .op(
        n3669) );
  mux2_1 U9319 ( .ip1(\ANSWER/mem[6][6][1] ), .ip2(n8900), .s(n9976), .op(
        n3668) );
  mux2_1 U9320 ( .ip1(\ANSWER/mem[6][7][1] ), .ip2(n8900), .s(n9977), .op(
        n3667) );
  mux2_1 U9321 ( .ip1(\ANSWER/mem[6][8][1] ), .ip2(n8900), .s(n9978), .op(
        n3666) );
  mux2_1 U9322 ( .ip1(\ANSWER/mem[6][9][1] ), .ip2(n8900), .s(n9979), .op(
        n3665) );
  mux2_1 U9323 ( .ip1(\ANSWER/mem[7][0][1] ), .ip2(n8900), .s(n9980), .op(
        n3664) );
  mux2_1 U9324 ( .ip1(\ANSWER/mem[7][1][1] ), .ip2(n8900), .s(n9981), .op(
        n3663) );
  buf_1 U9325 ( .ip(n8900), .op(n8901) );
  mux2_1 U9326 ( .ip1(\ANSWER/mem[7][2][1] ), .ip2(n8901), .s(n9983), .op(
        n3662) );
  mux2_1 U9327 ( .ip1(\ANSWER/mem[7][3][1] ), .ip2(n8901), .s(n9984), .op(
        n3661) );
  mux2_1 U9328 ( .ip1(\ANSWER/mem[7][4][1] ), .ip2(n8901), .s(n9985), .op(
        n3660) );
  mux2_1 U9329 ( .ip1(\ANSWER/mem[7][5][1] ), .ip2(n8901), .s(n9986), .op(
        n3659) );
  mux2_1 U9330 ( .ip1(\ANSWER/mem[7][6][1] ), .ip2(n8901), .s(n9987), .op(
        n3658) );
  mux2_1 U9331 ( .ip1(\ANSWER/mem[7][7][1] ), .ip2(n8901), .s(n9988), .op(
        n3657) );
  mux2_1 U9332 ( .ip1(\ANSWER/mem[7][8][1] ), .ip2(n8901), .s(n9989), .op(
        n3656) );
  mux2_1 U9333 ( .ip1(\ANSWER/mem[7][9][1] ), .ip2(n8900), .s(n9990), .op(
        n3655) );
  mux2_1 U9334 ( .ip1(\ANSWER/mem[8][0][1] ), .ip2(n8901), .s(n9991), .op(
        n3654) );
  mux2_1 U9335 ( .ip1(\ANSWER/mem[8][1][1] ), .ip2(n8901), .s(n9992), .op(
        n3653) );
  mux2_1 U9336 ( .ip1(\ANSWER/mem[8][2][1] ), .ip2(n8901), .s(n9993), .op(
        n3652) );
  mux2_1 U9337 ( .ip1(\ANSWER/mem[8][3][1] ), .ip2(n8901), .s(n9994), .op(
        n3651) );
  mux2_1 U9338 ( .ip1(\ANSWER/mem[8][4][1] ), .ip2(n8900), .s(n9996), .op(
        n3650) );
  mux2_1 U9339 ( .ip1(\ANSWER/mem[8][5][1] ), .ip2(n8900), .s(n9997), .op(
        n3649) );
  mux2_1 U9340 ( .ip1(\ANSWER/mem[8][6][1] ), .ip2(n8900), .s(n9998), .op(
        n3648) );
  mux2_1 U9341 ( .ip1(\ANSWER/mem[8][7][1] ), .ip2(n8900), .s(n9999), .op(
        n3647) );
  mux2_1 U9342 ( .ip1(\ANSWER/mem[8][8][1] ), .ip2(n8900), .s(n10000), .op(
        n3646) );
  mux2_1 U9343 ( .ip1(\ANSWER/mem[8][9][1] ), .ip2(n8900), .s(n10001), .op(
        n3645) );
  mux2_1 U9344 ( .ip1(\ANSWER/mem[9][0][1] ), .ip2(n8900), .s(n10002), .op(
        n3644) );
  mux2_1 U9345 ( .ip1(\ANSWER/mem[9][1][1] ), .ip2(n8900), .s(n10003), .op(
        n3643) );
  mux2_1 U9346 ( .ip1(\ANSWER/mem[9][2][1] ), .ip2(n8900), .s(n10004), .op(
        n3642) );
  mux2_1 U9347 ( .ip1(\ANSWER/mem[9][3][1] ), .ip2(n8900), .s(n10005), .op(
        n3641) );
  mux2_1 U9348 ( .ip1(\ANSWER/mem[9][4][1] ), .ip2(n8900), .s(n10006), .op(
        n3640) );
  mux2_1 U9349 ( .ip1(\ANSWER/mem[9][5][1] ), .ip2(n8900), .s(n10007), .op(
        n3639) );
  mux2_1 U9350 ( .ip1(\ANSWER/mem[9][6][1] ), .ip2(n8901), .s(n10008), .op(
        n3638) );
  mux2_1 U9351 ( .ip1(\ANSWER/mem[9][7][1] ), .ip2(n8901), .s(n10009), .op(
        n3637) );
  mux2_1 U9352 ( .ip1(\ANSWER/mem[9][8][1] ), .ip2(n8901), .s(n10010), .op(
        n3636) );
  mux2_1 U9353 ( .ip1(\ANSWER/mem[9][9][1] ), .ip2(n8901), .s(n10011), .op(
        n3635) );
  nor2_1 U9354 ( .ip1(\SIGMOID/lut_out [1]), .ip2(\SIGMOID/N64 ), .op(n8902)
         );
  nor2_1 U9355 ( .ip1(\SIGMOID/sign_bit ), .ip2(n8902), .op(n8903) );
  xor2_1 U9356 ( .ip1(\SIGMOID/lut_out [2]), .ip2(n8903), .op(n10264) );
  inv_1 U9357 ( .ip(n8904), .op(n8907) );
  nor2_1 U9358 ( .ip1(n8908), .ip2(n8907), .op(n8905) );
  or2_1 U9359 ( .ip1(n8906), .ip2(n8905), .op(n8910) );
  nand2_1 U9360 ( .ip1(n8908), .ip2(n8907), .op(n8909) );
  nand2_1 U9361 ( .ip1(n8910), .ip2(n8909), .op(n8960) );
  nand2_1 U9362 ( .ip1(m2DataIn[7]), .ip2(q_w2[3]), .op(n8911) );
  nand2_1 U9363 ( .ip1(m2DataIn[7]), .ip2(q_w2[4]), .op(n8982) );
  nor3_1 U9364 ( .ip1(n9467), .ip2(n9372), .ip3(n8982), .op(n9001) );
  or2_1 U9365 ( .ip1(n8911), .ip2(n9001), .op(n8914) );
  nand2_1 U9366 ( .ip1(m2DataIn[6]), .ip2(q_w2[4]), .op(n8912) );
  or2_1 U9367 ( .ip1(n8912), .ip2(n9001), .op(n8913) );
  nand2_1 U9368 ( .ip1(n8914), .ip2(n8913), .op(n9000) );
  nor2_1 U9369 ( .ip1(n9817), .ip2(n9499), .op(n9002) );
  xor2_1 U9370 ( .ip1(n9000), .ip2(n9002), .op(n9019) );
  nand2_1 U9371 ( .ip1(m2DataIn[4]), .ip2(q_w2[6]), .op(n8916) );
  nand2_1 U9372 ( .ip1(m2DataIn[5]), .ip2(q_w2[6]), .op(n8978) );
  nor2_1 U9373 ( .ip1(n8978), .ip2(n8915), .op(n8991) );
  or2_1 U9374 ( .ip1(n8916), .ip2(n8991), .op(n8919) );
  nand2_1 U9375 ( .ip1(m2DataIn[5]), .ip2(q_w2[5]), .op(n8917) );
  or2_1 U9376 ( .ip1(n8917), .ip2(n8991), .op(n8918) );
  nand2_1 U9377 ( .ip1(n8919), .ip2(n8918), .op(n8990) );
  inv_1 U9378 ( .ip(m2DataIn[9]), .op(n9790) );
  nor2_1 U9379 ( .ip1(n9790), .ip2(n9334), .op(n8992) );
  xor2_1 U9380 ( .ip1(n8990), .ip2(n8992), .op(n9018) );
  nor3_1 U9381 ( .ip1(n8920), .ip2(n9790), .ip3(n9141), .op(n8922) );
  or2_1 U9382 ( .ip1(n8922), .ip2(n8921), .op(n9017) );
  inv_1 U9383 ( .ip(n8923), .op(n9026) );
  or2_1 U9384 ( .ip1(rdata[1]), .ip2(n8924), .op(n8927) );
  or2_1 U9385 ( .ip1(n8925), .ip2(n8924), .op(n8926) );
  nand2_1 U9386 ( .ip1(n8927), .ip2(n8926), .op(n9023) );
  inv_1 U9387 ( .ip(rdata[2]), .op(n8933) );
  nand2_1 U9388 ( .ip1(m2DataIn[1]), .ip2(q_w2[9]), .op(n8929) );
  nand2_1 U9389 ( .ip1(m2DataIn[2]), .ip2(q_w2[9]), .op(n8996) );
  nor2_1 U9390 ( .ip1(n8996), .ip2(n8928), .op(n9008) );
  or2_1 U9391 ( .ip1(n8929), .ip2(n9008), .op(n8932) );
  nand2_1 U9392 ( .ip1(m2DataIn[2]), .ip2(q_w2[8]), .op(n8930) );
  or2_1 U9393 ( .ip1(n8930), .ip2(n9008), .op(n8931) );
  nand2_1 U9394 ( .ip1(n8932), .ip2(n8931), .op(n9009) );
  mux2_1 U9395 ( .ip1(n8933), .ip2(rdata[2]), .s(n9009), .op(n9022) );
  or2_1 U9396 ( .ip1(n8934), .ip2(n8935), .op(n8938) );
  or2_1 U9397 ( .ip1(n8936), .ip2(n8935), .op(n8937) );
  nand2_1 U9398 ( .ip1(n8938), .ip2(n8937), .op(n9021) );
  fulladder U9399 ( .a(n8941), .b(n8940), .ci(n8939), .co(n9024), .s(n8964) );
  inv_1 U9400 ( .ip(n8942), .op(n9034) );
  or2_1 U9401 ( .ip1(n8943), .ip2(n8944), .op(n8947) );
  or2_1 U9402 ( .ip1(n8945), .ip2(n8944), .op(n8946) );
  nand2_1 U9403 ( .ip1(n8947), .ip2(n8946), .op(n9007) );
  nand2_1 U9404 ( .ip1(m2DataIn[3]), .ip2(q_w2[7]), .op(n8949) );
  inv_1 U9405 ( .ip(q_w2[10]), .op(n9814) );
  nor3_1 U9406 ( .ip1(n9530), .ip2(n9814), .ip3(n8948), .op(n9013) );
  or2_1 U9407 ( .ip1(n8949), .ip2(n9013), .op(n8951) );
  nand2_1 U9408 ( .ip1(m2DataIn[0]), .ip2(q_w2[10]), .op(n9136) );
  or2_1 U9409 ( .ip1(n9136), .ip2(n9013), .op(n8950) );
  nand2_1 U9410 ( .ip1(n8951), .ip2(n8950), .op(n9012) );
  nor2_1 U9411 ( .ip1(n9792), .ip2(n9141), .op(n9014) );
  xnor2_1 U9412 ( .ip1(n9012), .ip2(n9014), .op(n9006) );
  fulladder U9413 ( .a(n8954), .b(n8953), .ci(n8952), .co(n9005), .s(n8879) );
  inv_1 U9414 ( .ip(n8955), .op(n9033) );
  fulladder U9415 ( .a(n8958), .b(n8957), .ci(n8956), .co(n9032), .s(n8891) );
  nor2_1 U9416 ( .ip1(n8960), .ip2(n8959), .op(n9028) );
  inv_1 U9417 ( .ip(n9028), .op(n8961) );
  nand2_1 U9418 ( .ip1(n8960), .ip2(n8959), .op(n9030) );
  nand2_1 U9419 ( .ip1(n8961), .ip2(n9030), .op(n8965) );
  fulladder U9420 ( .a(n8964), .b(n8963), .ci(n8962), .co(n9029), .s(n8904) );
  xor2_1 U9421 ( .ip1(n8965), .ip2(n9029), .op(n8966) );
  mux2_1 U9422 ( .ip1(n10264), .ip2(n8966), .s(n9445), .op(n8968) );
  buf_1 U9423 ( .ip(n8968), .op(n8967) );
  mux2_1 U9424 ( .ip1(\ANSWER/mem[0][0][2] ), .ip2(n8967), .s(n9910), .op(
        n3634) );
  mux2_1 U9425 ( .ip1(\ANSWER/mem[0][1][2] ), .ip2(n8967), .s(n9911), .op(
        n3633) );
  mux2_1 U9426 ( .ip1(\ANSWER/mem[0][2][2] ), .ip2(n8967), .s(n9912), .op(
        n3632) );
  mux2_1 U9427 ( .ip1(\ANSWER/mem[0][3][2] ), .ip2(n8967), .s(n9913), .op(
        n3631) );
  mux2_1 U9428 ( .ip1(\ANSWER/mem[0][4][2] ), .ip2(n8967), .s(n9914), .op(
        n3630) );
  mux2_1 U9429 ( .ip1(\ANSWER/mem[0][5][2] ), .ip2(n8967), .s(n9915), .op(
        n3629) );
  mux2_1 U9430 ( .ip1(\ANSWER/mem[0][6][2] ), .ip2(n8967), .s(n9916), .op(
        n3628) );
  mux2_1 U9431 ( .ip1(\ANSWER/mem[0][7][2] ), .ip2(n8967), .s(n9917), .op(
        n3627) );
  mux2_1 U9432 ( .ip1(\ANSWER/mem[0][8][2] ), .ip2(n8967), .s(n9918), .op(
        n3626) );
  mux2_1 U9433 ( .ip1(\ANSWER/mem[0][9][2] ), .ip2(n8967), .s(n9919), .op(
        n3625) );
  mux2_1 U9434 ( .ip1(\ANSWER/mem[1][0][2] ), .ip2(n8967), .s(n9920), .op(
        n3624) );
  mux2_1 U9435 ( .ip1(\ANSWER/mem[1][1][2] ), .ip2(n8967), .s(n9921), .op(
        n3623) );
  mux2_1 U9436 ( .ip1(\ANSWER/mem[1][2][2] ), .ip2(n8967), .s(n9922), .op(
        n3622) );
  mux2_1 U9437 ( .ip1(\ANSWER/mem[1][3][2] ), .ip2(n8967), .s(n9923), .op(
        n3621) );
  mux2_1 U9438 ( .ip1(\ANSWER/mem[1][4][2] ), .ip2(n8967), .s(n9924), .op(
        n3620) );
  mux2_1 U9439 ( .ip1(\ANSWER/mem[1][5][2] ), .ip2(n8967), .s(n9925), .op(
        n3619) );
  mux2_1 U9440 ( .ip1(\ANSWER/mem[1][6][2] ), .ip2(n8967), .s(n9926), .op(
        n3618) );
  mux2_1 U9441 ( .ip1(\ANSWER/mem[1][7][2] ), .ip2(n8967), .s(n9927), .op(
        n3617) );
  mux2_1 U9442 ( .ip1(\ANSWER/mem[1][8][2] ), .ip2(n8967), .s(n9928), .op(
        n3616) );
  mux2_1 U9443 ( .ip1(\ANSWER/mem[1][9][2] ), .ip2(n8967), .s(n9929), .op(
        n3615) );
  mux2_1 U9444 ( .ip1(\ANSWER/mem[2][0][2] ), .ip2(n8967), .s(n9930), .op(
        n3614) );
  mux2_1 U9445 ( .ip1(\ANSWER/mem[2][1][2] ), .ip2(n8967), .s(n9931), .op(
        n3613) );
  mux2_1 U9446 ( .ip1(\ANSWER/mem[2][2][2] ), .ip2(n8967), .s(n9932), .op(
        n3612) );
  mux2_1 U9447 ( .ip1(\ANSWER/mem[2][3][2] ), .ip2(n8967), .s(n9933), .op(
        n3611) );
  mux2_1 U9448 ( .ip1(\ANSWER/mem[2][4][2] ), .ip2(n8967), .s(n9934), .op(
        n3610) );
  mux2_1 U9449 ( .ip1(\ANSWER/mem[2][5][2] ), .ip2(n8967), .s(n9935), .op(
        n3609) );
  mux2_1 U9450 ( .ip1(\ANSWER/mem[2][6][2] ), .ip2(n8967), .s(n9936), .op(
        n3608) );
  mux2_1 U9451 ( .ip1(\ANSWER/mem[2][7][2] ), .ip2(n8967), .s(n9937), .op(
        n3607) );
  mux2_1 U9452 ( .ip1(\ANSWER/mem[2][8][2] ), .ip2(n8967), .s(n9938), .op(
        n3606) );
  mux2_1 U9453 ( .ip1(\ANSWER/mem[2][9][2] ), .ip2(n8967), .s(n9939), .op(
        n3605) );
  mux2_1 U9454 ( .ip1(\ANSWER/mem[3][0][2] ), .ip2(n8967), .s(n9940), .op(
        n3604) );
  mux2_1 U9455 ( .ip1(\ANSWER/mem[3][1][2] ), .ip2(n8967), .s(n9941), .op(
        n3603) );
  mux2_1 U9456 ( .ip1(\ANSWER/mem[3][2][2] ), .ip2(n8967), .s(n9942), .op(
        n3602) );
  mux2_1 U9457 ( .ip1(\ANSWER/mem[3][3][2] ), .ip2(n8967), .s(n9943), .op(
        n3601) );
  mux2_1 U9458 ( .ip1(\ANSWER/mem[3][4][2] ), .ip2(n8967), .s(n9944), .op(
        n3600) );
  mux2_1 U9459 ( .ip1(\ANSWER/mem[3][5][2] ), .ip2(n8967), .s(n9945), .op(
        n3599) );
  mux2_1 U9460 ( .ip1(\ANSWER/mem[3][6][2] ), .ip2(n8968), .s(n9946), .op(
        n3598) );
  mux2_1 U9461 ( .ip1(\ANSWER/mem[3][7][2] ), .ip2(n8968), .s(n9947), .op(
        n3597) );
  mux2_1 U9462 ( .ip1(\ANSWER/mem[3][8][2] ), .ip2(n8968), .s(n9948), .op(
        n3596) );
  mux2_1 U9463 ( .ip1(\ANSWER/mem[3][9][2] ), .ip2(n8968), .s(n9949), .op(
        n3595) );
  mux2_1 U9464 ( .ip1(\ANSWER/mem[4][0][2] ), .ip2(n8968), .s(n9950), .op(
        n3594) );
  mux2_1 U9465 ( .ip1(\ANSWER/mem[4][1][2] ), .ip2(n8968), .s(n9951), .op(
        n3593) );
  mux2_1 U9466 ( .ip1(\ANSWER/mem[4][2][2] ), .ip2(n8969), .s(n9952), .op(
        n3592) );
  mux2_1 U9467 ( .ip1(\ANSWER/mem[4][3][2] ), .ip2(n8969), .s(n9953), .op(
        n3591) );
  mux2_1 U9468 ( .ip1(\ANSWER/mem[4][4][2] ), .ip2(n8969), .s(n9954), .op(
        n3590) );
  mux2_1 U9469 ( .ip1(\ANSWER/mem[4][5][2] ), .ip2(n8969), .s(n9955), .op(
        n3589) );
  mux2_1 U9470 ( .ip1(\ANSWER/mem[4][6][2] ), .ip2(n8969), .s(n9956), .op(
        n3588) );
  mux2_1 U9471 ( .ip1(\ANSWER/mem[4][7][2] ), .ip2(n8969), .s(n9957), .op(
        n3587) );
  mux2_1 U9472 ( .ip1(\ANSWER/mem[4][8][2] ), .ip2(n8969), .s(n9958), .op(
        n3586) );
  mux2_1 U9473 ( .ip1(\ANSWER/mem[4][9][2] ), .ip2(n8969), .s(n9959), .op(
        n3585) );
  mux2_1 U9474 ( .ip1(\ANSWER/mem[5][0][2] ), .ip2(n8969), .s(n9960), .op(
        n3584) );
  mux2_1 U9475 ( .ip1(\ANSWER/mem[5][1][2] ), .ip2(n8968), .s(n9961), .op(
        n3583) );
  mux2_1 U9476 ( .ip1(\ANSWER/mem[5][2][2] ), .ip2(n8969), .s(n9962), .op(
        n3582) );
  mux2_1 U9477 ( .ip1(\ANSWER/mem[5][3][2] ), .ip2(n8968), .s(n9963), .op(
        n3581) );
  mux2_1 U9478 ( .ip1(\ANSWER/mem[5][4][2] ), .ip2(n8969), .s(n9964), .op(
        n3580) );
  mux2_1 U9479 ( .ip1(\ANSWER/mem[5][5][2] ), .ip2(n8968), .s(n9965), .op(
        n3579) );
  mux2_1 U9480 ( .ip1(\ANSWER/mem[5][6][2] ), .ip2(n8968), .s(n9966), .op(
        n3578) );
  mux2_1 U9481 ( .ip1(\ANSWER/mem[5][7][2] ), .ip2(n8968), .s(n9967), .op(
        n3577) );
  mux2_1 U9482 ( .ip1(\ANSWER/mem[5][8][2] ), .ip2(n8968), .s(n9968), .op(
        n3576) );
  mux2_1 U9483 ( .ip1(\ANSWER/mem[5][9][2] ), .ip2(n8968), .s(n9969), .op(
        n3575) );
  mux2_1 U9484 ( .ip1(\ANSWER/mem[6][0][2] ), .ip2(n8968), .s(n9970), .op(
        n3574) );
  mux2_1 U9485 ( .ip1(\ANSWER/mem[6][1][2] ), .ip2(n8968), .s(n9971), .op(
        n3573) );
  mux2_1 U9486 ( .ip1(\ANSWER/mem[6][2][2] ), .ip2(n8968), .s(n9972), .op(
        n3572) );
  mux2_1 U9487 ( .ip1(\ANSWER/mem[6][3][2] ), .ip2(n8968), .s(n9973), .op(
        n3571) );
  mux2_1 U9488 ( .ip1(\ANSWER/mem[6][4][2] ), .ip2(n8968), .s(n9974), .op(
        n3570) );
  mux2_1 U9489 ( .ip1(\ANSWER/mem[6][5][2] ), .ip2(n8968), .s(n9975), .op(
        n3569) );
  mux2_1 U9490 ( .ip1(\ANSWER/mem[6][6][2] ), .ip2(n8968), .s(n9976), .op(
        n3568) );
  mux2_1 U9491 ( .ip1(\ANSWER/mem[6][7][2] ), .ip2(n8968), .s(n9977), .op(
        n3567) );
  mux2_1 U9492 ( .ip1(\ANSWER/mem[6][8][2] ), .ip2(n8968), .s(n9978), .op(
        n3566) );
  mux2_1 U9493 ( .ip1(\ANSWER/mem[6][9][2] ), .ip2(n8968), .s(n9979), .op(
        n3565) );
  mux2_1 U9494 ( .ip1(\ANSWER/mem[7][0][2] ), .ip2(n8968), .s(n9980), .op(
        n3564) );
  mux2_1 U9495 ( .ip1(\ANSWER/mem[7][1][2] ), .ip2(n8968), .s(n9981), .op(
        n3563) );
  buf_1 U9496 ( .ip(n8968), .op(n8969) );
  mux2_1 U9497 ( .ip1(\ANSWER/mem[7][2][2] ), .ip2(n8969), .s(n9983), .op(
        n3562) );
  mux2_1 U9498 ( .ip1(\ANSWER/mem[7][3][2] ), .ip2(n8969), .s(n9984), .op(
        n3561) );
  mux2_1 U9499 ( .ip1(\ANSWER/mem[7][4][2] ), .ip2(n8969), .s(n9985), .op(
        n3560) );
  mux2_1 U9500 ( .ip1(\ANSWER/mem[7][5][2] ), .ip2(n8969), .s(n9986), .op(
        n3559) );
  mux2_1 U9501 ( .ip1(\ANSWER/mem[7][6][2] ), .ip2(n8969), .s(n9987), .op(
        n3558) );
  mux2_1 U9502 ( .ip1(\ANSWER/mem[7][7][2] ), .ip2(n8969), .s(n9988), .op(
        n3557) );
  mux2_1 U9503 ( .ip1(\ANSWER/mem[7][8][2] ), .ip2(n8969), .s(n9989), .op(
        n3556) );
  mux2_1 U9504 ( .ip1(\ANSWER/mem[7][9][2] ), .ip2(n8968), .s(n9990), .op(
        n3555) );
  mux2_1 U9505 ( .ip1(\ANSWER/mem[8][0][2] ), .ip2(n8969), .s(n9991), .op(
        n3554) );
  mux2_1 U9506 ( .ip1(\ANSWER/mem[8][1][2] ), .ip2(n8969), .s(n9992), .op(
        n3553) );
  mux2_1 U9507 ( .ip1(\ANSWER/mem[8][2][2] ), .ip2(n8969), .s(n9993), .op(
        n3552) );
  mux2_1 U9508 ( .ip1(\ANSWER/mem[8][3][2] ), .ip2(n8969), .s(n9994), .op(
        n3551) );
  mux2_1 U9509 ( .ip1(\ANSWER/mem[8][4][2] ), .ip2(n8968), .s(n9996), .op(
        n3550) );
  mux2_1 U9510 ( .ip1(\ANSWER/mem[8][5][2] ), .ip2(n8968), .s(n9997), .op(
        n3549) );
  mux2_1 U9511 ( .ip1(\ANSWER/mem[8][6][2] ), .ip2(n8968), .s(n9998), .op(
        n3548) );
  mux2_1 U9512 ( .ip1(\ANSWER/mem[8][7][2] ), .ip2(n8968), .s(n9999), .op(
        n3547) );
  mux2_1 U9513 ( .ip1(\ANSWER/mem[8][8][2] ), .ip2(n8968), .s(n10000), .op(
        n3546) );
  mux2_1 U9514 ( .ip1(\ANSWER/mem[8][9][2] ), .ip2(n8968), .s(n10001), .op(
        n3545) );
  mux2_1 U9515 ( .ip1(\ANSWER/mem[9][0][2] ), .ip2(n8968), .s(n10002), .op(
        n3544) );
  mux2_1 U9516 ( .ip1(\ANSWER/mem[9][1][2] ), .ip2(n8968), .s(n10003), .op(
        n3543) );
  mux2_1 U9517 ( .ip1(\ANSWER/mem[9][2][2] ), .ip2(n8968), .s(n10004), .op(
        n3542) );
  mux2_1 U9518 ( .ip1(\ANSWER/mem[9][3][2] ), .ip2(n8968), .s(n10005), .op(
        n3541) );
  mux2_1 U9519 ( .ip1(\ANSWER/mem[9][4][2] ), .ip2(n8968), .s(n10006), .op(
        n3540) );
  mux2_1 U9520 ( .ip1(\ANSWER/mem[9][5][2] ), .ip2(n8968), .s(n10007), .op(
        n3539) );
  mux2_1 U9521 ( .ip1(\ANSWER/mem[9][6][2] ), .ip2(n8969), .s(n10008), .op(
        n3538) );
  mux2_1 U9522 ( .ip1(\ANSWER/mem[9][7][2] ), .ip2(n8969), .s(n10009), .op(
        n3537) );
  mux2_1 U9523 ( .ip1(\ANSWER/mem[9][8][2] ), .ip2(n8969), .s(n10010), .op(
        n3536) );
  mux2_1 U9524 ( .ip1(\ANSWER/mem[9][9][2] ), .ip2(n8969), .s(n10011), .op(
        n3535) );
  inv_1 U9525 ( .ip(q_w2[11]), .op(n9791) );
  nor4_1 U9526 ( .ip1(n9530), .ip2(n9335), .ip3(n9788), .ip4(n9791), .op(n9082) );
  inv_1 U9527 ( .ip(n9082), .op(n8972) );
  nand2_1 U9528 ( .ip1(m2DataIn[0]), .ip2(q_w2[11]), .op(n9252) );
  nand2_1 U9529 ( .ip1(n9252), .ip2(n8970), .op(n8971) );
  nand2_1 U9530 ( .ip1(n8972), .ip2(n8971), .op(n8973) );
  inv_1 U9531 ( .ip(m2DataIn[11]), .op(n9735) );
  nor3_1 U9532 ( .ip1(n9735), .ip2(n9141), .ip3(n8973), .op(n9081) );
  or2_1 U9533 ( .ip1(n8973), .ip2(n9081), .op(n8976) );
  nand2_1 U9534 ( .ip1(m2DataIn[11]), .ip2(q_w2[0]), .op(n8974) );
  or2_1 U9535 ( .ip1(n8974), .ip2(n9081), .op(n8975) );
  nand2_1 U9536 ( .ip1(n8976), .ip2(n8975), .op(n9087) );
  nand2_1 U9537 ( .ip1(m2DataIn[4]), .ip2(q_w2[7]), .op(n9044) );
  nand4_1 U9538 ( .ip1(m2DataIn[5]), .ip2(m2DataIn[4]), .ip3(q_w2[6]), .ip4(
        q_w2[7]), .op(n9054) );
  inv_1 U9539 ( .ip(n9054), .op(n8977) );
  or2_1 U9540 ( .ip1(n9044), .ip2(n8977), .op(n8980) );
  or2_1 U9541 ( .ip1(n8978), .ip2(n8977), .op(n8979) );
  nand2_1 U9542 ( .ip1(n8980), .ip2(n8979), .op(n9052) );
  nor2_1 U9543 ( .ip1(n9792), .ip2(n9334), .op(n8981) );
  xor2_1 U9544 ( .ip1(n9052), .ip2(n8981), .op(n9086) );
  nor4_1 U9545 ( .ip1(n9467), .ip2(n9725), .ip3(n9638), .ip4(n9703), .op(n9084) );
  inv_1 U9546 ( .ip(n9084), .op(n8984) );
  nand2_1 U9547 ( .ip1(m2DataIn[6]), .ip2(q_w2[5]), .op(n9048) );
  nand2_1 U9548 ( .ip1(n9048), .ip2(n8982), .op(n8983) );
  nand2_1 U9549 ( .ip1(n8984), .ip2(n8983), .op(n8985) );
  nor3_1 U9550 ( .ip1(n9790), .ip2(n9499), .ip3(n8985), .op(n9083) );
  or2_1 U9551 ( .ip1(n8985), .ip2(n9083), .op(n8988) );
  nand2_1 U9552 ( .ip1(m2DataIn[9]), .ip2(q_w2[2]), .op(n8986) );
  or2_1 U9553 ( .ip1(n8986), .ip2(n9083), .op(n8987) );
  nand2_1 U9554 ( .ip1(n8988), .ip2(n8987), .op(n9085) );
  inv_1 U9555 ( .ip(n8989), .op(n9094) );
  or2_1 U9556 ( .ip1(n8990), .ip2(n8991), .op(n8994) );
  or2_1 U9557 ( .ip1(n8992), .ip2(n8991), .op(n8993) );
  nand2_1 U9558 ( .ip1(n8994), .ip2(n8993), .op(n9091) );
  nand2_1 U9559 ( .ip1(m2DataIn[1]), .ip2(q_w2[10]), .op(n9076) );
  nand4_1 U9560 ( .ip1(m2DataIn[2]), .ip2(m2DataIn[1]), .ip3(q_w2[9]), .ip4(
        q_w2[10]), .op(n9066) );
  inv_1 U9561 ( .ip(n9066), .op(n8995) );
  or2_1 U9562 ( .ip1(n9076), .ip2(n8995), .op(n8998) );
  or2_1 U9563 ( .ip1(n8996), .ip2(n8995), .op(n8997) );
  nand2_1 U9564 ( .ip1(n8998), .ip2(n8997), .op(n9064) );
  mux2_1 U9565 ( .ip1(n8999), .ip2(rdata[3]), .s(n9064), .op(n9090) );
  or2_1 U9566 ( .ip1(n9000), .ip2(n9001), .op(n9004) );
  or2_1 U9567 ( .ip1(n9002), .ip2(n9001), .op(n9003) );
  nand2_1 U9568 ( .ip1(n9004), .ip2(n9003), .op(n9089) );
  fulladder U9569 ( .a(n9007), .b(n9006), .ci(n9005), .co(n9092), .s(n8955) );
  nand2_1 U9570 ( .ip1(m2DataIn[8]), .ip2(q_w2[3]), .op(n9072) );
  or2_1 U9571 ( .ip1(rdata[2]), .ip2(n9008), .op(n9011) );
  or2_1 U9572 ( .ip1(n9009), .ip2(n9008), .op(n9010) );
  nand2_1 U9573 ( .ip1(n9011), .ip2(n9010), .op(n9071) );
  or2_1 U9574 ( .ip1(n9012), .ip2(n9013), .op(n9016) );
  or2_1 U9575 ( .ip1(n9014), .ip2(n9013), .op(n9015) );
  nand2_1 U9576 ( .ip1(n9016), .ip2(n9015), .op(n9070) );
  fulladder U9577 ( .a(n9019), .b(n9018), .ci(n9017), .co(n9020), .s(n8923) );
  inv_1 U9578 ( .ip(n9020), .op(n9074) );
  fulladder U9579 ( .a(n9023), .b(n9022), .ci(n9021), .co(n9073), .s(n9025) );
  fulladder U9580 ( .a(n9026), .b(n9025), .ci(n9024), .co(n9041), .s(n8942) );
  inv_1 U9581 ( .ip(n9027), .op(n9098) );
  or2_1 U9582 ( .ip1(n9029), .ip2(n9028), .op(n9031) );
  nand2_1 U9583 ( .ip1(n9031), .ip2(n9030), .op(n9097) );
  fulladder U9584 ( .a(n9034), .b(n9033), .ci(n9032), .co(n9096), .s(n8959) );
  nor3_1 U9585 ( .ip1(\SIGMOID/lut_out [2]), .ip2(\SIGMOID/lut_out [1]), .ip3(
        \SIGMOID/N64 ), .op(n9035) );
  nor2_1 U9586 ( .ip1(\SIGMOID/sign_bit ), .ip2(n9035), .op(n9036) );
  xor2_1 U9587 ( .ip1(\SIGMOID/lut_out [3]), .ip2(n9036), .op(n10296) );
  mux2_1 U9588 ( .ip1(n9037), .ip2(n10296), .s(n9907), .op(n9038) );
  buf_1 U9589 ( .ip(n9038), .op(n9039) );
  mux2_1 U9590 ( .ip1(\ANSWER/mem[0][0][3] ), .ip2(n9039), .s(n9910), .op(
        n3534) );
  mux2_1 U9591 ( .ip1(\ANSWER/mem[0][1][3] ), .ip2(n9039), .s(n9911), .op(
        n3533) );
  mux2_1 U9592 ( .ip1(\ANSWER/mem[0][2][3] ), .ip2(n9039), .s(n9912), .op(
        n3532) );
  mux2_1 U9593 ( .ip1(\ANSWER/mem[0][3][3] ), .ip2(n9039), .s(n9913), .op(
        n3531) );
  mux2_1 U9594 ( .ip1(\ANSWER/mem[0][4][3] ), .ip2(n9039), .s(n9914), .op(
        n3530) );
  mux2_1 U9595 ( .ip1(\ANSWER/mem[0][5][3] ), .ip2(n9039), .s(n9915), .op(
        n3529) );
  mux2_1 U9596 ( .ip1(\ANSWER/mem[0][6][3] ), .ip2(n9039), .s(n9916), .op(
        n3528) );
  mux2_1 U9597 ( .ip1(\ANSWER/mem[0][7][3] ), .ip2(n9039), .s(n9917), .op(
        n3527) );
  mux2_1 U9598 ( .ip1(\ANSWER/mem[0][8][3] ), .ip2(n9039), .s(n9918), .op(
        n3526) );
  mux2_1 U9599 ( .ip1(\ANSWER/mem[0][9][3] ), .ip2(n9039), .s(n9919), .op(
        n3525) );
  mux2_1 U9600 ( .ip1(\ANSWER/mem[1][0][3] ), .ip2(n9039), .s(n9920), .op(
        n3524) );
  mux2_1 U9601 ( .ip1(\ANSWER/mem[1][1][3] ), .ip2(n9039), .s(n9921), .op(
        n3523) );
  mux2_1 U9602 ( .ip1(\ANSWER/mem[1][2][3] ), .ip2(n9039), .s(n9922), .op(
        n3522) );
  buf_1 U9603 ( .ip(n9038), .op(n9040) );
  mux2_1 U9604 ( .ip1(\ANSWER/mem[1][3][3] ), .ip2(n9040), .s(n9923), .op(
        n3521) );
  mux2_1 U9605 ( .ip1(\ANSWER/mem[1][4][3] ), .ip2(n9040), .s(n9924), .op(
        n3520) );
  mux2_1 U9606 ( .ip1(\ANSWER/mem[1][5][3] ), .ip2(n9040), .s(n9925), .op(
        n3519) );
  mux2_1 U9607 ( .ip1(\ANSWER/mem[1][6][3] ), .ip2(n9040), .s(n9926), .op(
        n3518) );
  mux2_1 U9608 ( .ip1(\ANSWER/mem[1][7][3] ), .ip2(n9040), .s(n9927), .op(
        n3517) );
  mux2_1 U9609 ( .ip1(\ANSWER/mem[1][8][3] ), .ip2(n9040), .s(n9928), .op(
        n3516) );
  mux2_1 U9610 ( .ip1(\ANSWER/mem[1][9][3] ), .ip2(n9039), .s(n9929), .op(
        n3515) );
  mux2_1 U9611 ( .ip1(\ANSWER/mem[2][0][3] ), .ip2(n9040), .s(n9930), .op(
        n3514) );
  mux2_1 U9612 ( .ip1(\ANSWER/mem[2][1][3] ), .ip2(n9039), .s(n9931), .op(
        n3513) );
  mux2_1 U9613 ( .ip1(\ANSWER/mem[2][2][3] ), .ip2(n9040), .s(n9932), .op(
        n3512) );
  mux2_1 U9614 ( .ip1(\ANSWER/mem[2][3][3] ), .ip2(n9040), .s(n9933), .op(
        n3511) );
  mux2_1 U9615 ( .ip1(\ANSWER/mem[2][4][3] ), .ip2(n9039), .s(n9934), .op(
        n3510) );
  mux2_1 U9616 ( .ip1(\ANSWER/mem[2][5][3] ), .ip2(n9040), .s(n9935), .op(
        n3509) );
  mux2_1 U9617 ( .ip1(\ANSWER/mem[2][6][3] ), .ip2(n9038), .s(n9936), .op(
        n3508) );
  mux2_1 U9618 ( .ip1(\ANSWER/mem[2][7][3] ), .ip2(n9039), .s(n9937), .op(
        n3507) );
  mux2_1 U9619 ( .ip1(\ANSWER/mem[2][8][3] ), .ip2(n9038), .s(n9938), .op(
        n3506) );
  mux2_1 U9620 ( .ip1(\ANSWER/mem[2][9][3] ), .ip2(n9038), .s(n9939), .op(
        n3505) );
  mux2_1 U9621 ( .ip1(\ANSWER/mem[3][0][3] ), .ip2(n9038), .s(n9940), .op(
        n3504) );
  mux2_1 U9622 ( .ip1(\ANSWER/mem[3][1][3] ), .ip2(n9038), .s(n9941), .op(
        n3503) );
  mux2_1 U9623 ( .ip1(\ANSWER/mem[3][2][3] ), .ip2(n9040), .s(n9942), .op(
        n3502) );
  mux2_1 U9624 ( .ip1(\ANSWER/mem[3][3][3] ), .ip2(n9039), .s(n9943), .op(
        n3501) );
  mux2_1 U9625 ( .ip1(\ANSWER/mem[3][4][3] ), .ip2(n9038), .s(n9944), .op(
        n3500) );
  mux2_1 U9626 ( .ip1(\ANSWER/mem[3][5][3] ), .ip2(n9039), .s(n9945), .op(
        n3499) );
  mux2_1 U9627 ( .ip1(\ANSWER/mem[3][6][3] ), .ip2(n9040), .s(n9946), .op(
        n3498) );
  mux2_1 U9628 ( .ip1(\ANSWER/mem[3][7][3] ), .ip2(n9039), .s(n9947), .op(
        n3497) );
  mux2_1 U9629 ( .ip1(\ANSWER/mem[3][8][3] ), .ip2(n9038), .s(n9948), .op(
        n3496) );
  mux2_1 U9630 ( .ip1(\ANSWER/mem[3][9][3] ), .ip2(n9038), .s(n9949), .op(
        n3495) );
  mux2_1 U9631 ( .ip1(\ANSWER/mem[4][0][3] ), .ip2(n9038), .s(n9950), .op(
        n3494) );
  mux2_1 U9632 ( .ip1(\ANSWER/mem[4][1][3] ), .ip2(n9038), .s(n9951), .op(
        n3493) );
  mux2_1 U9633 ( .ip1(\ANSWER/mem[4][2][3] ), .ip2(n9038), .s(n9952), .op(
        n3492) );
  mux2_1 U9634 ( .ip1(\ANSWER/mem[4][3][3] ), .ip2(n9038), .s(n9953), .op(
        n3491) );
  mux2_1 U9635 ( .ip1(\ANSWER/mem[4][4][3] ), .ip2(n9040), .s(n9954), .op(
        n3490) );
  mux2_1 U9636 ( .ip1(\ANSWER/mem[4][5][3] ), .ip2(n9039), .s(n9955), .op(
        n3489) );
  mux2_1 U9637 ( .ip1(\ANSWER/mem[4][6][3] ), .ip2(n9040), .s(n9956), .op(
        n3488) );
  mux2_1 U9638 ( .ip1(\ANSWER/mem[4][7][3] ), .ip2(n9040), .s(n9957), .op(
        n3487) );
  mux2_1 U9639 ( .ip1(\ANSWER/mem[4][8][3] ), .ip2(n9038), .s(n9958), .op(
        n3486) );
  mux2_1 U9640 ( .ip1(\ANSWER/mem[4][9][3] ), .ip2(n9038), .s(n9959), .op(
        n3485) );
  mux2_1 U9641 ( .ip1(\ANSWER/mem[5][0][3] ), .ip2(n9038), .s(n9960), .op(
        n3484) );
  mux2_1 U9642 ( .ip1(\ANSWER/mem[5][1][3] ), .ip2(n9038), .s(n9961), .op(
        n3483) );
  mux2_1 U9643 ( .ip1(\ANSWER/mem[5][2][3] ), .ip2(n9038), .s(n9962), .op(
        n3482) );
  mux2_1 U9644 ( .ip1(\ANSWER/mem[5][3][3] ), .ip2(n9040), .s(n9963), .op(
        n3481) );
  mux2_1 U9645 ( .ip1(\ANSWER/mem[5][4][3] ), .ip2(n9038), .s(n9964), .op(
        n3480) );
  mux2_1 U9646 ( .ip1(\ANSWER/mem[5][5][3] ), .ip2(n9038), .s(n9965), .op(
        n3479) );
  mux2_1 U9647 ( .ip1(\ANSWER/mem[5][6][3] ), .ip2(n9038), .s(n9966), .op(
        n3478) );
  mux2_1 U9648 ( .ip1(\ANSWER/mem[5][7][3] ), .ip2(n9038), .s(n9967), .op(
        n3477) );
  mux2_1 U9649 ( .ip1(\ANSWER/mem[5][8][3] ), .ip2(n9038), .s(n9968), .op(
        n3476) );
  mux2_1 U9650 ( .ip1(\ANSWER/mem[5][9][3] ), .ip2(n9038), .s(n9969), .op(
        n3475) );
  mux2_1 U9651 ( .ip1(\ANSWER/mem[6][0][3] ), .ip2(n9038), .s(n9970), .op(
        n3474) );
  mux2_1 U9652 ( .ip1(\ANSWER/mem[6][1][3] ), .ip2(n9040), .s(n9971), .op(
        n3473) );
  mux2_1 U9653 ( .ip1(\ANSWER/mem[6][2][3] ), .ip2(n9040), .s(n9972), .op(
        n3472) );
  mux2_1 U9654 ( .ip1(\ANSWER/mem[6][3][3] ), .ip2(n9039), .s(n9973), .op(
        n3471) );
  mux2_1 U9655 ( .ip1(\ANSWER/mem[6][4][3] ), .ip2(n9040), .s(n9974), .op(
        n3470) );
  mux2_1 U9656 ( .ip1(\ANSWER/mem[6][5][3] ), .ip2(n9040), .s(n9975), .op(
        n3469) );
  mux2_1 U9657 ( .ip1(\ANSWER/mem[6][6][3] ), .ip2(n9039), .s(n9976), .op(
        n3468) );
  mux2_1 U9658 ( .ip1(\ANSWER/mem[6][7][3] ), .ip2(n9039), .s(n9977), .op(
        n3467) );
  mux2_1 U9659 ( .ip1(\ANSWER/mem[6][8][3] ), .ip2(n9038), .s(n9978), .op(
        n3466) );
  mux2_1 U9660 ( .ip1(\ANSWER/mem[6][9][3] ), .ip2(n9039), .s(n9979), .op(
        n3465) );
  mux2_1 U9661 ( .ip1(\ANSWER/mem[7][0][3] ), .ip2(n9038), .s(n9980), .op(
        n3464) );
  mux2_1 U9662 ( .ip1(\ANSWER/mem[7][1][3] ), .ip2(n9038), .s(n9981), .op(
        n3463) );
  mux2_1 U9663 ( .ip1(\ANSWER/mem[7][2][3] ), .ip2(n9038), .s(n9983), .op(
        n3462) );
  mux2_1 U9664 ( .ip1(\ANSWER/mem[7][3][3] ), .ip2(n9038), .s(n9984), .op(
        n3461) );
  mux2_1 U9665 ( .ip1(\ANSWER/mem[7][4][3] ), .ip2(n9038), .s(n9985), .op(
        n3460) );
  mux2_1 U9666 ( .ip1(\ANSWER/mem[7][5][3] ), .ip2(n9038), .s(n9986), .op(
        n3459) );
  mux2_1 U9667 ( .ip1(\ANSWER/mem[7][6][3] ), .ip2(n9038), .s(n9987), .op(
        n3458) );
  mux2_1 U9668 ( .ip1(\ANSWER/mem[7][7][3] ), .ip2(n9038), .s(n9988), .op(
        n3457) );
  mux2_1 U9669 ( .ip1(\ANSWER/mem[7][8][3] ), .ip2(n9038), .s(n9989), .op(
        n3456) );
  mux2_1 U9670 ( .ip1(\ANSWER/mem[7][9][3] ), .ip2(n9038), .s(n9990), .op(
        n3455) );
  mux2_1 U9671 ( .ip1(\ANSWER/mem[8][0][3] ), .ip2(n9038), .s(n9991), .op(
        n3454) );
  mux2_1 U9672 ( .ip1(\ANSWER/mem[8][1][3] ), .ip2(n9038), .s(n9992), .op(
        n3453) );
  mux2_1 U9673 ( .ip1(\ANSWER/mem[8][2][3] ), .ip2(n9038), .s(n9993), .op(
        n3452) );
  mux2_1 U9674 ( .ip1(\ANSWER/mem[8][3][3] ), .ip2(n9038), .s(n9994), .op(
        n3451) );
  mux2_1 U9675 ( .ip1(\ANSWER/mem[8][4][3] ), .ip2(n9039), .s(n9996), .op(
        n3450) );
  mux2_1 U9676 ( .ip1(\ANSWER/mem[8][5][3] ), .ip2(n9040), .s(n9997), .op(
        n3449) );
  mux2_1 U9677 ( .ip1(\ANSWER/mem[8][6][3] ), .ip2(n9039), .s(n9998), .op(
        n3448) );
  mux2_1 U9678 ( .ip1(\ANSWER/mem[8][7][3] ), .ip2(n9040), .s(n9999), .op(
        n3447) );
  mux2_1 U9679 ( .ip1(\ANSWER/mem[8][8][3] ), .ip2(n9040), .s(n10000), .op(
        n3446) );
  mux2_1 U9680 ( .ip1(\ANSWER/mem[8][9][3] ), .ip2(n9039), .s(n10001), .op(
        n3445) );
  mux2_1 U9681 ( .ip1(\ANSWER/mem[9][0][3] ), .ip2(n9039), .s(n10002), .op(
        n3444) );
  mux2_1 U9682 ( .ip1(\ANSWER/mem[9][1][3] ), .ip2(n9040), .s(n10003), .op(
        n3443) );
  mux2_1 U9683 ( .ip1(\ANSWER/mem[9][2][3] ), .ip2(n9039), .s(n10004), .op(
        n3442) );
  mux2_1 U9684 ( .ip1(\ANSWER/mem[9][3][3] ), .ip2(n9039), .s(n10005), .op(
        n3441) );
  mux2_1 U9685 ( .ip1(\ANSWER/mem[9][4][3] ), .ip2(n9040), .s(n10006), .op(
        n3440) );
  mux2_1 U9686 ( .ip1(\ANSWER/mem[9][5][3] ), .ip2(n9039), .s(n10007), .op(
        n3439) );
  mux2_1 U9687 ( .ip1(\ANSWER/mem[9][6][3] ), .ip2(n9040), .s(n10008), .op(
        n3438) );
  mux2_1 U9688 ( .ip1(\ANSWER/mem[9][7][3] ), .ip2(n9040), .s(n10009), .op(
        n3437) );
  mux2_1 U9689 ( .ip1(\ANSWER/mem[9][8][3] ), .ip2(n9040), .s(n10010), .op(
        n3436) );
  mux2_1 U9690 ( .ip1(\ANSWER/mem[9][9][3] ), .ip2(n9040), .s(n10011), .op(
        n3435) );
  fulladder U9691 ( .a(n9043), .b(n9042), .ci(n9041), .co(n9112), .s(n9027) );
  inv_1 U9692 ( .ip(n9112), .op(n9102) );
  nand2_1 U9693 ( .ip1(m2DataIn[5]), .ip2(q_w2[7]), .op(n9045) );
  nor3_1 U9694 ( .ip1(n9702), .ip2(n9788), .ip3(n9044), .op(n9156) );
  or2_1 U9695 ( .ip1(n9045), .ip2(n9156), .op(n9047) );
  nand2_1 U9696 ( .ip1(m2DataIn[4]), .ip2(q_w2[8]), .op(n9132) );
  or2_1 U9697 ( .ip1(n9132), .ip2(n9156), .op(n9046) );
  nand2_1 U9698 ( .ip1(n9047), .ip2(n9046), .op(n9155) );
  nor2_1 U9699 ( .ip1(n9735), .ip2(n9334), .op(n9157) );
  xor2_1 U9700 ( .ip1(n9155), .ip2(n9157), .op(n9124) );
  nand2_1 U9701 ( .ip1(m2DataIn[7]), .ip2(q_w2[5]), .op(n9049) );
  nor3_1 U9702 ( .ip1(n9725), .ip2(n9732), .ip3(n9048), .op(n9162) );
  or2_1 U9703 ( .ip1(n9049), .ip2(n9162), .op(n9051) );
  nand2_1 U9704 ( .ip1(m2DataIn[6]), .ip2(q_w2[6]), .op(n9142) );
  or2_1 U9705 ( .ip1(n9142), .ip2(n9162), .op(n9050) );
  nand2_1 U9706 ( .ip1(n9051), .ip2(n9050), .op(n9161) );
  nor2_1 U9707 ( .ip1(n9792), .ip2(n9499), .op(n9163) );
  xor2_1 U9708 ( .ip1(n9161), .ip2(n9163), .op(n9123) );
  nand3_1 U9709 ( .ip1(m2DataIn[10]), .ip2(q_w2[1]), .ip3(n9052), .op(n9053)
         );
  nand2_1 U9710 ( .ip1(n9054), .ip2(n9053), .op(n9122) );
  inv_1 U9711 ( .ip(n9055), .op(n9180) );
  nand2_1 U9712 ( .ip1(m2DataIn[3]), .ip2(q_w2[12]), .op(n9392) );
  nor3_1 U9713 ( .ip1(n9335), .ip2(n9864), .ip3(n9392), .op(n9154) );
  or2_1 U9714 ( .ip1(q_w2[12]), .ip2(n9056), .op(n9058) );
  or2_1 U9715 ( .ip1(m2DataIn[0]), .ip2(n9056), .op(n9057) );
  nand2_1 U9716 ( .ip1(n9058), .ip2(n9057), .op(n9152) );
  nor2_1 U9717 ( .ip1(n9154), .ip2(n9152), .op(n9059) );
  nand2_1 U9718 ( .ip1(m2DataIn[12]), .ip2(q_w2[0]), .op(n9151) );
  xor2_1 U9719 ( .ip1(n9059), .ip2(n9151), .op(n9128) );
  nand2_1 U9720 ( .ip1(m2DataIn[8]), .ip2(q_w2[4]), .op(n9147) );
  nand4_1 U9721 ( .ip1(m2DataIn[9]), .ip2(m2DataIn[8]), .ip3(q_w2[3]), .ip4(
        q_w2[4]), .op(n9121) );
  inv_1 U9722 ( .ip(n9121), .op(n9060) );
  or2_1 U9723 ( .ip1(n9147), .ip2(n9060), .op(n9063) );
  nand2_1 U9724 ( .ip1(m2DataIn[9]), .ip2(q_w2[3]), .op(n9061) );
  or2_1 U9725 ( .ip1(n9061), .ip2(n9060), .op(n9062) );
  nand2_1 U9726 ( .ip1(n9063), .ip2(n9062), .op(n9068) );
  nand2_1 U9727 ( .ip1(rdata[3]), .ip2(n9064), .op(n9065) );
  nand2_1 U9728 ( .ip1(n9066), .ip2(n9065), .op(n9067) );
  nand2_1 U9729 ( .ip1(n9068), .ip2(n9067), .op(n9120) );
  or2_1 U9730 ( .ip1(n9068), .ip2(n9067), .op(n9069) );
  nand2_1 U9731 ( .ip1(n9120), .ip2(n9069), .op(n9127) );
  fulladder U9732 ( .a(n9072), .b(n9071), .ci(n9070), .co(n9126), .s(n9075) );
  fulladder U9733 ( .a(n9075), .b(n9074), .ci(n9073), .co(n9178), .s(n9042) );
  inv_1 U9734 ( .ip(rdata[4]), .op(n9080) );
  nand2_1 U9735 ( .ip1(m2DataIn[2]), .ip2(q_w2[10]), .op(n9077) );
  nor3_1 U9736 ( .ip1(n9500), .ip2(n9791), .ip3(n9076), .op(n9172) );
  or2_1 U9737 ( .ip1(n9077), .ip2(n9172), .op(n9079) );
  nand2_1 U9738 ( .ip1(m2DataIn[1]), .ip2(q_w2[11]), .op(n9166) );
  or2_1 U9739 ( .ip1(n9166), .ip2(n9172), .op(n9078) );
  nand2_1 U9740 ( .ip1(n9079), .ip2(n9078), .op(n9173) );
  mux2_1 U9741 ( .ip1(n9080), .ip2(rdata[4]), .s(n9173), .op(n9118) );
  nor2_1 U9742 ( .ip1(n9082), .ip2(n9081), .op(n9117) );
  nor2_1 U9743 ( .ip1(n9084), .ip2(n9083), .op(n9116) );
  fulladder U9744 ( .a(n9087), .b(n9086), .ci(n9085), .co(n9088), .s(n8989) );
  inv_1 U9745 ( .ip(n9088), .op(n9130) );
  fulladder U9746 ( .a(n9091), .b(n9090), .ci(n9089), .co(n9129), .s(n9093) );
  fulladder U9747 ( .a(n9094), .b(n9093), .ci(n9092), .co(n9109), .s(n9043) );
  inv_1 U9748 ( .ip(n9095), .op(n9099) );
  fulladder U9749 ( .a(n9098), .b(n9097), .ci(n9096), .co(n9100), .s(n9037) );
  and2_1 U9750 ( .ip1(n9099), .ip2(n9100), .op(n9115) );
  nor2_1 U9751 ( .ip1(n9100), .ip2(n9099), .op(n9113) );
  nor2_1 U9752 ( .ip1(n9115), .ip2(n9113), .op(n9101) );
  mux2_1 U9753 ( .ip1(n9102), .ip2(n9112), .s(n9101), .op(n9105) );
  inv_1 U9754 ( .ip(\SIGMOID/lut_out [4]), .op(n9104) );
  or4_1 U9755 ( .ip1(\SIGMOID/lut_out [3]), .ip2(\SIGMOID/lut_out [2]), .ip3(
        \SIGMOID/lut_out [1]), .ip4(\SIGMOID/N64 ), .op(n9186) );
  nand2_1 U9756 ( .ip1(n9187), .ip2(n9186), .op(n9103) );
  mux2_1 U9757 ( .ip1(n9104), .ip2(\SIGMOID/lut_out [4]), .s(n9103), .op(
        n10328) );
  mux2_1 U9758 ( .ip1(n9105), .ip2(n10328), .s(n9907), .op(n9106) );
  mux2_1 U9759 ( .ip1(\ANSWER/mem[0][0][4] ), .ip2(n9106), .s(n9910), .op(
        n3434) );
  buf_1 U9760 ( .ip(n9106), .op(n9108) );
  mux2_1 U9761 ( .ip1(\ANSWER/mem[0][1][4] ), .ip2(n9108), .s(n9911), .op(
        n3433) );
  buf_1 U9762 ( .ip(n9106), .op(n9107) );
  mux2_1 U9763 ( .ip1(\ANSWER/mem[0][2][4] ), .ip2(n9107), .s(n9912), .op(
        n3432) );
  mux2_1 U9764 ( .ip1(\ANSWER/mem[0][3][4] ), .ip2(n9108), .s(n9913), .op(
        n3431) );
  mux2_1 U9765 ( .ip1(\ANSWER/mem[0][4][4] ), .ip2(n9107), .s(n9914), .op(
        n3430) );
  mux2_1 U9766 ( .ip1(\ANSWER/mem[0][5][4] ), .ip2(n9108), .s(n9915), .op(
        n3429) );
  mux2_1 U9767 ( .ip1(\ANSWER/mem[0][6][4] ), .ip2(n9107), .s(n9916), .op(
        n3428) );
  mux2_1 U9768 ( .ip1(\ANSWER/mem[0][7][4] ), .ip2(n9108), .s(n9917), .op(
        n3427) );
  mux2_1 U9769 ( .ip1(\ANSWER/mem[0][8][4] ), .ip2(n9107), .s(n9918), .op(
        n3426) );
  mux2_1 U9770 ( .ip1(\ANSWER/mem[0][9][4] ), .ip2(n9108), .s(n9919), .op(
        n3425) );
  mux2_1 U9771 ( .ip1(\ANSWER/mem[1][0][4] ), .ip2(n9107), .s(n9920), .op(
        n3424) );
  mux2_1 U9772 ( .ip1(\ANSWER/mem[1][1][4] ), .ip2(n9108), .s(n9921), .op(
        n3423) );
  mux2_1 U9773 ( .ip1(\ANSWER/mem[1][2][4] ), .ip2(n9106), .s(n9922), .op(
        n3422) );
  mux2_1 U9774 ( .ip1(\ANSWER/mem[1][3][4] ), .ip2(n9106), .s(n9923), .op(
        n3421) );
  mux2_1 U9775 ( .ip1(\ANSWER/mem[1][4][4] ), .ip2(n9106), .s(n9924), .op(
        n3420) );
  mux2_1 U9776 ( .ip1(\ANSWER/mem[1][5][4] ), .ip2(n9106), .s(n9925), .op(
        n3419) );
  mux2_1 U9777 ( .ip1(\ANSWER/mem[1][6][4] ), .ip2(n9106), .s(n9926), .op(
        n3418) );
  mux2_1 U9778 ( .ip1(\ANSWER/mem[1][7][4] ), .ip2(n9106), .s(n9927), .op(
        n3417) );
  mux2_1 U9779 ( .ip1(\ANSWER/mem[1][8][4] ), .ip2(n9106), .s(n9928), .op(
        n3416) );
  mux2_1 U9780 ( .ip1(\ANSWER/mem[1][9][4] ), .ip2(n9106), .s(n9929), .op(
        n3415) );
  mux2_1 U9781 ( .ip1(\ANSWER/mem[2][0][4] ), .ip2(n9107), .s(n9930), .op(
        n3414) );
  mux2_1 U9782 ( .ip1(\ANSWER/mem[2][1][4] ), .ip2(n9107), .s(n9931), .op(
        n3413) );
  mux2_1 U9783 ( .ip1(\ANSWER/mem[2][2][4] ), .ip2(n9108), .s(n9932), .op(
        n3412) );
  mux2_1 U9784 ( .ip1(\ANSWER/mem[2][3][4] ), .ip2(n9108), .s(n9933), .op(
        n3411) );
  mux2_1 U9785 ( .ip1(\ANSWER/mem[2][4][4] ), .ip2(n9106), .s(n9934), .op(
        n3410) );
  mux2_1 U9786 ( .ip1(\ANSWER/mem[2][5][4] ), .ip2(n9106), .s(n9935), .op(
        n3409) );
  mux2_1 U9787 ( .ip1(\ANSWER/mem[2][6][4] ), .ip2(n9106), .s(n9936), .op(
        n3408) );
  mux2_1 U9788 ( .ip1(\ANSWER/mem[2][7][4] ), .ip2(n9106), .s(n9937), .op(
        n3407) );
  mux2_1 U9789 ( .ip1(\ANSWER/mem[2][8][4] ), .ip2(n9106), .s(n9938), .op(
        n3406) );
  mux2_1 U9790 ( .ip1(\ANSWER/mem[2][9][4] ), .ip2(n9106), .s(n9939), .op(
        n3405) );
  mux2_1 U9791 ( .ip1(\ANSWER/mem[3][0][4] ), .ip2(n9106), .s(n9940), .op(
        n3404) );
  mux2_1 U9792 ( .ip1(\ANSWER/mem[3][1][4] ), .ip2(n9106), .s(n9941), .op(
        n3403) );
  mux2_1 U9793 ( .ip1(\ANSWER/mem[3][2][4] ), .ip2(n9106), .s(n9942), .op(
        n3402) );
  mux2_1 U9794 ( .ip1(\ANSWER/mem[3][3][4] ), .ip2(n9106), .s(n9943), .op(
        n3401) );
  mux2_1 U9795 ( .ip1(\ANSWER/mem[3][4][4] ), .ip2(n9106), .s(n9944), .op(
        n3400) );
  mux2_1 U9796 ( .ip1(\ANSWER/mem[3][5][4] ), .ip2(n9106), .s(n9945), .op(
        n3399) );
  mux2_1 U9797 ( .ip1(\ANSWER/mem[3][6][4] ), .ip2(n9107), .s(n9946), .op(
        n3398) );
  mux2_1 U9798 ( .ip1(\ANSWER/mem[3][7][4] ), .ip2(n9106), .s(n9947), .op(
        n3397) );
  mux2_1 U9799 ( .ip1(\ANSWER/mem[3][8][4] ), .ip2(n9106), .s(n9948), .op(
        n3396) );
  mux2_1 U9800 ( .ip1(\ANSWER/mem[3][9][4] ), .ip2(n9106), .s(n9949), .op(
        n3395) );
  mux2_1 U9801 ( .ip1(\ANSWER/mem[4][0][4] ), .ip2(n9106), .s(n9950), .op(
        n3394) );
  mux2_1 U9802 ( .ip1(\ANSWER/mem[4][1][4] ), .ip2(n9106), .s(n9951), .op(
        n3393) );
  mux2_1 U9803 ( .ip1(\ANSWER/mem[4][2][4] ), .ip2(n9106), .s(n9952), .op(
        n3392) );
  mux2_1 U9804 ( .ip1(\ANSWER/mem[4][3][4] ), .ip2(n9106), .s(n9953), .op(
        n3391) );
  mux2_1 U9805 ( .ip1(\ANSWER/mem[4][4][4] ), .ip2(n9106), .s(n9954), .op(
        n3390) );
  mux2_1 U9806 ( .ip1(\ANSWER/mem[4][5][4] ), .ip2(n9106), .s(n9955), .op(
        n3389) );
  mux2_1 U9807 ( .ip1(\ANSWER/mem[4][6][4] ), .ip2(n9106), .s(n9956), .op(
        n3388) );
  mux2_1 U9808 ( .ip1(\ANSWER/mem[4][7][4] ), .ip2(n9106), .s(n9957), .op(
        n3387) );
  mux2_1 U9809 ( .ip1(\ANSWER/mem[4][8][4] ), .ip2(n9108), .s(n9958), .op(
        n3386) );
  mux2_1 U9810 ( .ip1(\ANSWER/mem[4][9][4] ), .ip2(n9108), .s(n9959), .op(
        n3385) );
  mux2_1 U9811 ( .ip1(\ANSWER/mem[5][0][4] ), .ip2(n9108), .s(n9960), .op(
        n3384) );
  mux2_1 U9812 ( .ip1(\ANSWER/mem[5][1][4] ), .ip2(n9108), .s(n9961), .op(
        n3383) );
  mux2_1 U9813 ( .ip1(\ANSWER/mem[5][2][4] ), .ip2(n9107), .s(n9962), .op(
        n3382) );
  mux2_1 U9814 ( .ip1(\ANSWER/mem[5][3][4] ), .ip2(n9106), .s(n9963), .op(
        n3381) );
  mux2_1 U9815 ( .ip1(\ANSWER/mem[5][4][4] ), .ip2(n9108), .s(n9964), .op(
        n3380) );
  mux2_1 U9816 ( .ip1(\ANSWER/mem[5][5][4] ), .ip2(n9107), .s(n9965), .op(
        n3379) );
  mux2_1 U9817 ( .ip1(\ANSWER/mem[5][6][4] ), .ip2(n9106), .s(n9966), .op(
        n3378) );
  mux2_1 U9818 ( .ip1(\ANSWER/mem[5][7][4] ), .ip2(n9108), .s(n9967), .op(
        n3377) );
  mux2_1 U9819 ( .ip1(\ANSWER/mem[5][8][4] ), .ip2(n9107), .s(n9968), .op(
        n3376) );
  mux2_1 U9820 ( .ip1(\ANSWER/mem[5][9][4] ), .ip2(n9106), .s(n9969), .op(
        n3375) );
  mux2_1 U9821 ( .ip1(\ANSWER/mem[6][0][4] ), .ip2(n9106), .s(n9970), .op(
        n3374) );
  mux2_1 U9822 ( .ip1(\ANSWER/mem[6][1][4] ), .ip2(n9107), .s(n9971), .op(
        n3373) );
  mux2_1 U9823 ( .ip1(\ANSWER/mem[6][2][4] ), .ip2(n9108), .s(n9972), .op(
        n3372) );
  mux2_1 U9824 ( .ip1(\ANSWER/mem[6][3][4] ), .ip2(n9107), .s(n9973), .op(
        n3371) );
  mux2_1 U9825 ( .ip1(\ANSWER/mem[6][4][4] ), .ip2(n9108), .s(n9974), .op(
        n3370) );
  mux2_1 U9826 ( .ip1(\ANSWER/mem[6][5][4] ), .ip2(n9108), .s(n9975), .op(
        n3369) );
  mux2_1 U9827 ( .ip1(\ANSWER/mem[6][6][4] ), .ip2(n9106), .s(n9976), .op(
        n3368) );
  mux2_1 U9828 ( .ip1(\ANSWER/mem[6][7][4] ), .ip2(n9108), .s(n9977), .op(
        n3367) );
  mux2_1 U9829 ( .ip1(\ANSWER/mem[6][8][4] ), .ip2(n9108), .s(n9978), .op(
        n3366) );
  mux2_1 U9830 ( .ip1(\ANSWER/mem[6][9][4] ), .ip2(n9106), .s(n9979), .op(
        n3365) );
  mux2_1 U9831 ( .ip1(\ANSWER/mem[7][0][4] ), .ip2(n9108), .s(n9980), .op(
        n3364) );
  mux2_1 U9832 ( .ip1(\ANSWER/mem[7][1][4] ), .ip2(n9108), .s(n9981), .op(
        n3363) );
  mux2_1 U9833 ( .ip1(\ANSWER/mem[7][2][4] ), .ip2(n9107), .s(n9983), .op(
        n3362) );
  mux2_1 U9834 ( .ip1(\ANSWER/mem[7][3][4] ), .ip2(n9107), .s(n9984), .op(
        n3361) );
  mux2_1 U9835 ( .ip1(\ANSWER/mem[7][4][4] ), .ip2(n9108), .s(n9985), .op(
        n3360) );
  mux2_1 U9836 ( .ip1(\ANSWER/mem[7][5][4] ), .ip2(n9108), .s(n9986), .op(
        n3359) );
  mux2_1 U9837 ( .ip1(\ANSWER/mem[7][6][4] ), .ip2(n9108), .s(n9987), .op(
        n3358) );
  mux2_1 U9838 ( .ip1(\ANSWER/mem[7][7][4] ), .ip2(n9108), .s(n9988), .op(
        n3357) );
  mux2_1 U9839 ( .ip1(\ANSWER/mem[7][8][4] ), .ip2(n9108), .s(n9989), .op(
        n3356) );
  mux2_1 U9840 ( .ip1(\ANSWER/mem[7][9][4] ), .ip2(n9107), .s(n9990), .op(
        n3355) );
  mux2_1 U9841 ( .ip1(\ANSWER/mem[8][0][4] ), .ip2(n9107), .s(n9991), .op(
        n3354) );
  mux2_1 U9842 ( .ip1(\ANSWER/mem[8][1][4] ), .ip2(n9107), .s(n9992), .op(
        n3353) );
  mux2_1 U9843 ( .ip1(\ANSWER/mem[8][2][4] ), .ip2(n9106), .s(n9993), .op(
        n3352) );
  mux2_1 U9844 ( .ip1(\ANSWER/mem[8][3][4] ), .ip2(n9108), .s(n9994), .op(
        n3351) );
  mux2_1 U9845 ( .ip1(\ANSWER/mem[8][4][4] ), .ip2(n9107), .s(n9996), .op(
        n3350) );
  mux2_1 U9846 ( .ip1(\ANSWER/mem[8][5][4] ), .ip2(n9107), .s(n9997), .op(
        n3349) );
  mux2_1 U9847 ( .ip1(\ANSWER/mem[8][6][4] ), .ip2(n9107), .s(n9998), .op(
        n3348) );
  mux2_1 U9848 ( .ip1(\ANSWER/mem[8][7][4] ), .ip2(n9107), .s(n9999), .op(
        n3347) );
  mux2_1 U9849 ( .ip1(\ANSWER/mem[8][8][4] ), .ip2(n9107), .s(n10000), .op(
        n3346) );
  mux2_1 U9850 ( .ip1(\ANSWER/mem[8][9][4] ), .ip2(n9107), .s(n10001), .op(
        n3345) );
  mux2_1 U9851 ( .ip1(\ANSWER/mem[9][0][4] ), .ip2(n9107), .s(n10002), .op(
        n3344) );
  mux2_1 U9852 ( .ip1(\ANSWER/mem[9][1][4] ), .ip2(n9107), .s(n10003), .op(
        n3343) );
  mux2_1 U9853 ( .ip1(\ANSWER/mem[9][2][4] ), .ip2(n9107), .s(n10004), .op(
        n3342) );
  mux2_1 U9854 ( .ip1(\ANSWER/mem[9][3][4] ), .ip2(n9107), .s(n10005), .op(
        n3341) );
  mux2_1 U9855 ( .ip1(\ANSWER/mem[9][4][4] ), .ip2(n9107), .s(n10006), .op(
        n3340) );
  mux2_1 U9856 ( .ip1(\ANSWER/mem[9][5][4] ), .ip2(n9107), .s(n10007), .op(
        n3339) );
  mux2_1 U9857 ( .ip1(\ANSWER/mem[9][6][4] ), .ip2(n9108), .s(n10008), .op(
        n3338) );
  mux2_1 U9858 ( .ip1(\ANSWER/mem[9][7][4] ), .ip2(n9108), .s(n10009), .op(
        n3337) );
  mux2_1 U9859 ( .ip1(\ANSWER/mem[9][8][4] ), .ip2(n9108), .s(n10010), .op(
        n3336) );
  mux2_1 U9860 ( .ip1(\ANSWER/mem[9][9][4] ), .ip2(n9108), .s(n10011), .op(
        n3335) );
  fulladder U9861 ( .a(n9111), .b(n9110), .ci(n9109), .co(n9185), .s(n9095) );
  inv_1 U9862 ( .ip(n9185), .op(n9197) );
  nor2_1 U9863 ( .ip1(n9113), .ip2(n9112), .op(n9114) );
  nor2_1 U9864 ( .ip1(n9115), .ip2(n9114), .op(n9182) );
  fulladder U9865 ( .a(n9118), .b(n9117), .ci(n9116), .co(n9119), .s(n9131) );
  inv_1 U9866 ( .ip(n9119), .op(n9233) );
  nand2_1 U9867 ( .ip1(n9121), .ip2(n9120), .op(n9232) );
  fulladder U9868 ( .a(n9124), .b(n9123), .ci(n9122), .co(n9231), .s(n9055) );
  inv_1 U9869 ( .ip(n9125), .op(n9267) );
  fulladder U9870 ( .a(n9128), .b(n9127), .ci(n9126), .co(n9266), .s(n9179) );
  fulladder U9871 ( .a(n9131), .b(n9130), .ci(n9129), .co(n9265), .s(n9110) );
  nand2_1 U9872 ( .ip1(m2DataIn[5]), .ip2(q_w2[8]), .op(n9133) );
  nor3_1 U9873 ( .ip1(n9702), .ip2(n9864), .ip3(n9132), .op(n9218) );
  or2_1 U9874 ( .ip1(n9133), .ip2(n9218), .op(n9135) );
  nand2_1 U9875 ( .ip1(m2DataIn[4]), .ip2(q_w2[9]), .op(n9330) );
  or2_1 U9876 ( .ip1(n9330), .ip2(n9218), .op(n9134) );
  nand2_1 U9877 ( .ip1(n9135), .ip2(n9134), .op(n9217) );
  nor2_1 U9878 ( .ip1(n9815), .ip2(n9334), .op(n9219) );
  xor2_1 U9879 ( .ip1(n9217), .ip2(n9219), .op(n9263) );
  nand2_1 U9880 ( .ip1(m2DataIn[3]), .ip2(q_w2[10]), .op(n9137) );
  nand2_1 U9881 ( .ip1(m2DataIn[3]), .ip2(q_w2[13]), .op(n9460) );
  nor2_1 U9882 ( .ip1(n9136), .ip2(n9460), .op(n9243) );
  or2_1 U9883 ( .ip1(n9137), .ip2(n9243), .op(n9140) );
  nand2_1 U9884 ( .ip1(m2DataIn[0]), .ip2(q_w2[13]), .op(n9138) );
  or2_1 U9885 ( .ip1(n9138), .ip2(n9243), .op(n9139) );
  nand2_1 U9886 ( .ip1(n9140), .ip2(n9139), .op(n9245) );
  nor2_1 U9887 ( .ip1(n9799), .ip2(n9141), .op(n9244) );
  xor2_1 U9888 ( .ip1(n9245), .ip2(n9244), .op(n9262) );
  nand2_1 U9889 ( .ip1(m2DataIn[7]), .ip2(q_w2[6]), .op(n9144) );
  inv_1 U9890 ( .ip(q_w2[7]), .op(n9143) );
  nor3_1 U9891 ( .ip1(n9725), .ip2(n9143), .ip3(n9142), .op(n9223) );
  or2_1 U9892 ( .ip1(n9144), .ip2(n9223), .op(n9146) );
  nand2_1 U9893 ( .ip1(m2DataIn[6]), .ip2(q_w2[7]), .op(n9566) );
  or2_1 U9894 ( .ip1(n9566), .ip2(n9223), .op(n9145) );
  nand2_1 U9895 ( .ip1(n9146), .ip2(n9145), .op(n9222) );
  nor2_1 U9896 ( .ip1(n9735), .ip2(n9499), .op(n9224) );
  xor2_1 U9897 ( .ip1(n9222), .ip2(n9224), .op(n9261) );
  nand2_1 U9898 ( .ip1(m2DataIn[9]), .ip2(q_w2[4]), .op(n9235) );
  nor3_1 U9899 ( .ip1(n9790), .ip2(n9703), .ip3(n9147), .op(n9204) );
  or2_1 U9900 ( .ip1(n9235), .ip2(n9204), .op(n9150) );
  nand2_1 U9901 ( .ip1(m2DataIn[8]), .ip2(q_w2[5]), .op(n9148) );
  or2_1 U9902 ( .ip1(n9148), .ip2(n9204), .op(n9149) );
  nand2_1 U9903 ( .ip1(n9150), .ip2(n9149), .op(n9203) );
  nor2_1 U9904 ( .ip1(n9792), .ip2(n9372), .op(n9205) );
  xnor2_1 U9905 ( .ip1(n9203), .ip2(n9205), .op(n9229) );
  nor2_1 U9906 ( .ip1(n9152), .ip2(n9151), .op(n9153) );
  nor2_1 U9907 ( .ip1(n9154), .ip2(n9153), .op(n9228) );
  or2_1 U9908 ( .ip1(n9155), .ip2(n9156), .op(n9159) );
  or2_1 U9909 ( .ip1(n9157), .ip2(n9156), .op(n9158) );
  nand2_1 U9910 ( .ip1(n9159), .ip2(n9158), .op(n9227) );
  inv_1 U9911 ( .ip(n9160), .op(n9201) );
  or2_1 U9912 ( .ip1(n9161), .ip2(n9162), .op(n9165) );
  or2_1 U9913 ( .ip1(n9163), .ip2(n9162), .op(n9164) );
  nand2_1 U9914 ( .ip1(n9165), .ip2(n9164), .op(n9259) );
  inv_1 U9915 ( .ip(rdata[5]), .op(n9171) );
  nand2_1 U9916 ( .ip1(m2DataIn[1]), .ip2(q_w2[12]), .op(n9167) );
  nand2_1 U9917 ( .ip1(m2DataIn[2]), .ip2(q_w2[12]), .op(n9213) );
  nor2_1 U9918 ( .ip1(n9213), .ip2(n9166), .op(n9208) );
  or2_1 U9919 ( .ip1(n9167), .ip2(n9208), .op(n9170) );
  nand2_1 U9920 ( .ip1(m2DataIn[2]), .ip2(q_w2[11]), .op(n9168) );
  or2_1 U9921 ( .ip1(n9168), .ip2(n9208), .op(n9169) );
  nand2_1 U9922 ( .ip1(n9170), .ip2(n9169), .op(n9209) );
  mux2_1 U9923 ( .ip1(n9171), .ip2(rdata[5]), .s(n9209), .op(n9258) );
  or2_1 U9924 ( .ip1(rdata[4]), .ip2(n9172), .op(n9175) );
  or2_1 U9925 ( .ip1(n9173), .ip2(n9172), .op(n9174) );
  nand2_1 U9926 ( .ip1(n9175), .ip2(n9174), .op(n9257) );
  inv_1 U9927 ( .ip(n9176), .op(n9200) );
  inv_1 U9928 ( .ip(n9177), .op(n9272) );
  fulladder U9929 ( .a(n9180), .b(n9179), .ci(n9178), .co(n9271), .s(n9111) );
  nor2_1 U9930 ( .ip1(n9182), .ip2(n9181), .op(n9196) );
  nand2_1 U9931 ( .ip1(n9182), .ip2(n9181), .op(n9199) );
  inv_1 U9932 ( .ip(n9199), .op(n9183) );
  nor2_1 U9933 ( .ip1(n9196), .ip2(n9183), .op(n9184) );
  mux2_1 U9934 ( .ip1(n9197), .ip2(n9185), .s(n9184), .op(n9190) );
  inv_1 U9935 ( .ip(\SIGMOID/lut_out [5]), .op(n9189) );
  or2_1 U9936 ( .ip1(\SIGMOID/lut_out [4]), .ip2(n9186), .op(n9354) );
  nand2_1 U9937 ( .ip1(n9187), .ip2(n9354), .op(n9188) );
  mux2_1 U9938 ( .ip1(n9189), .ip2(\SIGMOID/lut_out [5]), .s(n9188), .op(
        n10360) );
  mux2_1 U9939 ( .ip1(n9190), .ip2(n10360), .s(n9907), .op(n9191) );
  mux2_1 U9940 ( .ip1(\ANSWER/mem[0][0][5] ), .ip2(n9191), .s(n9910), .op(
        n3334) );
  buf_1 U9941 ( .ip(n9191), .op(n9193) );
  mux2_1 U9942 ( .ip1(\ANSWER/mem[0][1][5] ), .ip2(n9193), .s(n9911), .op(
        n3333) );
  buf_1 U9943 ( .ip(n9191), .op(n9192) );
  mux2_1 U9944 ( .ip1(\ANSWER/mem[0][2][5] ), .ip2(n9192), .s(n9912), .op(
        n3332) );
  mux2_1 U9945 ( .ip1(\ANSWER/mem[0][3][5] ), .ip2(n9193), .s(n9913), .op(
        n3331) );
  mux2_1 U9946 ( .ip1(\ANSWER/mem[0][4][5] ), .ip2(n9192), .s(n9914), .op(
        n3330) );
  mux2_1 U9947 ( .ip1(\ANSWER/mem[0][5][5] ), .ip2(n9193), .s(n9915), .op(
        n3329) );
  mux2_1 U9948 ( .ip1(\ANSWER/mem[0][6][5] ), .ip2(n9192), .s(n9916), .op(
        n3328) );
  mux2_1 U9949 ( .ip1(\ANSWER/mem[0][7][5] ), .ip2(n9193), .s(n9917), .op(
        n3327) );
  mux2_1 U9950 ( .ip1(\ANSWER/mem[0][8][5] ), .ip2(n9192), .s(n9918), .op(
        n3326) );
  mux2_1 U9951 ( .ip1(\ANSWER/mem[0][9][5] ), .ip2(n9193), .s(n9919), .op(
        n3325) );
  mux2_1 U9952 ( .ip1(\ANSWER/mem[1][0][5] ), .ip2(n9192), .s(n9920), .op(
        n3324) );
  mux2_1 U9953 ( .ip1(\ANSWER/mem[1][1][5] ), .ip2(n9193), .s(n9921), .op(
        n3323) );
  mux2_1 U9954 ( .ip1(\ANSWER/mem[1][2][5] ), .ip2(n9191), .s(n9922), .op(
        n3322) );
  mux2_1 U9955 ( .ip1(\ANSWER/mem[1][3][5] ), .ip2(n9191), .s(n9923), .op(
        n3321) );
  mux2_1 U9956 ( .ip1(\ANSWER/mem[1][4][5] ), .ip2(n9191), .s(n9924), .op(
        n3320) );
  mux2_1 U9957 ( .ip1(\ANSWER/mem[1][5][5] ), .ip2(n9191), .s(n9925), .op(
        n3319) );
  mux2_1 U9958 ( .ip1(\ANSWER/mem[1][6][5] ), .ip2(n9191), .s(n9926), .op(
        n3318) );
  mux2_1 U9959 ( .ip1(\ANSWER/mem[1][7][5] ), .ip2(n9191), .s(n9927), .op(
        n3317) );
  mux2_1 U9960 ( .ip1(\ANSWER/mem[1][8][5] ), .ip2(n9191), .s(n9928), .op(
        n3316) );
  mux2_1 U9961 ( .ip1(\ANSWER/mem[1][9][5] ), .ip2(n9191), .s(n9929), .op(
        n3315) );
  mux2_1 U9962 ( .ip1(\ANSWER/mem[2][0][5] ), .ip2(n9192), .s(n9930), .op(
        n3314) );
  mux2_1 U9963 ( .ip1(\ANSWER/mem[2][1][5] ), .ip2(n9192), .s(n9931), .op(
        n3313) );
  mux2_1 U9964 ( .ip1(\ANSWER/mem[2][2][5] ), .ip2(n9193), .s(n9932), .op(
        n3312) );
  mux2_1 U9965 ( .ip1(\ANSWER/mem[2][3][5] ), .ip2(n9193), .s(n9933), .op(
        n3311) );
  mux2_1 U9966 ( .ip1(\ANSWER/mem[2][4][5] ), .ip2(n9191), .s(n9934), .op(
        n3310) );
  mux2_1 U9967 ( .ip1(\ANSWER/mem[2][5][5] ), .ip2(n9191), .s(n9935), .op(
        n3309) );
  mux2_1 U9968 ( .ip1(\ANSWER/mem[2][6][5] ), .ip2(n9191), .s(n9936), .op(
        n3308) );
  mux2_1 U9969 ( .ip1(\ANSWER/mem[2][7][5] ), .ip2(n9191), .s(n9937), .op(
        n3307) );
  mux2_1 U9970 ( .ip1(\ANSWER/mem[2][8][5] ), .ip2(n9191), .s(n9938), .op(
        n3306) );
  mux2_1 U9971 ( .ip1(\ANSWER/mem[2][9][5] ), .ip2(n9191), .s(n9939), .op(
        n3305) );
  mux2_1 U9972 ( .ip1(\ANSWER/mem[3][0][5] ), .ip2(n9191), .s(n9940), .op(
        n3304) );
  mux2_1 U9973 ( .ip1(\ANSWER/mem[3][1][5] ), .ip2(n9191), .s(n9941), .op(
        n3303) );
  mux2_1 U9974 ( .ip1(\ANSWER/mem[3][2][5] ), .ip2(n9191), .s(n9942), .op(
        n3302) );
  mux2_1 U9975 ( .ip1(\ANSWER/mem[3][3][5] ), .ip2(n9191), .s(n9943), .op(
        n3301) );
  mux2_1 U9976 ( .ip1(\ANSWER/mem[3][4][5] ), .ip2(n9191), .s(n9944), .op(
        n3300) );
  mux2_1 U9977 ( .ip1(\ANSWER/mem[3][5][5] ), .ip2(n9191), .s(n9945), .op(
        n3299) );
  mux2_1 U9978 ( .ip1(\ANSWER/mem[3][6][5] ), .ip2(n9192), .s(n9946), .op(
        n3298) );
  mux2_1 U9979 ( .ip1(\ANSWER/mem[3][7][5] ), .ip2(n9191), .s(n9947), .op(
        n3297) );
  mux2_1 U9980 ( .ip1(\ANSWER/mem[3][8][5] ), .ip2(n9191), .s(n9948), .op(
        n3296) );
  mux2_1 U9981 ( .ip1(\ANSWER/mem[3][9][5] ), .ip2(n9191), .s(n9949), .op(
        n3295) );
  mux2_1 U9982 ( .ip1(\ANSWER/mem[4][0][5] ), .ip2(n9191), .s(n9950), .op(
        n3294) );
  mux2_1 U9983 ( .ip1(\ANSWER/mem[4][1][5] ), .ip2(n9191), .s(n9951), .op(
        n3293) );
  mux2_1 U9984 ( .ip1(\ANSWER/mem[4][2][5] ), .ip2(n9191), .s(n9952), .op(
        n3292) );
  mux2_1 U9985 ( .ip1(\ANSWER/mem[4][3][5] ), .ip2(n9191), .s(n9953), .op(
        n3291) );
  mux2_1 U9986 ( .ip1(\ANSWER/mem[4][4][5] ), .ip2(n9191), .s(n9954), .op(
        n3290) );
  mux2_1 U9987 ( .ip1(\ANSWER/mem[4][5][5] ), .ip2(n9191), .s(n9955), .op(
        n3289) );
  mux2_1 U9988 ( .ip1(\ANSWER/mem[4][6][5] ), .ip2(n9191), .s(n9956), .op(
        n3288) );
  mux2_1 U9989 ( .ip1(\ANSWER/mem[4][7][5] ), .ip2(n9191), .s(n9957), .op(
        n3287) );
  mux2_1 U9990 ( .ip1(\ANSWER/mem[4][8][5] ), .ip2(n9193), .s(n9958), .op(
        n3286) );
  mux2_1 U9991 ( .ip1(\ANSWER/mem[4][9][5] ), .ip2(n9193), .s(n9959), .op(
        n3285) );
  mux2_1 U9992 ( .ip1(\ANSWER/mem[5][0][5] ), .ip2(n9193), .s(n9960), .op(
        n3284) );
  mux2_1 U9993 ( .ip1(\ANSWER/mem[5][1][5] ), .ip2(n9193), .s(n9961), .op(
        n3283) );
  mux2_1 U9994 ( .ip1(\ANSWER/mem[5][2][5] ), .ip2(n9192), .s(n9962), .op(
        n3282) );
  mux2_1 U9995 ( .ip1(\ANSWER/mem[5][3][5] ), .ip2(n9191), .s(n9963), .op(
        n3281) );
  mux2_1 U9996 ( .ip1(\ANSWER/mem[5][4][5] ), .ip2(n9193), .s(n9964), .op(
        n3280) );
  mux2_1 U9997 ( .ip1(\ANSWER/mem[5][5][5] ), .ip2(n9192), .s(n9965), .op(
        n3279) );
  mux2_1 U9998 ( .ip1(\ANSWER/mem[5][6][5] ), .ip2(n9191), .s(n9966), .op(
        n3278) );
  mux2_1 U9999 ( .ip1(\ANSWER/mem[5][7][5] ), .ip2(n9193), .s(n9967), .op(
        n3277) );
  mux2_1 U10000 ( .ip1(\ANSWER/mem[5][8][5] ), .ip2(n9192), .s(n9968), .op(
        n3276) );
  mux2_1 U10001 ( .ip1(\ANSWER/mem[5][9][5] ), .ip2(n9191), .s(n9969), .op(
        n3275) );
  mux2_1 U10002 ( .ip1(\ANSWER/mem[6][0][5] ), .ip2(n9191), .s(n9970), .op(
        n3274) );
  mux2_1 U10003 ( .ip1(\ANSWER/mem[6][1][5] ), .ip2(n9192), .s(n9971), .op(
        n3273) );
  mux2_1 U10004 ( .ip1(\ANSWER/mem[6][2][5] ), .ip2(n9193), .s(n9972), .op(
        n3272) );
  mux2_1 U10005 ( .ip1(\ANSWER/mem[6][3][5] ), .ip2(n9191), .s(n9973), .op(
        n3271) );
  mux2_1 U10006 ( .ip1(\ANSWER/mem[6][4][5] ), .ip2(n9193), .s(n9974), .op(
        n3270) );
  mux2_1 U10007 ( .ip1(\ANSWER/mem[6][5][5] ), .ip2(n9193), .s(n9975), .op(
        n3269) );
  mux2_1 U10008 ( .ip1(\ANSWER/mem[6][6][5] ), .ip2(n9192), .s(n9976), .op(
        n3268) );
  mux2_1 U10009 ( .ip1(\ANSWER/mem[6][7][5] ), .ip2(n9193), .s(n9977), .op(
        n3267) );
  mux2_1 U10010 ( .ip1(\ANSWER/mem[6][8][5] ), .ip2(n9193), .s(n9978), .op(
        n3266) );
  mux2_1 U10011 ( .ip1(\ANSWER/mem[6][9][5] ), .ip2(n9191), .s(n9979), .op(
        n3265) );
  mux2_1 U10012 ( .ip1(\ANSWER/mem[7][0][5] ), .ip2(n9193), .s(n9980), .op(
        n3264) );
  mux2_1 U10013 ( .ip1(\ANSWER/mem[7][1][5] ), .ip2(n9193), .s(n9981), .op(
        n3263) );
  mux2_1 U10014 ( .ip1(\ANSWER/mem[7][2][5] ), .ip2(n9192), .s(n9983), .op(
        n3262) );
  mux2_1 U10015 ( .ip1(\ANSWER/mem[7][3][5] ), .ip2(n9192), .s(n9984), .op(
        n3261) );
  mux2_1 U10016 ( .ip1(\ANSWER/mem[7][4][5] ), .ip2(n9193), .s(n9985), .op(
        n3260) );
  mux2_1 U10017 ( .ip1(\ANSWER/mem[7][5][5] ), .ip2(n9193), .s(n9986), .op(
        n3259) );
  mux2_1 U10018 ( .ip1(\ANSWER/mem[7][6][5] ), .ip2(n9193), .s(n9987), .op(
        n3258) );
  mux2_1 U10019 ( .ip1(\ANSWER/mem[7][7][5] ), .ip2(n9193), .s(n9988), .op(
        n3257) );
  mux2_1 U10020 ( .ip1(\ANSWER/mem[7][8][5] ), .ip2(n9193), .s(n9989), .op(
        n3256) );
  mux2_1 U10021 ( .ip1(\ANSWER/mem[7][9][5] ), .ip2(n9192), .s(n9990), .op(
        n3255) );
  mux2_1 U10022 ( .ip1(\ANSWER/mem[8][0][5] ), .ip2(n9192), .s(n9991), .op(
        n3254) );
  mux2_1 U10023 ( .ip1(\ANSWER/mem[8][1][5] ), .ip2(n9192), .s(n9992), .op(
        n3253) );
  mux2_1 U10024 ( .ip1(\ANSWER/mem[8][2][5] ), .ip2(n9191), .s(n9993), .op(
        n3252) );
  mux2_1 U10025 ( .ip1(\ANSWER/mem[8][3][5] ), .ip2(n9193), .s(n9994), .op(
        n3251) );
  mux2_1 U10026 ( .ip1(\ANSWER/mem[8][4][5] ), .ip2(n9192), .s(n9996), .op(
        n3250) );
  mux2_1 U10027 ( .ip1(\ANSWER/mem[8][5][5] ), .ip2(n9192), .s(n9997), .op(
        n3249) );
  mux2_1 U10028 ( .ip1(\ANSWER/mem[8][6][5] ), .ip2(n9192), .s(n9998), .op(
        n3248) );
  mux2_1 U10029 ( .ip1(\ANSWER/mem[8][7][5] ), .ip2(n9192), .s(n9999), .op(
        n3247) );
  mux2_1 U10030 ( .ip1(\ANSWER/mem[8][8][5] ), .ip2(n9192), .s(n10000), .op(
        n3246) );
  mux2_1 U10031 ( .ip1(\ANSWER/mem[8][9][5] ), .ip2(n9192), .s(n10001), .op(
        n3245) );
  mux2_1 U10032 ( .ip1(\ANSWER/mem[9][0][5] ), .ip2(n9192), .s(n10002), .op(
        n3244) );
  mux2_1 U10033 ( .ip1(\ANSWER/mem[9][1][5] ), .ip2(n9192), .s(n10003), .op(
        n3243) );
  mux2_1 U10034 ( .ip1(\ANSWER/mem[9][2][5] ), .ip2(n9192), .s(n10004), .op(
        n3242) );
  mux2_1 U10035 ( .ip1(\ANSWER/mem[9][3][5] ), .ip2(n9192), .s(n10005), .op(
        n3241) );
  mux2_1 U10036 ( .ip1(\ANSWER/mem[9][4][5] ), .ip2(n9192), .s(n10006), .op(
        n3240) );
  mux2_1 U10037 ( .ip1(\ANSWER/mem[9][5][5] ), .ip2(n9192), .s(n10007), .op(
        n3239) );
  mux2_1 U10038 ( .ip1(\ANSWER/mem[9][6][5] ), .ip2(n9193), .s(n10008), .op(
        n3238) );
  mux2_1 U10039 ( .ip1(\ANSWER/mem[9][7][5] ), .ip2(n9193), .s(n10009), .op(
        n3237) );
  mux2_1 U10040 ( .ip1(\ANSWER/mem[9][8][5] ), .ip2(n9193), .s(n10010), .op(
        n3236) );
  mux2_1 U10041 ( .ip1(\ANSWER/mem[9][9][5] ), .ip2(n9193), .s(n10011), .op(
        n3235) );
  nor2_1 U10042 ( .ip1(\SIGMOID/lut_out [5]), .ip2(n9354), .op(n9194) );
  nor2_1 U10043 ( .ip1(\SIGMOID/sign_bit ), .ip2(n9194), .op(n9195) );
  xor2_1 U10044 ( .ip1(\SIGMOID/lut_out [6]), .ip2(n9195), .op(n10394) );
  or2_1 U10045 ( .ip1(n9197), .ip2(n9196), .op(n9198) );
  nand2_1 U10046 ( .ip1(n9199), .ip2(n9198), .op(n9269) );
  fulladder U10047 ( .a(n9202), .b(n9201), .ci(n9200), .co(n9344), .s(n9177)
         );
  or2_1 U10048 ( .ip1(n9203), .ip2(n9204), .op(n9207) );
  or2_1 U10049 ( .ip1(n9205), .ip2(n9204), .op(n9206) );
  nand2_1 U10050 ( .ip1(n9207), .ip2(n9206), .op(n9322) );
  nand2_1 U10051 ( .ip1(m2DataIn[11]), .ip2(q_w2[3]), .op(n9419) );
  or2_1 U10052 ( .ip1(rdata[5]), .ip2(n9208), .op(n9211) );
  or2_1 U10053 ( .ip1(n9209), .ip2(n9208), .op(n9210) );
  nand2_1 U10054 ( .ip1(n9211), .ip2(n9210), .op(n9321) );
  nand2_1 U10055 ( .ip1(m2DataIn[1]), .ip2(q_w2[13]), .op(n9283) );
  nand4_1 U10056 ( .ip1(m2DataIn[2]), .ip2(m2DataIn[1]), .ip3(q_w2[12]), .ip4(
        q_w2[13]), .op(n9315) );
  inv_1 U10057 ( .ip(n9315), .op(n9212) );
  or2_1 U10058 ( .ip1(n9283), .ip2(n9212), .op(n9215) );
  or2_1 U10059 ( .ip1(n9213), .ip2(n9212), .op(n9214) );
  nand2_1 U10060 ( .ip1(n9215), .ip2(n9214), .op(n9313) );
  mux2_1 U10061 ( .ip1(n9216), .ip2(rdata[6]), .s(n9313), .op(n9320) );
  or2_1 U10062 ( .ip1(n9217), .ip2(n9218), .op(n9221) );
  or2_1 U10063 ( .ip1(n9219), .ip2(n9218), .op(n9220) );
  nand2_1 U10064 ( .ip1(n9221), .ip2(n9220), .op(n9319) );
  or2_1 U10065 ( .ip1(n9222), .ip2(n9223), .op(n9226) );
  or2_1 U10066 ( .ip1(n9224), .ip2(n9223), .op(n9225) );
  nand2_1 U10067 ( .ip1(n9226), .ip2(n9225), .op(n9318) );
  fulladder U10068 ( .a(n9229), .b(n9228), .ci(n9227), .co(n9327), .s(n9160)
         );
  inv_1 U10069 ( .ip(n9230), .op(n9343) );
  fulladder U10070 ( .a(n9233), .b(n9232), .ci(n9231), .co(n9342), .s(n9125)
         );
  inv_1 U10071 ( .ip(n9234), .op(n9353) );
  nor3_1 U10072 ( .ip1(n9792), .ip2(n9703), .ip3(n9235), .op(n9290) );
  nor2_1 U10073 ( .ip1(n9790), .ip2(n9703), .op(n9236) );
  or2_1 U10074 ( .ip1(q_w2[4]), .ip2(n9236), .op(n9238) );
  or2_1 U10075 ( .ip1(m2DataIn[10]), .ip2(n9236), .op(n9237) );
  nand2_1 U10076 ( .ip1(n9238), .ip2(n9237), .op(n9239) );
  nor2_1 U10077 ( .ip1(n9290), .ip2(n9239), .op(n9289) );
  nor2_1 U10078 ( .ip1(n9815), .ip2(n9499), .op(n9291) );
  xor2_1 U10079 ( .ip1(n9289), .ip2(n9291), .op(n9312) );
  nand2_1 U10080 ( .ip1(m2DataIn[7]), .ip2(q_w2[7]), .op(n9295) );
  nor3_1 U10081 ( .ip1(n9725), .ip2(n9788), .ip3(n9566), .op(n9305) );
  or2_1 U10082 ( .ip1(n9295), .ip2(n9305), .op(n9242) );
  nand2_1 U10083 ( .ip1(m2DataIn[6]), .ip2(q_w2[8]), .op(n9240) );
  or2_1 U10084 ( .ip1(n9240), .ip2(n9305), .op(n9241) );
  nand2_1 U10085 ( .ip1(n9242), .ip2(n9241), .op(n9304) );
  nor2_1 U10086 ( .ip1(n9799), .ip2(n9334), .op(n9306) );
  xor2_1 U10087 ( .ip1(n9304), .ip2(n9306), .op(n9311) );
  inv_1 U10088 ( .ip(n9243), .op(n9247) );
  nand2_1 U10089 ( .ip1(n9245), .ip2(n9244), .op(n9246) );
  nand2_1 U10090 ( .ip1(n9247), .ip2(n9246), .op(n9310) );
  nor2_1 U10091 ( .ip1(n9702), .ip2(n9814), .op(n9379) );
  and3_1 U10092 ( .ip1(m2DataIn[4]), .ip2(q_w2[9]), .ip3(n9379), .op(n9303) );
  nor2_1 U10093 ( .ip1(n9702), .ip2(n9864), .op(n9248) );
  or2_1 U10094 ( .ip1(q_w2[10]), .ip2(n9248), .op(n9250) );
  or2_1 U10095 ( .ip1(m2DataIn[4]), .ip2(n9248), .op(n9249) );
  nand2_1 U10096 ( .ip1(n9250), .ip2(n9249), .op(n9301) );
  nor2_1 U10097 ( .ip1(n9303), .ip2(n9301), .op(n9251) );
  nand2_1 U10098 ( .ip1(m2DataIn[8]), .ip2(q_w2[6]), .op(n9300) );
  xor2_1 U10099 ( .ip1(n9251), .ip2(n9300), .op(n9340) );
  nand2_1 U10100 ( .ip1(m2DataIn[3]), .ip2(q_w2[14]), .op(n9571) );
  nor2_1 U10101 ( .ip1(n9252), .ip2(n9571), .op(n9282) );
  nor2_1 U10102 ( .ip1(n9530), .ip2(n9791), .op(n9253) );
  or2_1 U10103 ( .ip1(q_w2[14]), .ip2(n9253), .op(n9255) );
  or2_1 U10104 ( .ip1(m2DataIn[0]), .ip2(n9253), .op(n9254) );
  nand2_1 U10105 ( .ip1(n9255), .ip2(n9254), .op(n9280) );
  nor2_1 U10106 ( .ip1(n9282), .ip2(n9280), .op(n9256) );
  nand2_1 U10107 ( .ip1(m2DataIn[14]), .ip2(q_w2[0]), .op(n9279) );
  xor2_1 U10108 ( .ip1(n9256), .ip2(n9279), .op(n9339) );
  fulladder U10109 ( .a(n9259), .b(n9258), .ci(n9257), .co(n9338), .s(n9176)
         );
  inv_1 U10110 ( .ip(n9260), .op(n9325) );
  fulladder U10111 ( .a(n9263), .b(n9262), .ci(n9261), .co(n9324), .s(n9202)
         );
  inv_1 U10112 ( .ip(n9264), .op(n9352) );
  fulladder U10113 ( .a(n9267), .b(n9266), .ci(n9265), .co(n9351), .s(n9273)
         );
  nor2_1 U10114 ( .ip1(n9269), .ip2(n9268), .op(n9347) );
  inv_1 U10115 ( .ip(n9347), .op(n9270) );
  nand2_1 U10116 ( .ip1(n9269), .ip2(n9268), .op(n9350) );
  nand2_1 U10117 ( .ip1(n9270), .ip2(n9350), .op(n9274) );
  fulladder U10118 ( .a(n9273), .b(n9272), .ci(n9271), .co(n9346), .s(n9181)
         );
  xor2_1 U10119 ( .ip1(n9274), .ip2(n9346), .op(n9275) );
  mux2_1 U10120 ( .ip1(n10394), .ip2(n9275), .s(n9445), .op(n9277) );
  buf_1 U10121 ( .ip(n9277), .op(n9276) );
  mux2_1 U10122 ( .ip1(\ANSWER/mem[0][0][6] ), .ip2(n9276), .s(n9910), .op(
        n3234) );
  mux2_1 U10123 ( .ip1(\ANSWER/mem[0][1][6] ), .ip2(n9276), .s(n9911), .op(
        n3233) );
  mux2_1 U10124 ( .ip1(\ANSWER/mem[0][2][6] ), .ip2(n9276), .s(n9912), .op(
        n3232) );
  mux2_1 U10125 ( .ip1(\ANSWER/mem[0][3][6] ), .ip2(n9276), .s(n9913), .op(
        n3231) );
  mux2_1 U10126 ( .ip1(\ANSWER/mem[0][4][6] ), .ip2(n9276), .s(n9914), .op(
        n3230) );
  mux2_1 U10127 ( .ip1(\ANSWER/mem[0][5][6] ), .ip2(n9276), .s(n9915), .op(
        n3229) );
  mux2_1 U10128 ( .ip1(\ANSWER/mem[0][6][6] ), .ip2(n9276), .s(n9916), .op(
        n3228) );
  mux2_1 U10129 ( .ip1(\ANSWER/mem[0][7][6] ), .ip2(n9276), .s(n9917), .op(
        n3227) );
  mux2_1 U10130 ( .ip1(\ANSWER/mem[0][8][6] ), .ip2(n9276), .s(n9918), .op(
        n3226) );
  mux2_1 U10131 ( .ip1(\ANSWER/mem[0][9][6] ), .ip2(n9276), .s(n9919), .op(
        n3225) );
  mux2_1 U10132 ( .ip1(\ANSWER/mem[1][0][6] ), .ip2(n9276), .s(n9920), .op(
        n3224) );
  mux2_1 U10133 ( .ip1(\ANSWER/mem[1][1][6] ), .ip2(n9276), .s(n9921), .op(
        n3223) );
  mux2_1 U10134 ( .ip1(\ANSWER/mem[1][2][6] ), .ip2(n9277), .s(n9922), .op(
        n3222) );
  buf_1 U10135 ( .ip(n9277), .op(n9278) );
  mux2_1 U10136 ( .ip1(\ANSWER/mem[1][3][6] ), .ip2(n9278), .s(n9923), .op(
        n3221) );
  mux2_1 U10137 ( .ip1(\ANSWER/mem[1][4][6] ), .ip2(n9278), .s(n9924), .op(
        n3220) );
  mux2_1 U10138 ( .ip1(\ANSWER/mem[1][5][6] ), .ip2(n9278), .s(n9925), .op(
        n3219) );
  mux2_1 U10139 ( .ip1(\ANSWER/mem[1][6][6] ), .ip2(n9277), .s(n9926), .op(
        n3218) );
  mux2_1 U10140 ( .ip1(\ANSWER/mem[1][7][6] ), .ip2(n9277), .s(n9927), .op(
        n3217) );
  mux2_1 U10141 ( .ip1(\ANSWER/mem[1][8][6] ), .ip2(n9277), .s(n9928), .op(
        n3216) );
  mux2_1 U10142 ( .ip1(\ANSWER/mem[1][9][6] ), .ip2(n9277), .s(n9929), .op(
        n3215) );
  mux2_1 U10143 ( .ip1(\ANSWER/mem[2][0][6] ), .ip2(n9277), .s(n9930), .op(
        n3214) );
  mux2_1 U10144 ( .ip1(\ANSWER/mem[2][1][6] ), .ip2(n9277), .s(n9931), .op(
        n3213) );
  mux2_1 U10145 ( .ip1(\ANSWER/mem[2][2][6] ), .ip2(n9277), .s(n9932), .op(
        n3212) );
  mux2_1 U10146 ( .ip1(\ANSWER/mem[2][3][6] ), .ip2(n9277), .s(n9933), .op(
        n3211) );
  mux2_1 U10147 ( .ip1(\ANSWER/mem[2][4][6] ), .ip2(n9276), .s(n9934), .op(
        n3210) );
  mux2_1 U10148 ( .ip1(\ANSWER/mem[2][5][6] ), .ip2(n9277), .s(n9935), .op(
        n3209) );
  mux2_1 U10149 ( .ip1(\ANSWER/mem[2][6][6] ), .ip2(n9278), .s(n9936), .op(
        n3208) );
  mux2_1 U10150 ( .ip1(\ANSWER/mem[2][7][6] ), .ip2(n9277), .s(n9937), .op(
        n3207) );
  mux2_1 U10151 ( .ip1(\ANSWER/mem[2][8][6] ), .ip2(n9277), .s(n9938), .op(
        n3206) );
  mux2_1 U10152 ( .ip1(\ANSWER/mem[2][9][6] ), .ip2(n9277), .s(n9939), .op(
        n3205) );
  mux2_1 U10153 ( .ip1(\ANSWER/mem[3][0][6] ), .ip2(n9277), .s(n9940), .op(
        n3204) );
  mux2_1 U10154 ( .ip1(\ANSWER/mem[3][1][6] ), .ip2(n9277), .s(n9941), .op(
        n3203) );
  mux2_1 U10155 ( .ip1(\ANSWER/mem[3][2][6] ), .ip2(n9277), .s(n9942), .op(
        n3202) );
  mux2_1 U10156 ( .ip1(\ANSWER/mem[3][3][6] ), .ip2(n9278), .s(n9943), .op(
        n3201) );
  mux2_1 U10157 ( .ip1(\ANSWER/mem[3][4][6] ), .ip2(n9277), .s(n9944), .op(
        n3200) );
  mux2_1 U10158 ( .ip1(\ANSWER/mem[3][5][6] ), .ip2(n9278), .s(n9945), .op(
        n3199) );
  mux2_1 U10159 ( .ip1(\ANSWER/mem[3][6][6] ), .ip2(n9276), .s(n9946), .op(
        n3198) );
  mux2_1 U10160 ( .ip1(\ANSWER/mem[3][7][6] ), .ip2(n9276), .s(n9947), .op(
        n3197) );
  mux2_1 U10161 ( .ip1(\ANSWER/mem[3][8][6] ), .ip2(n9276), .s(n9948), .op(
        n3196) );
  mux2_1 U10162 ( .ip1(\ANSWER/mem[3][9][6] ), .ip2(n9278), .s(n9949), .op(
        n3195) );
  mux2_1 U10163 ( .ip1(\ANSWER/mem[4][0][6] ), .ip2(n9276), .s(n9950), .op(
        n3194) );
  mux2_1 U10164 ( .ip1(\ANSWER/mem[4][1][6] ), .ip2(n9276), .s(n9951), .op(
        n3193) );
  mux2_1 U10165 ( .ip1(\ANSWER/mem[4][2][6] ), .ip2(n9278), .s(n9952), .op(
        n3192) );
  mux2_1 U10166 ( .ip1(\ANSWER/mem[4][3][6] ), .ip2(n9276), .s(n9953), .op(
        n3191) );
  mux2_1 U10167 ( .ip1(\ANSWER/mem[4][4][6] ), .ip2(n9277), .s(n9954), .op(
        n3190) );
  mux2_1 U10168 ( .ip1(\ANSWER/mem[4][5][6] ), .ip2(n9276), .s(n9955), .op(
        n3189) );
  mux2_1 U10169 ( .ip1(\ANSWER/mem[4][6][6] ), .ip2(n9277), .s(n9956), .op(
        n3188) );
  mux2_1 U10170 ( .ip1(\ANSWER/mem[4][7][6] ), .ip2(n9276), .s(n9957), .op(
        n3187) );
  mux2_1 U10171 ( .ip1(\ANSWER/mem[4][8][6] ), .ip2(n9278), .s(n9958), .op(
        n3186) );
  mux2_1 U10172 ( .ip1(\ANSWER/mem[4][9][6] ), .ip2(n9278), .s(n9959), .op(
        n3185) );
  mux2_1 U10173 ( .ip1(\ANSWER/mem[5][0][6] ), .ip2(n9278), .s(n9960), .op(
        n3184) );
  mux2_1 U10174 ( .ip1(\ANSWER/mem[5][1][6] ), .ip2(n9278), .s(n9961), .op(
        n3183) );
  mux2_1 U10175 ( .ip1(\ANSWER/mem[5][2][6] ), .ip2(n9278), .s(n9962), .op(
        n3182) );
  mux2_1 U10176 ( .ip1(\ANSWER/mem[5][3][6] ), .ip2(n9278), .s(n9963), .op(
        n3181) );
  mux2_1 U10177 ( .ip1(\ANSWER/mem[5][4][6] ), .ip2(n9278), .s(n9964), .op(
        n3180) );
  mux2_1 U10178 ( .ip1(\ANSWER/mem[5][5][6] ), .ip2(n9278), .s(n9965), .op(
        n3179) );
  mux2_1 U10179 ( .ip1(\ANSWER/mem[5][6][6] ), .ip2(n9278), .s(n9966), .op(
        n3178) );
  mux2_1 U10180 ( .ip1(\ANSWER/mem[5][7][6] ), .ip2(n9278), .s(n9967), .op(
        n3177) );
  mux2_1 U10181 ( .ip1(\ANSWER/mem[5][8][6] ), .ip2(n9278), .s(n9968), .op(
        n3176) );
  mux2_1 U10182 ( .ip1(\ANSWER/mem[5][9][6] ), .ip2(n9278), .s(n9969), .op(
        n3175) );
  mux2_1 U10183 ( .ip1(\ANSWER/mem[6][0][6] ), .ip2(n9277), .s(n9970), .op(
        n3174) );
  mux2_1 U10184 ( .ip1(\ANSWER/mem[6][1][6] ), .ip2(n9277), .s(n9971), .op(
        n3173) );
  mux2_1 U10185 ( .ip1(\ANSWER/mem[6][2][6] ), .ip2(n9277), .s(n9972), .op(
        n3172) );
  mux2_1 U10186 ( .ip1(\ANSWER/mem[6][3][6] ), .ip2(n9276), .s(n9973), .op(
        n3171) );
  mux2_1 U10187 ( .ip1(\ANSWER/mem[6][4][6] ), .ip2(n9278), .s(n9974), .op(
        n3170) );
  mux2_1 U10188 ( .ip1(\ANSWER/mem[6][5][6] ), .ip2(n9276), .s(n9975), .op(
        n3169) );
  mux2_1 U10189 ( .ip1(\ANSWER/mem[6][6][6] ), .ip2(n9278), .s(n9976), .op(
        n3168) );
  mux2_1 U10190 ( .ip1(\ANSWER/mem[6][7][6] ), .ip2(n9276), .s(n9977), .op(
        n3167) );
  mux2_1 U10191 ( .ip1(\ANSWER/mem[6][8][6] ), .ip2(n9278), .s(n9978), .op(
        n3166) );
  mux2_1 U10192 ( .ip1(\ANSWER/mem[6][9][6] ), .ip2(n9276), .s(n9979), .op(
        n3165) );
  mux2_1 U10193 ( .ip1(\ANSWER/mem[7][0][6] ), .ip2(n9276), .s(n9980), .op(
        n3164) );
  mux2_1 U10194 ( .ip1(\ANSWER/mem[7][1][6] ), .ip2(n9278), .s(n9981), .op(
        n3163) );
  mux2_1 U10195 ( .ip1(\ANSWER/mem[7][2][6] ), .ip2(n9277), .s(n9983), .op(
        n3162) );
  mux2_1 U10196 ( .ip1(\ANSWER/mem[7][3][6] ), .ip2(n9276), .s(n9984), .op(
        n3161) );
  mux2_1 U10197 ( .ip1(\ANSWER/mem[7][4][6] ), .ip2(n9277), .s(n9985), .op(
        n3160) );
  mux2_1 U10198 ( .ip1(\ANSWER/mem[7][5][6] ), .ip2(n9276), .s(n9986), .op(
        n3159) );
  mux2_1 U10199 ( .ip1(\ANSWER/mem[7][6][6] ), .ip2(n9278), .s(n9987), .op(
        n3158) );
  mux2_1 U10200 ( .ip1(\ANSWER/mem[7][7][6] ), .ip2(n9277), .s(n9988), .op(
        n3157) );
  mux2_1 U10201 ( .ip1(\ANSWER/mem[7][8][6] ), .ip2(n9277), .s(n9989), .op(
        n3156) );
  mux2_1 U10202 ( .ip1(\ANSWER/mem[7][9][6] ), .ip2(n9277), .s(n9990), .op(
        n3155) );
  mux2_1 U10203 ( .ip1(\ANSWER/mem[8][0][6] ), .ip2(n9277), .s(n9991), .op(
        n3154) );
  mux2_1 U10204 ( .ip1(\ANSWER/mem[8][1][6] ), .ip2(n9277), .s(n9992), .op(
        n3153) );
  mux2_1 U10205 ( .ip1(\ANSWER/mem[8][2][6] ), .ip2(n9277), .s(n9993), .op(
        n3152) );
  mux2_1 U10206 ( .ip1(\ANSWER/mem[8][3][6] ), .ip2(n9278), .s(n9994), .op(
        n3151) );
  mux2_1 U10207 ( .ip1(\ANSWER/mem[8][4][6] ), .ip2(n9276), .s(n9996), .op(
        n3150) );
  mux2_1 U10208 ( .ip1(\ANSWER/mem[8][5][6] ), .ip2(n9276), .s(n9997), .op(
        n3149) );
  mux2_1 U10209 ( .ip1(\ANSWER/mem[8][6][6] ), .ip2(n9278), .s(n9998), .op(
        n3148) );
  mux2_1 U10210 ( .ip1(\ANSWER/mem[8][7][6] ), .ip2(n9276), .s(n9999), .op(
        n3147) );
  mux2_1 U10211 ( .ip1(\ANSWER/mem[8][8][6] ), .ip2(n9277), .s(n10000), .op(
        n3146) );
  mux2_1 U10212 ( .ip1(\ANSWER/mem[8][9][6] ), .ip2(n9277), .s(n10001), .op(
        n3145) );
  mux2_1 U10213 ( .ip1(\ANSWER/mem[9][0][6] ), .ip2(n9277), .s(n10002), .op(
        n3144) );
  mux2_1 U10214 ( .ip1(\ANSWER/mem[9][1][6] ), .ip2(n9277), .s(n10003), .op(
        n3143) );
  mux2_1 U10215 ( .ip1(\ANSWER/mem[9][2][6] ), .ip2(n9277), .s(n10004), .op(
        n3142) );
  mux2_1 U10216 ( .ip1(\ANSWER/mem[9][3][6] ), .ip2(n9278), .s(n10005), .op(
        n3141) );
  mux2_1 U10217 ( .ip1(\ANSWER/mem[9][4][6] ), .ip2(n9277), .s(n10006), .op(
        n3140) );
  mux2_1 U10218 ( .ip1(\ANSWER/mem[9][5][6] ), .ip2(n9277), .s(n10007), .op(
        n3139) );
  mux2_1 U10219 ( .ip1(\ANSWER/mem[9][6][6] ), .ip2(n9277), .s(n10008), .op(
        n3138) );
  mux2_1 U10220 ( .ip1(\ANSWER/mem[9][7][6] ), .ip2(n9277), .s(n10009), .op(
        n3137) );
  mux2_1 U10221 ( .ip1(\ANSWER/mem[9][8][6] ), .ip2(n9278), .s(n10010), .op(
        n3136) );
  mux2_1 U10222 ( .ip1(\ANSWER/mem[9][9][6] ), .ip2(n9278), .s(n10011), .op(
        n3135) );
  nor2_1 U10223 ( .ip1(n9280), .ip2(n9279), .op(n9281) );
  nor2_1 U10224 ( .ip1(n9282), .ip2(n9281), .op(n9412) );
  inv_1 U10225 ( .ip(rdata[7]), .op(n9288) );
  nand2_1 U10226 ( .ip1(m2DataIn[2]), .ip2(q_w2[13]), .op(n9284) );
  inv_1 U10227 ( .ip(q_w2[14]), .op(n9816) );
  nor3_1 U10228 ( .ip1(n9500), .ip2(n9816), .ip3(n9283), .op(n9403) );
  or2_1 U10229 ( .ip1(n9284), .ip2(n9403), .op(n9287) );
  nand2_1 U10230 ( .ip1(m2DataIn[1]), .ip2(q_w2[14]), .op(n9285) );
  or2_1 U10231 ( .ip1(n9285), .ip2(n9403), .op(n9286) );
  nand2_1 U10232 ( .ip1(n9287), .ip2(n9286), .op(n9404) );
  mux2_1 U10233 ( .ip1(n9288), .ip2(rdata[7]), .s(n9404), .op(n9411) );
  or2_1 U10234 ( .ip1(n9289), .ip2(n9290), .op(n9293) );
  or2_1 U10235 ( .ip1(n9291), .ip2(n9290), .op(n9292) );
  nand2_1 U10236 ( .ip1(n9293), .ip2(n9292), .op(n9410) );
  inv_1 U10237 ( .ip(n9294), .op(n9428) );
  nor3_1 U10238 ( .ip1(n9817), .ip2(n9788), .ip3(n9295), .op(n9402) );
  nor2_1 U10239 ( .ip1(n9725), .ip2(n9788), .op(n9296) );
  or2_1 U10240 ( .ip1(q_w2[7]), .ip2(n9296), .op(n9298) );
  or2_1 U10241 ( .ip1(m2DataIn[8]), .ip2(n9296), .op(n9297) );
  nand2_1 U10242 ( .ip1(n9298), .ip2(n9297), .op(n9400) );
  nor2_1 U10243 ( .ip1(n9402), .ip2(n9400), .op(n9299) );
  nand2_1 U10244 ( .ip1(m2DataIn[13]), .ip2(q_w2[2]), .op(n9399) );
  xor2_1 U10245 ( .ip1(n9299), .ip2(n9399), .op(n9409) );
  nor2_1 U10246 ( .ip1(n9301), .ip2(n9300), .op(n9302) );
  nor2_1 U10247 ( .ip1(n9303), .ip2(n9302), .op(n9408) );
  or2_1 U10248 ( .ip1(n9304), .ip2(n9305), .op(n9308) );
  or2_1 U10249 ( .ip1(n9306), .ip2(n9305), .op(n9307) );
  nand2_1 U10250 ( .ip1(n9308), .ip2(n9307), .op(n9407) );
  inv_1 U10251 ( .ip(n9309), .op(n9427) );
  fulladder U10252 ( .a(n9312), .b(n9311), .ci(n9310), .co(n9426), .s(n9326)
         );
  nand2_1 U10253 ( .ip1(rdata[6]), .ip2(n9313), .op(n9314) );
  nand2_1 U10254 ( .ip1(n9315), .ip2(n9314), .op(n9421) );
  nand2_1 U10255 ( .ip1(q_w2[4]), .ip2(m2DataIn[11]), .op(n9317) );
  nor2_1 U10256 ( .ip1(n9372), .ip2(n9815), .op(n9316) );
  xor2_1 U10257 ( .ip1(n9317), .ip2(n9316), .op(n9420) );
  xor2_1 U10258 ( .ip1(n9421), .ip2(n9420), .op(n9432) );
  fulladder U10259 ( .a(n9320), .b(n9319), .ci(n9318), .co(n9431), .s(n9328)
         );
  fulladder U10260 ( .a(n9322), .b(n9419), .ci(n9321), .co(n9430), .s(n9329)
         );
  inv_1 U10261 ( .ip(n9323), .op(n9435) );
  fulladder U10262 ( .a(n9326), .b(n9325), .ci(n9324), .co(n9434), .s(n9264)
         );
  fulladder U10263 ( .a(n9329), .b(n9328), .ci(n9327), .co(n9415), .s(n9230)
         );
  nor3_1 U10264 ( .ip1(n9467), .ip2(n9791), .ip3(n9330), .op(n9382) );
  nor2_1 U10265 ( .ip1(n9467), .ip2(n9864), .op(n9373) );
  or2_1 U10266 ( .ip1(q_w2[11]), .ip2(n9373), .op(n9332) );
  or2_1 U10267 ( .ip1(m2DataIn[4]), .ip2(n9373), .op(n9331) );
  nand2_1 U10268 ( .ip1(n9332), .ip2(n9331), .op(n9333) );
  nor2_1 U10269 ( .ip1(n9382), .ip2(n9333), .op(n9381) );
  nor2_1 U10270 ( .ip1(n9863), .ip2(n9334), .op(n9383) );
  xor2_1 U10271 ( .ip1(n9381), .ip2(n9383), .op(n9397) );
  nor2_1 U10272 ( .ip1(n9792), .ip2(n9703), .op(n9380) );
  nand2_1 U10273 ( .ip1(m2DataIn[15]), .ip2(q_w2[0]), .op(n9378) );
  inv_1 U10274 ( .ip(q_w2[15]), .op(n9701) );
  nor2_1 U10275 ( .ip1(n9335), .ip2(n9701), .op(n9393) );
  nand2_1 U10276 ( .ip1(m2DataIn[9]), .ip2(q_w2[6]), .op(n9391) );
  inv_1 U10277 ( .ip(n9336), .op(n9395) );
  inv_1 U10278 ( .ip(n9337), .op(n9414) );
  fulladder U10279 ( .a(n9340), .b(n9339), .ci(n9338), .co(n9413), .s(n9260)
         );
  inv_1 U10280 ( .ip(n9341), .op(n9442) );
  fulladder U10281 ( .a(n9344), .b(n9343), .ci(n9342), .co(n9441), .s(n9234)
         );
  inv_1 U10282 ( .ip(n9345), .op(n9367) );
  inv_1 U10283 ( .ip(n9346), .op(n9348) );
  or2_1 U10284 ( .ip1(n9348), .ip2(n9347), .op(n9349) );
  nand2_1 U10285 ( .ip1(n9350), .ip2(n9349), .op(n9366) );
  fulladder U10286 ( .a(n9353), .b(n9352), .ci(n9351), .co(n9365), .s(n9268)
         );
  nor3_1 U10287 ( .ip1(\SIGMOID/lut_out [6]), .ip2(\SIGMOID/lut_out [5]), 
        .ip3(n9354), .op(n9363) );
  nor2_1 U10288 ( .ip1(\SIGMOID/sign_bit ), .ip2(n9363), .op(n9355) );
  xor2_1 U10289 ( .ip1(\SIGMOID/lut_out [7]), .ip2(n9355), .op(n10433) );
  nor2_1 U10290 ( .ip1(n10433), .ip2(n9445), .op(n9357) );
  or2_1 U10291 ( .ip1(n9356), .ip2(n9357), .op(n9359) );
  or2_1 U10292 ( .ip1(n9445), .ip2(n9357), .op(n9358) );
  nand2_1 U10293 ( .ip1(n9359), .ip2(n9358), .op(n9361) );
  buf_1 U10294 ( .ip(n9361), .op(n9360) );
  mux2_1 U10295 ( .ip1(\ANSWER/mem[0][0][7] ), .ip2(n9360), .s(n9910), .op(
        n3134) );
  mux2_1 U10296 ( .ip1(\ANSWER/mem[0][1][7] ), .ip2(n9360), .s(n9911), .op(
        n3133) );
  mux2_1 U10297 ( .ip1(\ANSWER/mem[0][2][7] ), .ip2(n9360), .s(n9912), .op(
        n3132) );
  mux2_1 U10298 ( .ip1(\ANSWER/mem[0][3][7] ), .ip2(n9360), .s(n9913), .op(
        n3131) );
  mux2_1 U10299 ( .ip1(\ANSWER/mem[0][4][7] ), .ip2(n9360), .s(n9914), .op(
        n3130) );
  mux2_1 U10300 ( .ip1(\ANSWER/mem[0][5][7] ), .ip2(n9360), .s(n9915), .op(
        n3129) );
  mux2_1 U10301 ( .ip1(\ANSWER/mem[0][6][7] ), .ip2(n9360), .s(n9916), .op(
        n3128) );
  mux2_1 U10302 ( .ip1(\ANSWER/mem[0][7][7] ), .ip2(n9360), .s(n9917), .op(
        n3127) );
  mux2_1 U10303 ( .ip1(\ANSWER/mem[0][8][7] ), .ip2(n9360), .s(n9918), .op(
        n3126) );
  mux2_1 U10304 ( .ip1(\ANSWER/mem[0][9][7] ), .ip2(n9360), .s(n9919), .op(
        n3125) );
  mux2_1 U10305 ( .ip1(\ANSWER/mem[1][0][7] ), .ip2(n9360), .s(n9920), .op(
        n3124) );
  mux2_1 U10306 ( .ip1(\ANSWER/mem[1][1][7] ), .ip2(n9360), .s(n9921), .op(
        n3123) );
  mux2_1 U10307 ( .ip1(\ANSWER/mem[1][2][7] ), .ip2(n9360), .s(n9922), .op(
        n3122) );
  mux2_1 U10308 ( .ip1(\ANSWER/mem[1][3][7] ), .ip2(n9360), .s(n9923), .op(
        n3121) );
  mux2_1 U10309 ( .ip1(\ANSWER/mem[1][4][7] ), .ip2(n9360), .s(n9924), .op(
        n3120) );
  mux2_1 U10310 ( .ip1(\ANSWER/mem[1][5][7] ), .ip2(n9360), .s(n9925), .op(
        n3119) );
  mux2_1 U10311 ( .ip1(\ANSWER/mem[1][6][7] ), .ip2(n9360), .s(n9926), .op(
        n3118) );
  mux2_1 U10312 ( .ip1(\ANSWER/mem[1][7][7] ), .ip2(n9360), .s(n9927), .op(
        n3117) );
  mux2_1 U10313 ( .ip1(\ANSWER/mem[1][8][7] ), .ip2(n9360), .s(n9928), .op(
        n3116) );
  mux2_1 U10314 ( .ip1(\ANSWER/mem[1][9][7] ), .ip2(n9360), .s(n9929), .op(
        n3115) );
  mux2_1 U10315 ( .ip1(\ANSWER/mem[2][0][7] ), .ip2(n9360), .s(n9930), .op(
        n3114) );
  mux2_1 U10316 ( .ip1(\ANSWER/mem[2][1][7] ), .ip2(n9360), .s(n9931), .op(
        n3113) );
  mux2_1 U10317 ( .ip1(\ANSWER/mem[2][2][7] ), .ip2(n9360), .s(n9932), .op(
        n3112) );
  mux2_1 U10318 ( .ip1(\ANSWER/mem[2][3][7] ), .ip2(n9360), .s(n9933), .op(
        n3111) );
  mux2_1 U10319 ( .ip1(\ANSWER/mem[2][4][7] ), .ip2(n9360), .s(n9934), .op(
        n3110) );
  mux2_1 U10320 ( .ip1(\ANSWER/mem[2][5][7] ), .ip2(n9360), .s(n9935), .op(
        n3109) );
  mux2_1 U10321 ( .ip1(\ANSWER/mem[2][6][7] ), .ip2(n9360), .s(n9936), .op(
        n3108) );
  mux2_1 U10322 ( .ip1(\ANSWER/mem[2][7][7] ), .ip2(n9360), .s(n9937), .op(
        n3107) );
  mux2_1 U10323 ( .ip1(\ANSWER/mem[2][8][7] ), .ip2(n9360), .s(n9938), .op(
        n3106) );
  mux2_1 U10324 ( .ip1(\ANSWER/mem[2][9][7] ), .ip2(n9360), .s(n9939), .op(
        n3105) );
  mux2_1 U10325 ( .ip1(\ANSWER/mem[3][0][7] ), .ip2(n9360), .s(n9940), .op(
        n3104) );
  mux2_1 U10326 ( .ip1(\ANSWER/mem[3][1][7] ), .ip2(n9360), .s(n9941), .op(
        n3103) );
  mux2_1 U10327 ( .ip1(\ANSWER/mem[3][2][7] ), .ip2(n9360), .s(n9942), .op(
        n3102) );
  mux2_1 U10328 ( .ip1(\ANSWER/mem[3][3][7] ), .ip2(n9360), .s(n9943), .op(
        n3101) );
  mux2_1 U10329 ( .ip1(\ANSWER/mem[3][4][7] ), .ip2(n9360), .s(n9944), .op(
        n3100) );
  mux2_1 U10330 ( .ip1(\ANSWER/mem[3][5][7] ), .ip2(n9360), .s(n9945), .op(
        n3099) );
  mux2_1 U10331 ( .ip1(\ANSWER/mem[3][6][7] ), .ip2(n9361), .s(n9946), .op(
        n3098) );
  mux2_1 U10332 ( .ip1(\ANSWER/mem[3][7][7] ), .ip2(n9361), .s(n9947), .op(
        n3097) );
  mux2_1 U10333 ( .ip1(\ANSWER/mem[3][8][7] ), .ip2(n9361), .s(n9948), .op(
        n3096) );
  mux2_1 U10334 ( .ip1(\ANSWER/mem[3][9][7] ), .ip2(n9361), .s(n9949), .op(
        n3095) );
  mux2_1 U10335 ( .ip1(\ANSWER/mem[4][0][7] ), .ip2(n9361), .s(n9950), .op(
        n3094) );
  mux2_1 U10336 ( .ip1(\ANSWER/mem[4][1][7] ), .ip2(n9362), .s(n9951), .op(
        n3093) );
  mux2_1 U10337 ( .ip1(\ANSWER/mem[4][2][7] ), .ip2(n9362), .s(n9952), .op(
        n3092) );
  mux2_1 U10338 ( .ip1(\ANSWER/mem[4][3][7] ), .ip2(n9362), .s(n9953), .op(
        n3091) );
  mux2_1 U10339 ( .ip1(\ANSWER/mem[4][4][7] ), .ip2(n9362), .s(n9954), .op(
        n3090) );
  mux2_1 U10340 ( .ip1(\ANSWER/mem[4][5][7] ), .ip2(n9362), .s(n9955), .op(
        n3089) );
  mux2_1 U10341 ( .ip1(\ANSWER/mem[4][6][7] ), .ip2(n9362), .s(n9956), .op(
        n3088) );
  mux2_1 U10342 ( .ip1(\ANSWER/mem[4][7][7] ), .ip2(n9362), .s(n9957), .op(
        n3087) );
  mux2_1 U10343 ( .ip1(\ANSWER/mem[4][8][7] ), .ip2(n9362), .s(n9958), .op(
        n3086) );
  mux2_1 U10344 ( .ip1(\ANSWER/mem[4][9][7] ), .ip2(n9362), .s(n9959), .op(
        n3085) );
  mux2_1 U10345 ( .ip1(\ANSWER/mem[5][0][7] ), .ip2(n9362), .s(n9960), .op(
        n3084) );
  mux2_1 U10346 ( .ip1(\ANSWER/mem[5][1][7] ), .ip2(n9361), .s(n9961), .op(
        n3083) );
  mux2_1 U10347 ( .ip1(\ANSWER/mem[5][2][7] ), .ip2(n9362), .s(n9962), .op(
        n3082) );
  mux2_1 U10348 ( .ip1(\ANSWER/mem[5][3][7] ), .ip2(n9361), .s(n9963), .op(
        n3081) );
  mux2_1 U10349 ( .ip1(\ANSWER/mem[5][4][7] ), .ip2(n9362), .s(n9964), .op(
        n3080) );
  mux2_1 U10350 ( .ip1(\ANSWER/mem[5][5][7] ), .ip2(n9361), .s(n9965), .op(
        n3079) );
  mux2_1 U10351 ( .ip1(\ANSWER/mem[5][6][7] ), .ip2(n9361), .s(n9966), .op(
        n3078) );
  mux2_1 U10352 ( .ip1(\ANSWER/mem[5][7][7] ), .ip2(n9361), .s(n9967), .op(
        n3077) );
  mux2_1 U10353 ( .ip1(\ANSWER/mem[5][8][7] ), .ip2(n9361), .s(n9968), .op(
        n3076) );
  mux2_1 U10354 ( .ip1(\ANSWER/mem[5][9][7] ), .ip2(n9361), .s(n9969), .op(
        n3075) );
  mux2_1 U10355 ( .ip1(\ANSWER/mem[6][0][7] ), .ip2(n9361), .s(n9970), .op(
        n3074) );
  mux2_1 U10356 ( .ip1(\ANSWER/mem[6][1][7] ), .ip2(n9361), .s(n9971), .op(
        n3073) );
  mux2_1 U10357 ( .ip1(\ANSWER/mem[6][2][7] ), .ip2(n9361), .s(n9972), .op(
        n3072) );
  mux2_1 U10358 ( .ip1(\ANSWER/mem[6][3][7] ), .ip2(n9361), .s(n9973), .op(
        n3071) );
  mux2_1 U10359 ( .ip1(\ANSWER/mem[6][4][7] ), .ip2(n9361), .s(n9974), .op(
        n3070) );
  mux2_1 U10360 ( .ip1(\ANSWER/mem[6][5][7] ), .ip2(n9361), .s(n9975), .op(
        n3069) );
  mux2_1 U10361 ( .ip1(\ANSWER/mem[6][6][7] ), .ip2(n9361), .s(n9976), .op(
        n3068) );
  mux2_1 U10362 ( .ip1(\ANSWER/mem[6][7][7] ), .ip2(n9361), .s(n9977), .op(
        n3067) );
  mux2_1 U10363 ( .ip1(\ANSWER/mem[6][8][7] ), .ip2(n9361), .s(n9978), .op(
        n3066) );
  mux2_1 U10364 ( .ip1(\ANSWER/mem[6][9][7] ), .ip2(n9361), .s(n9979), .op(
        n3065) );
  mux2_1 U10365 ( .ip1(\ANSWER/mem[7][0][7] ), .ip2(n9361), .s(n9980), .op(
        n3064) );
  mux2_1 U10366 ( .ip1(\ANSWER/mem[7][1][7] ), .ip2(n9361), .s(n9981), .op(
        n3063) );
  buf_1 U10367 ( .ip(n9361), .op(n9362) );
  mux2_1 U10368 ( .ip1(\ANSWER/mem[7][2][7] ), .ip2(n9362), .s(n9983), .op(
        n3062) );
  mux2_1 U10369 ( .ip1(\ANSWER/mem[7][3][7] ), .ip2(n9362), .s(n9984), .op(
        n3061) );
  mux2_1 U10370 ( .ip1(\ANSWER/mem[7][4][7] ), .ip2(n9362), .s(n9985), .op(
        n3060) );
  mux2_1 U10371 ( .ip1(\ANSWER/mem[7][5][7] ), .ip2(n9362), .s(n9986), .op(
        n3059) );
  mux2_1 U10372 ( .ip1(\ANSWER/mem[7][6][7] ), .ip2(n9362), .s(n9987), .op(
        n3058) );
  mux2_1 U10373 ( .ip1(\ANSWER/mem[7][7][7] ), .ip2(n9362), .s(n9988), .op(
        n3057) );
  mux2_1 U10374 ( .ip1(\ANSWER/mem[7][8][7] ), .ip2(n9362), .s(n9989), .op(
        n3056) );
  mux2_1 U10375 ( .ip1(\ANSWER/mem[7][9][7] ), .ip2(n9361), .s(n9990), .op(
        n3055) );
  mux2_1 U10376 ( .ip1(\ANSWER/mem[8][0][7] ), .ip2(n9361), .s(n9991), .op(
        n3054) );
  mux2_1 U10377 ( .ip1(\ANSWER/mem[8][1][7] ), .ip2(n9362), .s(n9992), .op(
        n3053) );
  mux2_1 U10378 ( .ip1(\ANSWER/mem[8][2][7] ), .ip2(n9362), .s(n9993), .op(
        n3052) );
  mux2_1 U10379 ( .ip1(\ANSWER/mem[8][3][7] ), .ip2(n9362), .s(n9994), .op(
        n3051) );
  mux2_1 U10380 ( .ip1(\ANSWER/mem[8][4][7] ), .ip2(n9361), .s(n9996), .op(
        n3050) );
  mux2_1 U10381 ( .ip1(\ANSWER/mem[8][5][7] ), .ip2(n9361), .s(n9997), .op(
        n3049) );
  mux2_1 U10382 ( .ip1(\ANSWER/mem[8][6][7] ), .ip2(n9361), .s(n9998), .op(
        n3048) );
  mux2_1 U10383 ( .ip1(\ANSWER/mem[8][7][7] ), .ip2(n9361), .s(n9999), .op(
        n3047) );
  mux2_1 U10384 ( .ip1(\ANSWER/mem[8][8][7] ), .ip2(n9361), .s(n10000), .op(
        n3046) );
  mux2_1 U10385 ( .ip1(\ANSWER/mem[8][9][7] ), .ip2(n9361), .s(n10001), .op(
        n3045) );
  mux2_1 U10386 ( .ip1(\ANSWER/mem[9][0][7] ), .ip2(n9361), .s(n10002), .op(
        n3044) );
  mux2_1 U10387 ( .ip1(\ANSWER/mem[9][1][7] ), .ip2(n9361), .s(n10003), .op(
        n3043) );
  mux2_1 U10388 ( .ip1(\ANSWER/mem[9][2][7] ), .ip2(n9361), .s(n10004), .op(
        n3042) );
  mux2_1 U10389 ( .ip1(\ANSWER/mem[9][3][7] ), .ip2(n9361), .s(n10005), .op(
        n3041) );
  mux2_1 U10390 ( .ip1(\ANSWER/mem[9][4][7] ), .ip2(n9361), .s(n10006), .op(
        n3040) );
  mux2_1 U10391 ( .ip1(\ANSWER/mem[9][5][7] ), .ip2(n9361), .s(n10007), .op(
        n3039) );
  mux2_1 U10392 ( .ip1(\ANSWER/mem[9][6][7] ), .ip2(n9362), .s(n10008), .op(
        n3038) );
  mux2_1 U10393 ( .ip1(\ANSWER/mem[9][7][7] ), .ip2(n9362), .s(n10009), .op(
        n3037) );
  mux2_1 U10394 ( .ip1(\ANSWER/mem[9][8][7] ), .ip2(n9362), .s(n10010), .op(
        n3036) );
  mux2_1 U10395 ( .ip1(\ANSWER/mem[9][9][7] ), .ip2(n9362), .s(n10011), .op(
        n3035) );
  inv_1 U10396 ( .ip(n9363), .op(n9364) );
  nor3_1 U10397 ( .ip1(\SIGMOID/sign_bit ), .ip2(\SIGMOID/lut_out [7]), .ip3(
        n9364), .op(n10019) );
  fulladder U10398 ( .a(n9367), .b(n9366), .ci(n9365), .co(n9439), .s(n9356)
         );
  and3_1 U10399 ( .ip1(m2DataIn[11]), .ip2(q_w2[6]), .ip3(n9380), .op(n9480)
         );
  nor2_1 U10400 ( .ip1(n9792), .ip2(n9732), .op(n9368) );
  or2_1 U10401 ( .ip1(q_w2[5]), .ip2(n9368), .op(n9370) );
  or2_1 U10402 ( .ip1(m2DataIn[11]), .ip2(n9368), .op(n9369) );
  nand2_1 U10403 ( .ip1(n9370), .ip2(n9369), .op(n9371) );
  nor2_1 U10404 ( .ip1(n9480), .ip2(n9371), .op(n9479) );
  nor2_1 U10405 ( .ip1(n9799), .ip2(n9372), .op(n9481) );
  xor2_1 U10406 ( .ip1(n9479), .ip2(n9481), .op(n9491) );
  and3_1 U10407 ( .ip1(m2DataIn[7]), .ip2(q_w2[10]), .ip3(n9373), .op(n9454)
         );
  nor2_1 U10408 ( .ip1(n9467), .ip2(n9814), .op(n9374) );
  or2_1 U10409 ( .ip1(q_w2[9]), .ip2(n9374), .op(n9376) );
  or2_1 U10410 ( .ip1(m2DataIn[7]), .ip2(n9374), .op(n9375) );
  nand2_1 U10411 ( .ip1(n9376), .ip2(n9375), .op(n9377) );
  nor2_1 U10412 ( .ip1(n9454), .ip2(n9377), .op(n9453) );
  nor2_1 U10413 ( .ip1(n9702), .ip2(n9791), .op(n9455) );
  xor2_1 U10414 ( .ip1(n9453), .ip2(n9455), .op(n9490) );
  fulladder U10415 ( .a(n9380), .b(n9379), .ci(n9378), .co(n9489), .s(n9396)
         );
  or2_1 U10416 ( .ip1(n9381), .ip2(n9382), .op(n9385) );
  or2_1 U10417 ( .ip1(n9383), .ip2(n9382), .op(n9384) );
  nand2_1 U10418 ( .ip1(n9385), .ip2(n9384), .op(n9495) );
  nand2_1 U10419 ( .ip1(m2DataIn[2]), .ip2(q_w2[14]), .op(n9387) );
  nand2_1 U10420 ( .ip1(m2DataIn[9]), .ip2(q_w2[14]), .op(n9862) );
  nor2_1 U10421 ( .ip1(n9862), .ip2(n9386), .op(n9485) );
  or2_1 U10422 ( .ip1(n9387), .ip2(n9485), .op(n9390) );
  nand2_1 U10423 ( .ip1(m2DataIn[9]), .ip2(q_w2[7]), .op(n9388) );
  or2_1 U10424 ( .ip1(n9388), .ip2(n9485), .op(n9389) );
  nand2_1 U10425 ( .ip1(n9390), .ip2(n9389), .op(n9484) );
  mux2_1 U10426 ( .ip1(rdata[8]), .ip2(n9486), .s(n9484), .op(n9494) );
  fulladder U10427 ( .a(n9393), .b(n9392), .ci(n9391), .co(n9493), .s(n9336)
         );
  inv_1 U10428 ( .ip(n9394), .op(n9505) );
  fulladder U10429 ( .a(n9397), .b(n9396), .ci(n9395), .co(n9504), .s(n9337)
         );
  inv_1 U10430 ( .ip(n9398), .op(n9513) );
  nor2_1 U10431 ( .ip1(n9400), .ip2(n9399), .op(n9401) );
  nor2_1 U10432 ( .ip1(n9402), .ip2(n9401), .op(n9503) );
  nand2_1 U10433 ( .ip1(m2DataIn[12]), .ip2(q_w2[4]), .op(n9502) );
  or2_1 U10434 ( .ip1(rdata[7]), .ip2(n9403), .op(n9406) );
  or2_1 U10435 ( .ip1(n9404), .ip2(n9403), .op(n9405) );
  nand2_1 U10436 ( .ip1(n9406), .ip2(n9405), .op(n9501) );
  fulladder U10437 ( .a(n9409), .b(n9408), .ci(n9407), .co(n9509), .s(n9309)
         );
  fulladder U10438 ( .a(n9412), .b(n9411), .ci(n9410), .co(n9508), .s(n9294)
         );
  fulladder U10439 ( .a(n9415), .b(n9414), .ci(n9413), .co(n9511), .s(n9341)
         );
  inv_1 U10440 ( .ip(n9416), .op(n9452) );
  nor2_1 U10441 ( .ip1(n9417), .ip2(n9701), .op(n9461) );
  nand2_1 U10442 ( .ip1(m2DataIn[14]), .ip2(q_w2[2]), .op(n9459) );
  inv_1 U10443 ( .ip(n9418), .op(n9477) );
  nor2_1 U10444 ( .ip1(n9817), .ip2(n9788), .op(n9474) );
  inv_1 U10445 ( .ip(q_w2[12]), .op(n9724) );
  nor2_1 U10446 ( .ip1(n9640), .ip2(n9724), .op(n9473) );
  nand2_1 U10447 ( .ip1(m2DataIn[15]), .ip2(q_w2[1]), .op(n9472) );
  or2_1 U10448 ( .ip1(n9502), .ip2(n9419), .op(n9424) );
  inv_1 U10449 ( .ip(n9420), .op(n9422) );
  nand2_1 U10450 ( .ip1(n9422), .ip2(n9421), .op(n9423) );
  nand2_1 U10451 ( .ip1(n9424), .ip2(n9423), .op(n9475) );
  inv_1 U10452 ( .ip(n9425), .op(n9498) );
  fulladder U10453 ( .a(n9428), .b(n9427), .ci(n9426), .co(n9429), .s(n9436)
         );
  inv_1 U10454 ( .ip(n9429), .op(n9497) );
  fulladder U10455 ( .a(n9432), .b(n9431), .ci(n9430), .co(n9496), .s(n9323)
         );
  inv_1 U10456 ( .ip(n9433), .op(n9451) );
  fulladder U10457 ( .a(n9436), .b(n9435), .ci(n9434), .co(n9450), .s(n9443)
         );
  inv_1 U10458 ( .ip(n9437), .op(n9438) );
  nand2_1 U10459 ( .ip1(n9439), .ip2(n9438), .op(n9517) );
  inv_1 U10460 ( .ip(n9517), .op(n9440) );
  nor2_1 U10461 ( .ip1(n9439), .ip2(n9438), .op(n9515) );
  nor2_1 U10462 ( .ip1(n9440), .ip2(n9515), .op(n9444) );
  fulladder U10463 ( .a(n9443), .b(n9442), .ci(n9441), .co(n9514), .s(n9345)
         );
  xor2_1 U10464 ( .ip1(n9444), .ip2(n9514), .op(n9446) );
  mux2_1 U10465 ( .ip1(n10019), .ip2(n9446), .s(n9445), .op(n9448) );
  buf_1 U10466 ( .ip(n9448), .op(n9447) );
  mux2_1 U10467 ( .ip1(\ANSWER/mem[0][0][8] ), .ip2(n9447), .s(n9910), .op(
        n3034) );
  mux2_1 U10468 ( .ip1(\ANSWER/mem[0][1][8] ), .ip2(n9447), .s(n9911), .op(
        n3033) );
  mux2_1 U10469 ( .ip1(\ANSWER/mem[0][2][8] ), .ip2(n9447), .s(n9912), .op(
        n3032) );
  mux2_1 U10470 ( .ip1(\ANSWER/mem[0][3][8] ), .ip2(n9447), .s(n9913), .op(
        n3031) );
  mux2_1 U10471 ( .ip1(\ANSWER/mem[0][4][8] ), .ip2(n9447), .s(n9914), .op(
        n3030) );
  mux2_1 U10472 ( .ip1(\ANSWER/mem[0][5][8] ), .ip2(n9447), .s(n9915), .op(
        n3029) );
  mux2_1 U10473 ( .ip1(\ANSWER/mem[0][6][8] ), .ip2(n9447), .s(n9916), .op(
        n3028) );
  mux2_1 U10474 ( .ip1(\ANSWER/mem[0][7][8] ), .ip2(n9447), .s(n9917), .op(
        n3027) );
  mux2_1 U10475 ( .ip1(\ANSWER/mem[0][8][8] ), .ip2(n9447), .s(n9918), .op(
        n3026) );
  mux2_1 U10476 ( .ip1(\ANSWER/mem[0][9][8] ), .ip2(n9447), .s(n9919), .op(
        n3025) );
  mux2_1 U10477 ( .ip1(\ANSWER/mem[1][0][8] ), .ip2(n9447), .s(n9920), .op(
        n3024) );
  mux2_1 U10478 ( .ip1(\ANSWER/mem[1][1][8] ), .ip2(n9447), .s(n9921), .op(
        n3023) );
  mux2_1 U10479 ( .ip1(\ANSWER/mem[1][2][8] ), .ip2(n9447), .s(n9922), .op(
        n3022) );
  mux2_1 U10480 ( .ip1(\ANSWER/mem[1][3][8] ), .ip2(n9447), .s(n9923), .op(
        n3021) );
  mux2_1 U10481 ( .ip1(\ANSWER/mem[1][4][8] ), .ip2(n9447), .s(n9924), .op(
        n3020) );
  mux2_1 U10482 ( .ip1(\ANSWER/mem[1][5][8] ), .ip2(n9447), .s(n9925), .op(
        n3019) );
  mux2_1 U10483 ( .ip1(\ANSWER/mem[1][6][8] ), .ip2(n9447), .s(n9926), .op(
        n3018) );
  mux2_1 U10484 ( .ip1(\ANSWER/mem[1][7][8] ), .ip2(n9447), .s(n9927), .op(
        n3017) );
  mux2_1 U10485 ( .ip1(\ANSWER/mem[1][8][8] ), .ip2(n9447), .s(n9928), .op(
        n3016) );
  mux2_1 U10486 ( .ip1(\ANSWER/mem[1][9][8] ), .ip2(n9447), .s(n9929), .op(
        n3015) );
  mux2_1 U10487 ( .ip1(\ANSWER/mem[2][0][8] ), .ip2(n9447), .s(n9930), .op(
        n3014) );
  mux2_1 U10488 ( .ip1(\ANSWER/mem[2][1][8] ), .ip2(n9447), .s(n9931), .op(
        n3013) );
  mux2_1 U10489 ( .ip1(\ANSWER/mem[2][2][8] ), .ip2(n9447), .s(n9932), .op(
        n3012) );
  mux2_1 U10490 ( .ip1(\ANSWER/mem[2][3][8] ), .ip2(n9447), .s(n9933), .op(
        n3011) );
  mux2_1 U10491 ( .ip1(\ANSWER/mem[2][4][8] ), .ip2(n9447), .s(n9934), .op(
        n3010) );
  mux2_1 U10492 ( .ip1(\ANSWER/mem[2][5][8] ), .ip2(n9447), .s(n9935), .op(
        n3009) );
  mux2_1 U10493 ( .ip1(\ANSWER/mem[2][6][8] ), .ip2(n9447), .s(n9936), .op(
        n3008) );
  mux2_1 U10494 ( .ip1(\ANSWER/mem[2][7][8] ), .ip2(n9447), .s(n9937), .op(
        n3007) );
  mux2_1 U10495 ( .ip1(\ANSWER/mem[2][8][8] ), .ip2(n9447), .s(n9938), .op(
        n3006) );
  mux2_1 U10496 ( .ip1(\ANSWER/mem[2][9][8] ), .ip2(n9447), .s(n9939), .op(
        n3005) );
  mux2_1 U10497 ( .ip1(\ANSWER/mem[3][0][8] ), .ip2(n9447), .s(n9940), .op(
        n3004) );
  mux2_1 U10498 ( .ip1(\ANSWER/mem[3][1][8] ), .ip2(n9447), .s(n9941), .op(
        n3003) );
  mux2_1 U10499 ( .ip1(\ANSWER/mem[3][2][8] ), .ip2(n9447), .s(n9942), .op(
        n3002) );
  mux2_1 U10500 ( .ip1(\ANSWER/mem[3][3][8] ), .ip2(n9447), .s(n9943), .op(
        n3001) );
  mux2_1 U10501 ( .ip1(\ANSWER/mem[3][4][8] ), .ip2(n9447), .s(n9944), .op(
        n3000) );
  mux2_1 U10502 ( .ip1(\ANSWER/mem[3][5][8] ), .ip2(n9447), .s(n9945), .op(
        n2999) );
  mux2_1 U10503 ( .ip1(\ANSWER/mem[3][6][8] ), .ip2(n9448), .s(n9946), .op(
        n2998) );
  mux2_1 U10504 ( .ip1(\ANSWER/mem[3][7][8] ), .ip2(n9448), .s(n9947), .op(
        n2997) );
  mux2_1 U10505 ( .ip1(\ANSWER/mem[3][8][8] ), .ip2(n9448), .s(n9948), .op(
        n2996) );
  mux2_1 U10506 ( .ip1(\ANSWER/mem[3][9][8] ), .ip2(n9448), .s(n9949), .op(
        n2995) );
  mux2_1 U10507 ( .ip1(\ANSWER/mem[4][0][8] ), .ip2(n9448), .s(n9950), .op(
        n2994) );
  mux2_1 U10508 ( .ip1(\ANSWER/mem[4][1][8] ), .ip2(n9448), .s(n9951), .op(
        n2993) );
  mux2_1 U10509 ( .ip1(\ANSWER/mem[4][2][8] ), .ip2(n9449), .s(n9952), .op(
        n2992) );
  mux2_1 U10510 ( .ip1(\ANSWER/mem[4][3][8] ), .ip2(n9449), .s(n9953), .op(
        n2991) );
  mux2_1 U10511 ( .ip1(\ANSWER/mem[4][4][8] ), .ip2(n9449), .s(n9954), .op(
        n2990) );
  mux2_1 U10512 ( .ip1(\ANSWER/mem[4][5][8] ), .ip2(n9449), .s(n9955), .op(
        n2989) );
  mux2_1 U10513 ( .ip1(\ANSWER/mem[4][6][8] ), .ip2(n9449), .s(n9956), .op(
        n2988) );
  mux2_1 U10514 ( .ip1(\ANSWER/mem[4][7][8] ), .ip2(n9449), .s(n9957), .op(
        n2987) );
  mux2_1 U10515 ( .ip1(\ANSWER/mem[4][8][8] ), .ip2(n9449), .s(n9958), .op(
        n2986) );
  mux2_1 U10516 ( .ip1(\ANSWER/mem[4][9][8] ), .ip2(n9449), .s(n9959), .op(
        n2985) );
  mux2_1 U10517 ( .ip1(\ANSWER/mem[5][0][8] ), .ip2(n9449), .s(n9960), .op(
        n2984) );
  mux2_1 U10518 ( .ip1(\ANSWER/mem[5][1][8] ), .ip2(n9448), .s(n9961), .op(
        n2983) );
  mux2_1 U10519 ( .ip1(\ANSWER/mem[5][2][8] ), .ip2(n9449), .s(n9962), .op(
        n2982) );
  mux2_1 U10520 ( .ip1(\ANSWER/mem[5][3][8] ), .ip2(n9448), .s(n9963), .op(
        n2981) );
  mux2_1 U10521 ( .ip1(\ANSWER/mem[5][4][8] ), .ip2(n9449), .s(n9964), .op(
        n2980) );
  mux2_1 U10522 ( .ip1(\ANSWER/mem[5][5][8] ), .ip2(n9448), .s(n9965), .op(
        n2979) );
  mux2_1 U10523 ( .ip1(\ANSWER/mem[5][6][8] ), .ip2(n9448), .s(n9966), .op(
        n2978) );
  mux2_1 U10524 ( .ip1(\ANSWER/mem[5][7][8] ), .ip2(n9448), .s(n9967), .op(
        n2977) );
  mux2_1 U10525 ( .ip1(\ANSWER/mem[5][8][8] ), .ip2(n9448), .s(n9968), .op(
        n2976) );
  mux2_1 U10526 ( .ip1(\ANSWER/mem[5][9][8] ), .ip2(n9448), .s(n9969), .op(
        n2975) );
  mux2_1 U10527 ( .ip1(\ANSWER/mem[6][0][8] ), .ip2(n9448), .s(n9970), .op(
        n2974) );
  mux2_1 U10528 ( .ip1(\ANSWER/mem[6][1][8] ), .ip2(n9448), .s(n9971), .op(
        n2973) );
  mux2_1 U10529 ( .ip1(\ANSWER/mem[6][2][8] ), .ip2(n9448), .s(n9972), .op(
        n2972) );
  mux2_1 U10530 ( .ip1(\ANSWER/mem[6][3][8] ), .ip2(n9448), .s(n9973), .op(
        n2971) );
  mux2_1 U10531 ( .ip1(\ANSWER/mem[6][4][8] ), .ip2(n9448), .s(n9974), .op(
        n2970) );
  mux2_1 U10532 ( .ip1(\ANSWER/mem[6][5][8] ), .ip2(n9448), .s(n9975), .op(
        n2969) );
  mux2_1 U10533 ( .ip1(\ANSWER/mem[6][6][8] ), .ip2(n9448), .s(n9976), .op(
        n2968) );
  mux2_1 U10534 ( .ip1(\ANSWER/mem[6][7][8] ), .ip2(n9448), .s(n9977), .op(
        n2967) );
  mux2_1 U10535 ( .ip1(\ANSWER/mem[6][8][8] ), .ip2(n9448), .s(n9978), .op(
        n2966) );
  mux2_1 U10536 ( .ip1(\ANSWER/mem[6][9][8] ), .ip2(n9448), .s(n9979), .op(
        n2965) );
  mux2_1 U10537 ( .ip1(\ANSWER/mem[7][0][8] ), .ip2(n9448), .s(n9980), .op(
        n2964) );
  mux2_1 U10538 ( .ip1(\ANSWER/mem[7][1][8] ), .ip2(n9448), .s(n9981), .op(
        n2963) );
  buf_1 U10539 ( .ip(n9448), .op(n9449) );
  mux2_1 U10540 ( .ip1(\ANSWER/mem[7][2][8] ), .ip2(n9449), .s(n9983), .op(
        n2962) );
  mux2_1 U10541 ( .ip1(\ANSWER/mem[7][3][8] ), .ip2(n9449), .s(n9984), .op(
        n2961) );
  mux2_1 U10542 ( .ip1(\ANSWER/mem[7][4][8] ), .ip2(n9449), .s(n9985), .op(
        n2960) );
  mux2_1 U10543 ( .ip1(\ANSWER/mem[7][5][8] ), .ip2(n9449), .s(n9986), .op(
        n2959) );
  mux2_1 U10544 ( .ip1(\ANSWER/mem[7][6][8] ), .ip2(n9449), .s(n9987), .op(
        n2958) );
  mux2_1 U10545 ( .ip1(\ANSWER/mem[7][7][8] ), .ip2(n9449), .s(n9988), .op(
        n2957) );
  mux2_1 U10546 ( .ip1(\ANSWER/mem[7][8][8] ), .ip2(n9449), .s(n9989), .op(
        n2956) );
  mux2_1 U10547 ( .ip1(\ANSWER/mem[7][9][8] ), .ip2(n9448), .s(n9990), .op(
        n2955) );
  mux2_1 U10548 ( .ip1(\ANSWER/mem[8][0][8] ), .ip2(n9449), .s(n9991), .op(
        n2954) );
  mux2_1 U10549 ( .ip1(\ANSWER/mem[8][1][8] ), .ip2(n9449), .s(n9992), .op(
        n2953) );
  mux2_1 U10550 ( .ip1(\ANSWER/mem[8][2][8] ), .ip2(n9449), .s(n9993), .op(
        n2952) );
  mux2_1 U10551 ( .ip1(\ANSWER/mem[8][3][8] ), .ip2(n9449), .s(n9994), .op(
        n2951) );
  mux2_1 U10552 ( .ip1(\ANSWER/mem[8][4][8] ), .ip2(n9448), .s(n9996), .op(
        n2950) );
  mux2_1 U10553 ( .ip1(\ANSWER/mem[8][5][8] ), .ip2(n9448), .s(n9997), .op(
        n2949) );
  mux2_1 U10554 ( .ip1(\ANSWER/mem[8][6][8] ), .ip2(n9448), .s(n9998), .op(
        n2948) );
  mux2_1 U10555 ( .ip1(\ANSWER/mem[8][7][8] ), .ip2(n9448), .s(n9999), .op(
        n2947) );
  mux2_1 U10556 ( .ip1(\ANSWER/mem[8][8][8] ), .ip2(n9448), .s(n10000), .op(
        n2946) );
  mux2_1 U10557 ( .ip1(\ANSWER/mem[8][9][8] ), .ip2(n9448), .s(n10001), .op(
        n2945) );
  mux2_1 U10558 ( .ip1(\ANSWER/mem[9][0][8] ), .ip2(n9448), .s(n10002), .op(
        n2944) );
  mux2_1 U10559 ( .ip1(\ANSWER/mem[9][1][8] ), .ip2(n9448), .s(n10003), .op(
        n2943) );
  mux2_1 U10560 ( .ip1(\ANSWER/mem[9][2][8] ), .ip2(n9448), .s(n10004), .op(
        n2942) );
  mux2_1 U10561 ( .ip1(\ANSWER/mem[9][3][8] ), .ip2(n9448), .s(n10005), .op(
        n2941) );
  mux2_1 U10562 ( .ip1(\ANSWER/mem[9][4][8] ), .ip2(n9448), .s(n10006), .op(
        n2940) );
  mux2_1 U10563 ( .ip1(\ANSWER/mem[9][5][8] ), .ip2(n9448), .s(n10007), .op(
        n2939) );
  mux2_1 U10564 ( .ip1(\ANSWER/mem[9][6][8] ), .ip2(n9449), .s(n10008), .op(
        n2938) );
  mux2_1 U10565 ( .ip1(\ANSWER/mem[9][7][8] ), .ip2(n9449), .s(n10009), .op(
        n2937) );
  mux2_1 U10566 ( .ip1(\ANSWER/mem[9][8][8] ), .ip2(n9449), .s(n10010), .op(
        n2936) );
  mux2_1 U10567 ( .ip1(\ANSWER/mem[9][9][8] ), .ip2(n9449), .s(n10011), .op(
        n2935) );
  fulladder U10568 ( .a(n9452), .b(n9451), .ci(n9450), .co(n9582), .s(n9437)
         );
  or2_1 U10569 ( .ip1(n9453), .ip2(n9454), .op(n9457) );
  or2_1 U10570 ( .ip1(n9455), .ip2(n9454), .op(n9456) );
  nand2_1 U10571 ( .ip1(n9457), .ip2(n9456), .op(n9542) );
  nor2_1 U10572 ( .ip1(n9790), .ip2(n9788), .op(n9533) );
  inv_1 U10573 ( .ip(n9458), .op(n9541) );
  fulladder U10574 ( .a(n9461), .b(n9460), .ci(n9459), .co(n9540), .s(n9418)
         );
  inv_1 U10575 ( .ip(n9462), .op(n9548) );
  nand2_1 U10576 ( .ip1(m2DataIn[11]), .ip2(q_w2[7]), .op(n9694) );
  nor3_1 U10577 ( .ip1(n9792), .ip2(n9732), .ip3(n9694), .op(n9562) );
  nor2_1 U10578 ( .ip1(n9735), .ip2(n9732), .op(n9463) );
  or2_1 U10579 ( .ip1(q_w2[7]), .ip2(n9463), .op(n9465) );
  or2_1 U10580 ( .ip1(m2DataIn[10]), .ip2(n9463), .op(n9464) );
  nand2_1 U10581 ( .ip1(n9465), .ip2(n9464), .op(n9466) );
  nor2_1 U10582 ( .ip1(n9562), .ip2(n9466), .op(n9561) );
  nor2_1 U10583 ( .ip1(n9799), .ip2(n9638), .op(n9563) );
  xor2_1 U10584 ( .ip1(n9561), .ip2(n9563), .op(n9538) );
  nand2_1 U10585 ( .ip1(m2DataIn[6]), .ip2(q_w2[11]), .op(n9468) );
  nand2_1 U10586 ( .ip1(m2DataIn[7]), .ip2(q_w2[11]), .op(n9625) );
  nor3_1 U10587 ( .ip1(n9467), .ip2(n9814), .ip3(n9625), .op(n9551) );
  or2_1 U10588 ( .ip1(n9468), .ip2(n9551), .op(n9471) );
  nand2_1 U10589 ( .ip1(m2DataIn[7]), .ip2(q_w2[10]), .op(n9469) );
  or2_1 U10590 ( .ip1(n9469), .ip2(n9551), .op(n9470) );
  nand2_1 U10591 ( .ip1(n9471), .ip2(n9470), .op(n9550) );
  nor2_1 U10592 ( .ip1(n9702), .ip2(n9724), .op(n9552) );
  xor2_1 U10593 ( .ip1(n9550), .ip2(n9552), .op(n9537) );
  fulladder U10594 ( .a(n9474), .b(n9473), .ci(n9472), .co(n9536), .s(n9476)
         );
  fulladder U10595 ( .a(n9477), .b(n9476), .ci(n9475), .co(n9546), .s(n9425)
         );
  inv_1 U10596 ( .ip(n9478), .op(n9581) );
  nand2_1 U10597 ( .ip1(m2DataIn[12]), .ip2(q_w2[5]), .op(n9600) );
  or2_1 U10598 ( .ip1(n9479), .ip2(n9480), .op(n9483) );
  or2_1 U10599 ( .ip1(n9481), .ip2(n9480), .op(n9482) );
  nand2_1 U10600 ( .ip1(n9483), .ip2(n9482), .op(n9532) );
  or2_1 U10601 ( .ip1(n9484), .ip2(n9485), .op(n9488) );
  or2_1 U10602 ( .ip1(n9486), .ip2(n9485), .op(n9487) );
  nand2_1 U10603 ( .ip1(n9488), .ip2(n9487), .op(n9531) );
  fulladder U10604 ( .a(n9491), .b(n9490), .ci(n9489), .co(n9492), .s(n9506)
         );
  inv_1 U10605 ( .ip(n9492), .op(n9544) );
  fulladder U10606 ( .a(n9495), .b(n9494), .ci(n9493), .co(n9543), .s(n9394)
         );
  fulladder U10607 ( .a(n9498), .b(n9497), .ci(n9496), .co(n9579), .s(n9433)
         );
  inv_1 U10608 ( .ip(m2DataIn[15]), .op(n9704) );
  nor2_1 U10609 ( .ip1(n9704), .ip2(n9499), .op(n9560) );
  nand2_1 U10610 ( .ip1(m2DataIn[4]), .ip2(q_w2[13]), .op(n9559) );
  nand2_1 U10611 ( .ip1(m2DataIn[8]), .ip2(q_w2[9]), .op(n9558) );
  nor2_1 U10612 ( .ip1(n9500), .ip2(n9701), .op(n9572) );
  nand2_1 U10613 ( .ip1(m2DataIn[14]), .ip2(q_w2[3]), .op(n9570) );
  fulladder U10614 ( .a(n9503), .b(n9502), .ci(n9501), .co(n9573), .s(n9510)
         );
  fulladder U10615 ( .a(n9506), .b(n9505), .ci(n9504), .co(n9507), .s(n9398)
         );
  inv_1 U10616 ( .ip(n9507), .op(n9577) );
  fulladder U10617 ( .a(n9510), .b(n9509), .ci(n9508), .co(n9576), .s(n9512)
         );
  fulladder U10618 ( .a(n9513), .b(n9512), .ci(n9511), .co(n9526), .s(n9416)
         );
  or2_1 U10619 ( .ip1(n9515), .ip2(n9514), .op(n9516) );
  nand2_1 U10620 ( .ip1(n9517), .ip2(n9516), .op(n9518) );
  nand2_1 U10621 ( .ip1(n9519), .ip2(n9518), .op(n9585) );
  inv_1 U10622 ( .ip(n9585), .op(n9520) );
  nor2_1 U10623 ( .ip1(n9519), .ip2(n9518), .op(n9583) );
  nor2_1 U10624 ( .ip1(n9520), .ip2(n9583), .op(n9522) );
  nor2_1 U10625 ( .ip1(n9582), .ip2(n9522), .op(n9521) );
  not_ab_or_c_or_d U10626 ( .ip1(n9582), .ip2(n9522), .ip3(n9907), .ip4(n9521), 
        .op(n9524) );
  buf_1 U10627 ( .ip(n9524), .op(n9523) );
  mux2_1 U10628 ( .ip1(\ANSWER/mem[0][0][9] ), .ip2(n9523), .s(n9910), .op(
        n2934) );
  mux2_1 U10629 ( .ip1(\ANSWER/mem[0][1][9] ), .ip2(n9523), .s(n9911), .op(
        n2933) );
  mux2_1 U10630 ( .ip1(\ANSWER/mem[0][2][9] ), .ip2(n9523), .s(n9912), .op(
        n2932) );
  mux2_1 U10631 ( .ip1(\ANSWER/mem[0][3][9] ), .ip2(n9523), .s(n9913), .op(
        n2931) );
  mux2_1 U10632 ( .ip1(\ANSWER/mem[0][4][9] ), .ip2(n9523), .s(n9914), .op(
        n2930) );
  mux2_1 U10633 ( .ip1(\ANSWER/mem[0][5][9] ), .ip2(n9523), .s(n9915), .op(
        n2929) );
  mux2_1 U10634 ( .ip1(\ANSWER/mem[0][6][9] ), .ip2(n9523), .s(n9916), .op(
        n2928) );
  mux2_1 U10635 ( .ip1(\ANSWER/mem[0][7][9] ), .ip2(n9523), .s(n9917), .op(
        n2927) );
  mux2_1 U10636 ( .ip1(\ANSWER/mem[0][8][9] ), .ip2(n9523), .s(n9918), .op(
        n2926) );
  mux2_1 U10637 ( .ip1(\ANSWER/mem[0][9][9] ), .ip2(n9523), .s(n9919), .op(
        n2925) );
  mux2_1 U10638 ( .ip1(\ANSWER/mem[1][0][9] ), .ip2(n9523), .s(n9920), .op(
        n2924) );
  mux2_1 U10639 ( .ip1(\ANSWER/mem[1][1][9] ), .ip2(n9523), .s(n9921), .op(
        n2923) );
  buf_1 U10640 ( .ip(n9524), .op(n9525) );
  mux2_1 U10641 ( .ip1(\ANSWER/mem[1][2][9] ), .ip2(n9525), .s(n9922), .op(
        n2922) );
  mux2_1 U10642 ( .ip1(\ANSWER/mem[1][3][9] ), .ip2(n9525), .s(n9923), .op(
        n2921) );
  mux2_1 U10643 ( .ip1(\ANSWER/mem[1][4][9] ), .ip2(n9525), .s(n9924), .op(
        n2920) );
  mux2_1 U10644 ( .ip1(\ANSWER/mem[1][5][9] ), .ip2(n9525), .s(n9925), .op(
        n2919) );
  mux2_1 U10645 ( .ip1(\ANSWER/mem[1][6][9] ), .ip2(n9525), .s(n9926), .op(
        n2918) );
  mux2_1 U10646 ( .ip1(\ANSWER/mem[1][7][9] ), .ip2(n9525), .s(n9927), .op(
        n2917) );
  mux2_1 U10647 ( .ip1(\ANSWER/mem[1][8][9] ), .ip2(n9525), .s(n9928), .op(
        n2916) );
  mux2_1 U10648 ( .ip1(\ANSWER/mem[1][9][9] ), .ip2(n9525), .s(n9929), .op(
        n2915) );
  mux2_1 U10649 ( .ip1(\ANSWER/mem[2][0][9] ), .ip2(n9525), .s(n9930), .op(
        n2914) );
  mux2_1 U10650 ( .ip1(\ANSWER/mem[2][1][9] ), .ip2(n9525), .s(n9931), .op(
        n2913) );
  mux2_1 U10651 ( .ip1(\ANSWER/mem[2][2][9] ), .ip2(n9525), .s(n9932), .op(
        n2912) );
  mux2_1 U10652 ( .ip1(\ANSWER/mem[2][3][9] ), .ip2(n9525), .s(n9933), .op(
        n2911) );
  mux2_1 U10653 ( .ip1(\ANSWER/mem[2][4][9] ), .ip2(n9523), .s(n9934), .op(
        n2910) );
  mux2_1 U10654 ( .ip1(\ANSWER/mem[2][5][9] ), .ip2(n9523), .s(n9935), .op(
        n2909) );
  mux2_1 U10655 ( .ip1(\ANSWER/mem[2][6][9] ), .ip2(n9523), .s(n9936), .op(
        n2908) );
  mux2_1 U10656 ( .ip1(\ANSWER/mem[2][7][9] ), .ip2(n9523), .s(n9937), .op(
        n2907) );
  mux2_1 U10657 ( .ip1(\ANSWER/mem[2][8][9] ), .ip2(n9523), .s(n9938), .op(
        n2906) );
  mux2_1 U10658 ( .ip1(\ANSWER/mem[2][9][9] ), .ip2(n9523), .s(n9939), .op(
        n2905) );
  mux2_1 U10659 ( .ip1(\ANSWER/mem[3][0][9] ), .ip2(n9523), .s(n9940), .op(
        n2904) );
  mux2_1 U10660 ( .ip1(\ANSWER/mem[3][1][9] ), .ip2(n9523), .s(n9941), .op(
        n2903) );
  mux2_1 U10661 ( .ip1(\ANSWER/mem[3][2][9] ), .ip2(n9523), .s(n9942), .op(
        n2902) );
  mux2_1 U10662 ( .ip1(\ANSWER/mem[3][3][9] ), .ip2(n9523), .s(n9943), .op(
        n2901) );
  mux2_1 U10663 ( .ip1(\ANSWER/mem[3][4][9] ), .ip2(n9523), .s(n9944), .op(
        n2900) );
  mux2_1 U10664 ( .ip1(\ANSWER/mem[3][5][9] ), .ip2(n9523), .s(n9945), .op(
        n2899) );
  mux2_1 U10665 ( .ip1(\ANSWER/mem[3][6][9] ), .ip2(n9525), .s(n9946), .op(
        n2898) );
  mux2_1 U10666 ( .ip1(\ANSWER/mem[3][7][9] ), .ip2(n9525), .s(n9947), .op(
        n2897) );
  mux2_1 U10667 ( .ip1(\ANSWER/mem[3][8][9] ), .ip2(n9525), .s(n9948), .op(
        n2896) );
  mux2_1 U10668 ( .ip1(\ANSWER/mem[3][9][9] ), .ip2(n9525), .s(n9949), .op(
        n2895) );
  mux2_1 U10669 ( .ip1(\ANSWER/mem[4][0][9] ), .ip2(n9525), .s(n9950), .op(
        n2894) );
  mux2_1 U10670 ( .ip1(\ANSWER/mem[4][1][9] ), .ip2(n9525), .s(n9951), .op(
        n2893) );
  mux2_1 U10671 ( .ip1(\ANSWER/mem[4][2][9] ), .ip2(n9525), .s(n9952), .op(
        n2892) );
  mux2_1 U10672 ( .ip1(\ANSWER/mem[4][3][9] ), .ip2(n9525), .s(n9953), .op(
        n2891) );
  mux2_1 U10673 ( .ip1(\ANSWER/mem[4][4][9] ), .ip2(n9525), .s(n9954), .op(
        n2890) );
  mux2_1 U10674 ( .ip1(\ANSWER/mem[4][5][9] ), .ip2(n9525), .s(n9955), .op(
        n2889) );
  mux2_1 U10675 ( .ip1(\ANSWER/mem[4][6][9] ), .ip2(n9525), .s(n9956), .op(
        n2888) );
  mux2_1 U10676 ( .ip1(\ANSWER/mem[4][7][9] ), .ip2(n9524), .s(n9957), .op(
        n2887) );
  mux2_1 U10677 ( .ip1(\ANSWER/mem[4][8][9] ), .ip2(n9524), .s(n9958), .op(
        n2886) );
  mux2_1 U10678 ( .ip1(\ANSWER/mem[4][9][9] ), .ip2(n9524), .s(n9959), .op(
        n2885) );
  mux2_1 U10679 ( .ip1(\ANSWER/mem[5][0][9] ), .ip2(n9524), .s(n9960), .op(
        n2884) );
  mux2_1 U10680 ( .ip1(\ANSWER/mem[5][1][9] ), .ip2(n9524), .s(n9961), .op(
        n2883) );
  mux2_1 U10681 ( .ip1(\ANSWER/mem[5][2][9] ), .ip2(n9524), .s(n9962), .op(
        n2882) );
  mux2_1 U10682 ( .ip1(\ANSWER/mem[5][3][9] ), .ip2(n9524), .s(n9963), .op(
        n2881) );
  mux2_1 U10683 ( .ip1(\ANSWER/mem[5][4][9] ), .ip2(n9524), .s(n9964), .op(
        n2880) );
  mux2_1 U10684 ( .ip1(\ANSWER/mem[5][5][9] ), .ip2(n9524), .s(n9965), .op(
        n2879) );
  mux2_1 U10685 ( .ip1(\ANSWER/mem[5][6][9] ), .ip2(n9524), .s(n9966), .op(
        n2878) );
  mux2_1 U10686 ( .ip1(\ANSWER/mem[5][7][9] ), .ip2(n9524), .s(n9967), .op(
        n2877) );
  mux2_1 U10687 ( .ip1(\ANSWER/mem[5][8][9] ), .ip2(n9524), .s(n9968), .op(
        n2876) );
  mux2_1 U10688 ( .ip1(\ANSWER/mem[5][9][9] ), .ip2(n9524), .s(n9969), .op(
        n2875) );
  mux2_1 U10689 ( .ip1(\ANSWER/mem[6][0][9] ), .ip2(n9524), .s(n9970), .op(
        n2874) );
  mux2_1 U10690 ( .ip1(\ANSWER/mem[6][1][9] ), .ip2(n9524), .s(n9971), .op(
        n2873) );
  mux2_1 U10691 ( .ip1(\ANSWER/mem[6][2][9] ), .ip2(n9524), .s(n9972), .op(
        n2872) );
  mux2_1 U10692 ( .ip1(\ANSWER/mem[6][3][9] ), .ip2(n9524), .s(n9973), .op(
        n2871) );
  mux2_1 U10693 ( .ip1(\ANSWER/mem[6][4][9] ), .ip2(n9524), .s(n9974), .op(
        n2870) );
  mux2_1 U10694 ( .ip1(\ANSWER/mem[6][5][9] ), .ip2(n9524), .s(n9975), .op(
        n2869) );
  mux2_1 U10695 ( .ip1(\ANSWER/mem[6][6][9] ), .ip2(n9524), .s(n9976), .op(
        n2868) );
  mux2_1 U10696 ( .ip1(\ANSWER/mem[6][7][9] ), .ip2(n9524), .s(n9977), .op(
        n2867) );
  mux2_1 U10697 ( .ip1(\ANSWER/mem[6][8][9] ), .ip2(n9524), .s(n9978), .op(
        n2866) );
  mux2_1 U10698 ( .ip1(\ANSWER/mem[6][9][9] ), .ip2(n9524), .s(n9979), .op(
        n2865) );
  mux2_1 U10699 ( .ip1(\ANSWER/mem[7][0][9] ), .ip2(n9524), .s(n9980), .op(
        n2864) );
  mux2_1 U10700 ( .ip1(\ANSWER/mem[7][1][9] ), .ip2(n9524), .s(n9981), .op(
        n2863) );
  mux2_1 U10701 ( .ip1(\ANSWER/mem[7][2][9] ), .ip2(n9524), .s(n9983), .op(
        n2862) );
  mux2_1 U10702 ( .ip1(\ANSWER/mem[7][3][9] ), .ip2(n9524), .s(n9984), .op(
        n2861) );
  mux2_1 U10703 ( .ip1(\ANSWER/mem[7][4][9] ), .ip2(n9524), .s(n9985), .op(
        n2860) );
  mux2_1 U10704 ( .ip1(\ANSWER/mem[7][5][9] ), .ip2(n9524), .s(n9986), .op(
        n2859) );
  mux2_1 U10705 ( .ip1(\ANSWER/mem[7][6][9] ), .ip2(n9524), .s(n9987), .op(
        n2858) );
  mux2_1 U10706 ( .ip1(\ANSWER/mem[7][7][9] ), .ip2(n9524), .s(n9988), .op(
        n2857) );
  mux2_1 U10707 ( .ip1(\ANSWER/mem[7][8][9] ), .ip2(n9524), .s(n9989), .op(
        n2856) );
  mux2_1 U10708 ( .ip1(\ANSWER/mem[7][9][9] ), .ip2(n9524), .s(n9990), .op(
        n2855) );
  mux2_1 U10709 ( .ip1(\ANSWER/mem[8][0][9] ), .ip2(n9524), .s(n9991), .op(
        n2854) );
  mux2_1 U10710 ( .ip1(\ANSWER/mem[8][1][9] ), .ip2(n9524), .s(n9992), .op(
        n2853) );
  mux2_1 U10711 ( .ip1(\ANSWER/mem[8][2][9] ), .ip2(n9524), .s(n9993), .op(
        n2852) );
  mux2_1 U10712 ( .ip1(\ANSWER/mem[8][3][9] ), .ip2(n9524), .s(n9994), .op(
        n2851) );
  mux2_1 U10713 ( .ip1(\ANSWER/mem[8][4][9] ), .ip2(n9525), .s(n9996), .op(
        n2850) );
  mux2_1 U10714 ( .ip1(\ANSWER/mem[8][5][9] ), .ip2(n9525), .s(n9997), .op(
        n2849) );
  mux2_1 U10715 ( .ip1(\ANSWER/mem[8][6][9] ), .ip2(n9525), .s(n9998), .op(
        n2848) );
  mux2_1 U10716 ( .ip1(\ANSWER/mem[8][7][9] ), .ip2(n9525), .s(n9999), .op(
        n2847) );
  mux2_1 U10717 ( .ip1(\ANSWER/mem[8][8][9] ), .ip2(n9525), .s(n10000), .op(
        n2846) );
  mux2_1 U10718 ( .ip1(\ANSWER/mem[8][9][9] ), .ip2(n9525), .s(n10001), .op(
        n2845) );
  mux2_1 U10719 ( .ip1(\ANSWER/mem[9][0][9] ), .ip2(n9525), .s(n10002), .op(
        n2844) );
  mux2_1 U10720 ( .ip1(\ANSWER/mem[9][1][9] ), .ip2(n9525), .s(n10003), .op(
        n2843) );
  mux2_1 U10721 ( .ip1(\ANSWER/mem[9][2][9] ), .ip2(n9525), .s(n10004), .op(
        n2842) );
  mux2_1 U10722 ( .ip1(\ANSWER/mem[9][3][9] ), .ip2(n9525), .s(n10005), .op(
        n2841) );
  mux2_1 U10723 ( .ip1(\ANSWER/mem[9][4][9] ), .ip2(n9525), .s(n10006), .op(
        n2840) );
  mux2_1 U10724 ( .ip1(\ANSWER/mem[9][5][9] ), .ip2(n9525), .s(n10007), .op(
        n2839) );
  mux2_1 U10725 ( .ip1(\ANSWER/mem[9][6][9] ), .ip2(n9523), .s(n10008), .op(
        n2838) );
  mux2_1 U10726 ( .ip1(\ANSWER/mem[9][7][9] ), .ip2(n9523), .s(n10009), .op(
        n2837) );
  mux2_1 U10727 ( .ip1(\ANSWER/mem[9][8][9] ), .ip2(n9524), .s(n10010), .op(
        n2836) );
  mux2_1 U10728 ( .ip1(\ANSWER/mem[9][9][9] ), .ip2(n9525), .s(n10011), .op(
        n2835) );
  fulladder U10729 ( .a(n9528), .b(n9527), .ci(n9526), .co(n9594), .s(n9519)
         );
  inv_1 U10730 ( .ip(q_w2[13]), .op(n9789) );
  nor2_1 U10731 ( .ip1(n9702), .ip2(n9789), .op(n9636) );
  nor2_1 U10732 ( .ip1(n9790), .ip2(n9864), .op(n9635) );
  nand2_1 U10733 ( .ip1(m2DataIn[15]), .ip2(q_w2[3]), .op(n9634) );
  inv_1 U10734 ( .ip(n9529), .op(n9599) );
  nand2_1 U10735 ( .ip1(m2DataIn[4]), .ip2(q_w2[14]), .op(n9627) );
  nor2_1 U10736 ( .ip1(n9530), .ip2(n9701), .op(n9626) );
  fulladder U10737 ( .a(n9600), .b(n9532), .ci(n9531), .co(n9597), .s(n9545)
         );
  fulladder U10738 ( .a(rdata[9]), .b(rdata[8]), .ci(n9533), .co(n9601), .s(
        n9458) );
  nand2_1 U10739 ( .ip1(q_w2[6]), .ip2(m2DataIn[12]), .op(n9535) );
  nor2_1 U10740 ( .ip1(n9703), .ip2(n9799), .op(n9534) );
  xor2_1 U10741 ( .ip1(n9535), .ip2(n9534), .op(n9602) );
  xor2_1 U10742 ( .ip1(n9601), .ip2(n9602), .op(n9621) );
  fulladder U10743 ( .a(n9538), .b(n9537), .ci(n9536), .co(n9539), .s(n9547)
         );
  inv_1 U10744 ( .ip(n9539), .op(n9620) );
  fulladder U10745 ( .a(n9542), .b(n9541), .ci(n9540), .co(n9619), .s(n9462)
         );
  fulladder U10746 ( .a(n9545), .b(n9544), .ci(n9543), .co(n9648), .s(n9580)
         );
  fulladder U10747 ( .a(n9548), .b(n9547), .ci(n9546), .co(n9549), .s(n9478)
         );
  inv_1 U10748 ( .ip(n9549), .op(n9653) );
  or2_1 U10749 ( .ip1(n9550), .ip2(n9551), .op(n9554) );
  or2_1 U10750 ( .ip1(n9552), .ip2(n9551), .op(n9553) );
  nand2_1 U10751 ( .ip1(n9554), .ip2(n9553), .op(n9618) );
  nand2_1 U10752 ( .ip1(q_w2[10]), .ip2(m2DataIn[8]), .op(n9556) );
  nand2_1 U10753 ( .ip1(q_w2[8]), .ip2(m2DataIn[10]), .op(n9555) );
  xor2_1 U10754 ( .ip1(n9556), .ip2(n9555), .op(n9613) );
  mux2_1 U10755 ( .ip1(n9557), .ip2(rdata[10]), .s(n9613), .op(n9617) );
  fulladder U10756 ( .a(n9560), .b(n9559), .ci(n9558), .co(n9616), .s(n9575)
         );
  or2_1 U10757 ( .ip1(n9561), .ip2(n9562), .op(n9565) );
  or2_1 U10758 ( .ip1(n9563), .ip2(n9562), .op(n9564) );
  nand2_1 U10759 ( .ip1(n9565), .ip2(n9564), .op(n9647) );
  nand2_1 U10760 ( .ip1(m2DataIn[11]), .ip2(q_w2[12]), .op(n9898) );
  nor2_1 U10761 ( .ip1(n9898), .ip2(n9566), .op(n9608) );
  or2_1 U10762 ( .ip1(n9694), .ip2(n9608), .op(n9569) );
  nand2_1 U10763 ( .ip1(m2DataIn[6]), .ip2(q_w2[12]), .op(n9567) );
  or2_1 U10764 ( .ip1(n9567), .ip2(n9608), .op(n9568) );
  nand2_1 U10765 ( .ip1(n9569), .ip2(n9568), .op(n9607) );
  nor2_1 U10766 ( .ip1(n9863), .ip2(n9638), .op(n9609) );
  xnor2_1 U10767 ( .ip1(n9607), .ip2(n9609), .op(n9646) );
  fulladder U10768 ( .a(n9572), .b(n9571), .ci(n9570), .co(n9645), .s(n9574)
         );
  fulladder U10769 ( .a(n9575), .b(n9574), .ci(n9573), .co(n9622), .s(n9578)
         );
  fulladder U10770 ( .a(n9578), .b(n9577), .ci(n9576), .co(n9651), .s(n9527)
         );
  fulladder U10771 ( .a(n9581), .b(n9580), .ci(n9579), .co(n9654), .s(n9528)
         );
  or2_1 U10772 ( .ip1(n9583), .ip2(n9582), .op(n9584) );
  nand2_1 U10773 ( .ip1(n9585), .ip2(n9584), .op(n9586) );
  nand2_1 U10774 ( .ip1(n9587), .ip2(n9586), .op(n9596) );
  or2_1 U10775 ( .ip1(n9587), .ip2(n9586), .op(n9593) );
  nand2_1 U10776 ( .ip1(n9596), .ip2(n9593), .op(n9589) );
  nor2_1 U10777 ( .ip1(n9594), .ip2(n9589), .op(n9588) );
  not_ab_or_c_or_d U10778 ( .ip1(n9594), .ip2(n9589), .ip3(n9907), .ip4(n9588), 
        .op(n9591) );
  buf_1 U10779 ( .ip(n9591), .op(n9590) );
  mux2_1 U10780 ( .ip1(\ANSWER/mem[0][0][10] ), .ip2(n9590), .s(n9910), .op(
        n2834) );
  mux2_1 U10781 ( .ip1(\ANSWER/mem[0][1][10] ), .ip2(n9590), .s(n9911), .op(
        n2833) );
  mux2_1 U10782 ( .ip1(\ANSWER/mem[0][2][10] ), .ip2(n9590), .s(n9912), .op(
        n2832) );
  mux2_1 U10783 ( .ip1(\ANSWER/mem[0][3][10] ), .ip2(n9590), .s(n9913), .op(
        n2831) );
  mux2_1 U10784 ( .ip1(\ANSWER/mem[0][4][10] ), .ip2(n9590), .s(n9914), .op(
        n2830) );
  mux2_1 U10785 ( .ip1(\ANSWER/mem[0][5][10] ), .ip2(n9590), .s(n9915), .op(
        n2829) );
  mux2_1 U10786 ( .ip1(\ANSWER/mem[0][6][10] ), .ip2(n9590), .s(n9916), .op(
        n2828) );
  mux2_1 U10787 ( .ip1(\ANSWER/mem[0][7][10] ), .ip2(n9590), .s(n9917), .op(
        n2827) );
  mux2_1 U10788 ( .ip1(\ANSWER/mem[0][8][10] ), .ip2(n9590), .s(n9918), .op(
        n2826) );
  mux2_1 U10789 ( .ip1(\ANSWER/mem[0][9][10] ), .ip2(n9590), .s(n9919), .op(
        n2825) );
  mux2_1 U10790 ( .ip1(\ANSWER/mem[1][0][10] ), .ip2(n9590), .s(n9920), .op(
        n2824) );
  mux2_1 U10791 ( .ip1(\ANSWER/mem[1][1][10] ), .ip2(n9590), .s(n9921), .op(
        n2823) );
  mux2_1 U10792 ( .ip1(\ANSWER/mem[1][2][10] ), .ip2(n9590), .s(n9922), .op(
        n2822) );
  mux2_1 U10793 ( .ip1(\ANSWER/mem[1][3][10] ), .ip2(n9590), .s(n9923), .op(
        n2821) );
  mux2_1 U10794 ( .ip1(\ANSWER/mem[1][4][10] ), .ip2(n9590), .s(n9924), .op(
        n2820) );
  mux2_1 U10795 ( .ip1(\ANSWER/mem[1][5][10] ), .ip2(n9590), .s(n9925), .op(
        n2819) );
  mux2_1 U10796 ( .ip1(\ANSWER/mem[1][6][10] ), .ip2(n9590), .s(n9926), .op(
        n2818) );
  mux2_1 U10797 ( .ip1(\ANSWER/mem[1][7][10] ), .ip2(n9590), .s(n9927), .op(
        n2817) );
  mux2_1 U10798 ( .ip1(\ANSWER/mem[1][8][10] ), .ip2(n9590), .s(n9928), .op(
        n2816) );
  mux2_1 U10799 ( .ip1(\ANSWER/mem[1][9][10] ), .ip2(n9590), .s(n9929), .op(
        n2815) );
  mux2_1 U10800 ( .ip1(\ANSWER/mem[2][0][10] ), .ip2(n9590), .s(n9930), .op(
        n2814) );
  mux2_1 U10801 ( .ip1(\ANSWER/mem[2][1][10] ), .ip2(n9590), .s(n9931), .op(
        n2813) );
  mux2_1 U10802 ( .ip1(\ANSWER/mem[2][2][10] ), .ip2(n9590), .s(n9932), .op(
        n2812) );
  mux2_1 U10803 ( .ip1(\ANSWER/mem[2][3][10] ), .ip2(n9590), .s(n9933), .op(
        n2811) );
  mux2_1 U10804 ( .ip1(\ANSWER/mem[2][4][10] ), .ip2(n9590), .s(n9934), .op(
        n2810) );
  mux2_1 U10805 ( .ip1(\ANSWER/mem[2][5][10] ), .ip2(n9590), .s(n9935), .op(
        n2809) );
  mux2_1 U10806 ( .ip1(\ANSWER/mem[2][6][10] ), .ip2(n9590), .s(n9936), .op(
        n2808) );
  mux2_1 U10807 ( .ip1(\ANSWER/mem[2][7][10] ), .ip2(n9590), .s(n9937), .op(
        n2807) );
  mux2_1 U10808 ( .ip1(\ANSWER/mem[2][8][10] ), .ip2(n9590), .s(n9938), .op(
        n2806) );
  mux2_1 U10809 ( .ip1(\ANSWER/mem[2][9][10] ), .ip2(n9590), .s(n9939), .op(
        n2805) );
  mux2_1 U10810 ( .ip1(\ANSWER/mem[3][0][10] ), .ip2(n9590), .s(n9940), .op(
        n2804) );
  mux2_1 U10811 ( .ip1(\ANSWER/mem[3][1][10] ), .ip2(n9590), .s(n9941), .op(
        n2803) );
  mux2_1 U10812 ( .ip1(\ANSWER/mem[3][2][10] ), .ip2(n9590), .s(n9942), .op(
        n2802) );
  mux2_1 U10813 ( .ip1(\ANSWER/mem[3][3][10] ), .ip2(n9590), .s(n9943), .op(
        n2801) );
  mux2_1 U10814 ( .ip1(\ANSWER/mem[3][4][10] ), .ip2(n9590), .s(n9944), .op(
        n2800) );
  mux2_1 U10815 ( .ip1(\ANSWER/mem[3][5][10] ), .ip2(n9590), .s(n9945), .op(
        n2799) );
  mux2_1 U10816 ( .ip1(\ANSWER/mem[3][6][10] ), .ip2(n9591), .s(n9946), .op(
        n2798) );
  mux2_1 U10817 ( .ip1(\ANSWER/mem[3][7][10] ), .ip2(n9591), .s(n9947), .op(
        n2797) );
  mux2_1 U10818 ( .ip1(\ANSWER/mem[3][8][10] ), .ip2(n9591), .s(n9948), .op(
        n2796) );
  mux2_1 U10819 ( .ip1(\ANSWER/mem[3][9][10] ), .ip2(n9591), .s(n9949), .op(
        n2795) );
  mux2_1 U10820 ( .ip1(\ANSWER/mem[4][0][10] ), .ip2(n9591), .s(n9950), .op(
        n2794) );
  mux2_1 U10821 ( .ip1(\ANSWER/mem[4][1][10] ), .ip2(n9591), .s(n9951), .op(
        n2793) );
  mux2_1 U10822 ( .ip1(\ANSWER/mem[4][2][10] ), .ip2(n9591), .s(n9952), .op(
        n2792) );
  mux2_1 U10823 ( .ip1(\ANSWER/mem[4][3][10] ), .ip2(n9591), .s(n9953), .op(
        n2791) );
  mux2_1 U10824 ( .ip1(\ANSWER/mem[4][4][10] ), .ip2(n9591), .s(n9954), .op(
        n2790) );
  mux2_1 U10825 ( .ip1(\ANSWER/mem[4][5][10] ), .ip2(n9591), .s(n9955), .op(
        n2789) );
  mux2_1 U10826 ( .ip1(\ANSWER/mem[4][6][10] ), .ip2(n9591), .s(n9956), .op(
        n2788) );
  mux2_1 U10827 ( .ip1(\ANSWER/mem[4][7][10] ), .ip2(n9592), .s(n9957), .op(
        n2787) );
  mux2_1 U10828 ( .ip1(\ANSWER/mem[4][8][10] ), .ip2(n9592), .s(n9958), .op(
        n2786) );
  mux2_1 U10829 ( .ip1(\ANSWER/mem[4][9][10] ), .ip2(n9592), .s(n9959), .op(
        n2785) );
  mux2_1 U10830 ( .ip1(\ANSWER/mem[5][0][10] ), .ip2(n9592), .s(n9960), .op(
        n2784) );
  mux2_1 U10831 ( .ip1(\ANSWER/mem[5][1][10] ), .ip2(n9592), .s(n9961), .op(
        n2783) );
  mux2_1 U10832 ( .ip1(\ANSWER/mem[5][2][10] ), .ip2(n9592), .s(n9962), .op(
        n2782) );
  mux2_1 U10833 ( .ip1(\ANSWER/mem[5][3][10] ), .ip2(n9592), .s(n9963), .op(
        n2781) );
  mux2_1 U10834 ( .ip1(\ANSWER/mem[5][4][10] ), .ip2(n9592), .s(n9964), .op(
        n2780) );
  mux2_1 U10835 ( .ip1(\ANSWER/mem[5][5][10] ), .ip2(n9592), .s(n9965), .op(
        n2779) );
  mux2_1 U10836 ( .ip1(\ANSWER/mem[5][6][10] ), .ip2(n9592), .s(n9966), .op(
        n2778) );
  mux2_1 U10837 ( .ip1(\ANSWER/mem[5][7][10] ), .ip2(n9591), .s(n9967), .op(
        n2777) );
  mux2_1 U10838 ( .ip1(\ANSWER/mem[5][8][10] ), .ip2(n9591), .s(n9968), .op(
        n2776) );
  mux2_1 U10839 ( .ip1(\ANSWER/mem[5][9][10] ), .ip2(n9591), .s(n9969), .op(
        n2775) );
  mux2_1 U10840 ( .ip1(\ANSWER/mem[6][0][10] ), .ip2(n9592), .s(n9970), .op(
        n2774) );
  mux2_1 U10841 ( .ip1(\ANSWER/mem[6][1][10] ), .ip2(n9591), .s(n9971), .op(
        n2773) );
  mux2_1 U10842 ( .ip1(\ANSWER/mem[6][2][10] ), .ip2(n9591), .s(n9972), .op(
        n2772) );
  mux2_1 U10843 ( .ip1(\ANSWER/mem[6][3][10] ), .ip2(n9591), .s(n9973), .op(
        n2771) );
  mux2_1 U10844 ( .ip1(\ANSWER/mem[6][4][10] ), .ip2(n9591), .s(n9974), .op(
        n2770) );
  mux2_1 U10845 ( .ip1(\ANSWER/mem[6][5][10] ), .ip2(n9591), .s(n9975), .op(
        n2769) );
  mux2_1 U10846 ( .ip1(\ANSWER/mem[6][6][10] ), .ip2(n9591), .s(n9976), .op(
        n2768) );
  mux2_1 U10847 ( .ip1(\ANSWER/mem[6][7][10] ), .ip2(n9591), .s(n9977), .op(
        n2767) );
  mux2_1 U10848 ( .ip1(\ANSWER/mem[6][8][10] ), .ip2(n9591), .s(n9978), .op(
        n2766) );
  mux2_1 U10849 ( .ip1(\ANSWER/mem[6][9][10] ), .ip2(n9591), .s(n9979), .op(
        n2765) );
  mux2_1 U10850 ( .ip1(\ANSWER/mem[7][0][10] ), .ip2(n9591), .s(n9980), .op(
        n2764) );
  mux2_1 U10851 ( .ip1(\ANSWER/mem[7][1][10] ), .ip2(n9591), .s(n9981), .op(
        n2763) );
  buf_1 U10852 ( .ip(n9591), .op(n9592) );
  mux2_1 U10853 ( .ip1(\ANSWER/mem[7][2][10] ), .ip2(n9592), .s(n9983), .op(
        n2762) );
  mux2_1 U10854 ( .ip1(\ANSWER/mem[7][3][10] ), .ip2(n9592), .s(n9984), .op(
        n2761) );
  mux2_1 U10855 ( .ip1(\ANSWER/mem[7][4][10] ), .ip2(n9592), .s(n9985), .op(
        n2760) );
  mux2_1 U10856 ( .ip1(\ANSWER/mem[7][5][10] ), .ip2(n9592), .s(n9986), .op(
        n2759) );
  mux2_1 U10857 ( .ip1(\ANSWER/mem[7][6][10] ), .ip2(n9592), .s(n9987), .op(
        n2758) );
  mux2_1 U10858 ( .ip1(\ANSWER/mem[7][7][10] ), .ip2(n9592), .s(n9988), .op(
        n2757) );
  mux2_1 U10859 ( .ip1(\ANSWER/mem[7][8][10] ), .ip2(n9592), .s(n9989), .op(
        n2756) );
  mux2_1 U10860 ( .ip1(\ANSWER/mem[7][9][10] ), .ip2(n9592), .s(n9990), .op(
        n2755) );
  mux2_1 U10861 ( .ip1(\ANSWER/mem[8][0][10] ), .ip2(n9591), .s(n9991), .op(
        n2754) );
  mux2_1 U10862 ( .ip1(\ANSWER/mem[8][1][10] ), .ip2(n9592), .s(n9992), .op(
        n2753) );
  mux2_1 U10863 ( .ip1(\ANSWER/mem[8][2][10] ), .ip2(n9592), .s(n9993), .op(
        n2752) );
  mux2_1 U10864 ( .ip1(\ANSWER/mem[8][3][10] ), .ip2(n9592), .s(n9994), .op(
        n2751) );
  mux2_1 U10865 ( .ip1(\ANSWER/mem[8][4][10] ), .ip2(n9591), .s(n9996), .op(
        n2750) );
  mux2_1 U10866 ( .ip1(\ANSWER/mem[8][5][10] ), .ip2(n9591), .s(n9997), .op(
        n2749) );
  mux2_1 U10867 ( .ip1(\ANSWER/mem[8][6][10] ), .ip2(n9591), .s(n9998), .op(
        n2748) );
  mux2_1 U10868 ( .ip1(\ANSWER/mem[8][7][10] ), .ip2(n9591), .s(n9999), .op(
        n2747) );
  mux2_1 U10869 ( .ip1(\ANSWER/mem[8][8][10] ), .ip2(n9591), .s(n10000), .op(
        n2746) );
  mux2_1 U10870 ( .ip1(\ANSWER/mem[8][9][10] ), .ip2(n9591), .s(n10001), .op(
        n2745) );
  mux2_1 U10871 ( .ip1(\ANSWER/mem[9][0][10] ), .ip2(n9591), .s(n10002), .op(
        n2744) );
  mux2_1 U10872 ( .ip1(\ANSWER/mem[9][1][10] ), .ip2(n9591), .s(n10003), .op(
        n2743) );
  mux2_1 U10873 ( .ip1(\ANSWER/mem[9][2][10] ), .ip2(n9591), .s(n10004), .op(
        n2742) );
  mux2_1 U10874 ( .ip1(\ANSWER/mem[9][3][10] ), .ip2(n9591), .s(n10005), .op(
        n2741) );
  mux2_1 U10875 ( .ip1(\ANSWER/mem[9][4][10] ), .ip2(n9591), .s(n10006), .op(
        n2740) );
  mux2_1 U10876 ( .ip1(\ANSWER/mem[9][5][10] ), .ip2(n9591), .s(n10007), .op(
        n2739) );
  mux2_1 U10877 ( .ip1(\ANSWER/mem[9][6][10] ), .ip2(n9592), .s(n10008), .op(
        n2738) );
  mux2_1 U10878 ( .ip1(\ANSWER/mem[9][7][10] ), .ip2(n9592), .s(n10009), .op(
        n2737) );
  mux2_1 U10879 ( .ip1(\ANSWER/mem[9][8][10] ), .ip2(n9592), .s(n10010), .op(
        n2736) );
  mux2_1 U10880 ( .ip1(\ANSWER/mem[9][9][10] ), .ip2(n9592), .s(n10011), .op(
        n2735) );
  nand2_1 U10881 ( .ip1(n9594), .ip2(n9593), .op(n9595) );
  nand2_1 U10882 ( .ip1(n9596), .ip2(n9595), .op(n9716) );
  fulladder U10883 ( .a(n9599), .b(n9598), .ci(n9597), .co(n9686), .s(n9650)
         );
  nand2_1 U10884 ( .ip1(m2DataIn[13]), .ip2(q_w2[6]), .op(n9706) );
  nor2_1 U10885 ( .ip1(n9706), .ip2(n9600), .op(n9603) );
  or2_1 U10886 ( .ip1(n9601), .ip2(n9603), .op(n9606) );
  inv_1 U10887 ( .ip(n9602), .op(n9604) );
  or2_1 U10888 ( .ip1(n9604), .ip2(n9603), .op(n9605) );
  nand2_1 U10889 ( .ip1(n9606), .ip2(n9605), .op(n9710) );
  or2_1 U10890 ( .ip1(n9607), .ip2(n9608), .op(n9611) );
  or2_1 U10891 ( .ip1(n9609), .ip2(n9608), .op(n9610) );
  nand2_1 U10892 ( .ip1(n9611), .ip2(n9610), .op(n9707) );
  nand2_1 U10893 ( .ip1(m2DataIn[10]), .ip2(q_w2[10]), .op(n9736) );
  nor3_1 U10894 ( .ip1(n9817), .ip2(n9788), .ip3(n9736), .op(n9612) );
  or2_1 U10895 ( .ip1(rdata[10]), .ip2(n9612), .op(n9615) );
  or2_1 U10896 ( .ip1(n9613), .ip2(n9612), .op(n9614) );
  nand2_1 U10897 ( .ip1(n9615), .ip2(n9614), .op(n9705) );
  fulladder U10898 ( .a(n9618), .b(n9617), .ci(n9616), .co(n9708), .s(n9624)
         );
  fulladder U10899 ( .a(n9621), .b(n9620), .ci(n9619), .co(n9684), .s(n9649)
         );
  fulladder U10900 ( .a(n9624), .b(n9623), .ci(n9622), .co(n9713), .s(n9652)
         );
  fulladder U10901 ( .a(n9627), .b(n9626), .ci(n9625), .co(n9628), .s(n9598)
         );
  inv_1 U10902 ( .ip(n9628), .op(n9679) );
  inv_1 U10903 ( .ip(rdata[11]), .op(n9633) );
  nand2_1 U10904 ( .ip1(m2DataIn[9]), .ip2(q_w2[10]), .op(n9629) );
  nor3_1 U10905 ( .ip1(n9790), .ip2(n9864), .ip3(n9736), .op(n9669) );
  or2_1 U10906 ( .ip1(n9629), .ip2(n9669), .op(n9632) );
  nand2_1 U10907 ( .ip1(m2DataIn[10]), .ip2(q_w2[9]), .op(n9630) );
  or2_1 U10908 ( .ip1(n9630), .ip2(n9669), .op(n9631) );
  nand2_1 U10909 ( .ip1(n9632), .ip2(n9631), .op(n9670) );
  mux2_1 U10910 ( .ip1(rdata[11]), .ip2(n9633), .s(n9670), .op(n9678) );
  fulladder U10911 ( .a(n9636), .b(n9635), .ci(n9634), .co(n9677), .s(n9529)
         );
  inv_1 U10912 ( .ip(n9637), .op(n9683) );
  nand2_1 U10913 ( .ip1(m2DataIn[6]), .ip2(q_w2[13]), .op(n9668) );
  nor2_1 U10914 ( .ip1(n9704), .ip2(n9638), .op(n9667) );
  nand2_1 U10915 ( .ip1(m2DataIn[8]), .ip2(q_w2[11]), .op(n9666) );
  inv_1 U10916 ( .ip(n9639), .op(n9676) );
  nor2_1 U10917 ( .ip1(n9640), .ip2(n9701), .op(n9700) );
  nand2_1 U10918 ( .ip1(m2DataIn[7]), .ip2(q_w2[12]), .op(n9699) );
  nand2_1 U10919 ( .ip1(m2DataIn[5]), .ip2(q_w2[14]), .op(n9698) );
  inv_1 U10920 ( .ip(n9641), .op(n9675) );
  nand2_1 U10921 ( .ip1(q_w2[7]), .ip2(m2DataIn[12]), .op(n9643) );
  nand2_1 U10922 ( .ip1(q_w2[8]), .ip2(m2DataIn[11]), .op(n9642) );
  xor2_1 U10923 ( .ip1(n9643), .ip2(n9642), .op(n9687) );
  nor2_1 U10924 ( .ip1(n9863), .ip2(n9703), .op(n9689) );
  xor2_1 U10925 ( .ip1(n9687), .ip2(n9689), .op(n9674) );
  inv_1 U10926 ( .ip(n9644), .op(n9682) );
  fulladder U10927 ( .a(n9647), .b(n9646), .ci(n9645), .co(n9681), .s(n9623)
         );
  fulladder U10928 ( .a(n9650), .b(n9649), .ci(n9648), .co(n9711), .s(n9656)
         );
  fulladder U10929 ( .a(n9653), .b(n9652), .ci(n9651), .co(n9661), .s(n9655)
         );
  fulladder U10930 ( .a(n9656), .b(n9655), .ci(n9654), .co(n9714), .s(n9587)
         );
  nor2_1 U10931 ( .ip1(n9907), .ip2(n9657), .op(n9659) );
  buf_1 U10932 ( .ip(n9659), .op(n9658) );
  mux2_1 U10933 ( .ip1(\ANSWER/mem[0][0][11] ), .ip2(n9658), .s(n9910), .op(
        n2734) );
  mux2_1 U10934 ( .ip1(\ANSWER/mem[0][1][11] ), .ip2(n9658), .s(n9911), .op(
        n2733) );
  mux2_1 U10935 ( .ip1(\ANSWER/mem[0][2][11] ), .ip2(n9658), .s(n9912), .op(
        n2732) );
  mux2_1 U10936 ( .ip1(\ANSWER/mem[0][3][11] ), .ip2(n9658), .s(n9913), .op(
        n2731) );
  mux2_1 U10937 ( .ip1(\ANSWER/mem[0][4][11] ), .ip2(n9658), .s(n9914), .op(
        n2730) );
  mux2_1 U10938 ( .ip1(\ANSWER/mem[0][5][11] ), .ip2(n9658), .s(n9915), .op(
        n2729) );
  mux2_1 U10939 ( .ip1(\ANSWER/mem[0][6][11] ), .ip2(n9658), .s(n9916), .op(
        n2728) );
  mux2_1 U10940 ( .ip1(\ANSWER/mem[0][7][11] ), .ip2(n9658), .s(n9917), .op(
        n2727) );
  mux2_1 U10941 ( .ip1(\ANSWER/mem[0][8][11] ), .ip2(n9658), .s(n9918), .op(
        n2726) );
  mux2_1 U10942 ( .ip1(\ANSWER/mem[0][9][11] ), .ip2(n9658), .s(n9919), .op(
        n2725) );
  mux2_1 U10943 ( .ip1(\ANSWER/mem[1][0][11] ), .ip2(n9658), .s(n9920), .op(
        n2724) );
  mux2_1 U10944 ( .ip1(\ANSWER/mem[1][1][11] ), .ip2(n9658), .s(n9921), .op(
        n2723) );
  mux2_1 U10945 ( .ip1(\ANSWER/mem[1][2][11] ), .ip2(n9658), .s(n9922), .op(
        n2722) );
  mux2_1 U10946 ( .ip1(\ANSWER/mem[1][3][11] ), .ip2(n9658), .s(n9923), .op(
        n2721) );
  mux2_1 U10947 ( .ip1(\ANSWER/mem[1][4][11] ), .ip2(n9658), .s(n9924), .op(
        n2720) );
  mux2_1 U10948 ( .ip1(\ANSWER/mem[1][5][11] ), .ip2(n9658), .s(n9925), .op(
        n2719) );
  mux2_1 U10949 ( .ip1(\ANSWER/mem[1][6][11] ), .ip2(n9658), .s(n9926), .op(
        n2718) );
  mux2_1 U10950 ( .ip1(\ANSWER/mem[1][7][11] ), .ip2(n9658), .s(n9927), .op(
        n2717) );
  mux2_1 U10951 ( .ip1(\ANSWER/mem[1][8][11] ), .ip2(n9658), .s(n9928), .op(
        n2716) );
  mux2_1 U10952 ( .ip1(\ANSWER/mem[1][9][11] ), .ip2(n9658), .s(n9929), .op(
        n2715) );
  mux2_1 U10953 ( .ip1(\ANSWER/mem[2][0][11] ), .ip2(n9658), .s(n9930), .op(
        n2714) );
  mux2_1 U10954 ( .ip1(\ANSWER/mem[2][1][11] ), .ip2(n9658), .s(n9931), .op(
        n2713) );
  mux2_1 U10955 ( .ip1(\ANSWER/mem[2][2][11] ), .ip2(n9658), .s(n9932), .op(
        n2712) );
  mux2_1 U10956 ( .ip1(\ANSWER/mem[2][3][11] ), .ip2(n9658), .s(n9933), .op(
        n2711) );
  mux2_1 U10957 ( .ip1(\ANSWER/mem[2][4][11] ), .ip2(n9658), .s(n9934), .op(
        n2710) );
  mux2_1 U10958 ( .ip1(\ANSWER/mem[2][5][11] ), .ip2(n9658), .s(n9935), .op(
        n2709) );
  mux2_1 U10959 ( .ip1(\ANSWER/mem[2][6][11] ), .ip2(n9658), .s(n9936), .op(
        n2708) );
  mux2_1 U10960 ( .ip1(\ANSWER/mem[2][7][11] ), .ip2(n9658), .s(n9937), .op(
        n2707) );
  mux2_1 U10961 ( .ip1(\ANSWER/mem[2][8][11] ), .ip2(n9658), .s(n9938), .op(
        n2706) );
  mux2_1 U10962 ( .ip1(\ANSWER/mem[2][9][11] ), .ip2(n9658), .s(n9939), .op(
        n2705) );
  mux2_1 U10963 ( .ip1(\ANSWER/mem[3][0][11] ), .ip2(n9658), .s(n9940), .op(
        n2704) );
  mux2_1 U10964 ( .ip1(\ANSWER/mem[3][1][11] ), .ip2(n9658), .s(n9941), .op(
        n2703) );
  mux2_1 U10965 ( .ip1(\ANSWER/mem[3][2][11] ), .ip2(n9658), .s(n9942), .op(
        n2702) );
  mux2_1 U10966 ( .ip1(\ANSWER/mem[3][3][11] ), .ip2(n9658), .s(n9943), .op(
        n2701) );
  mux2_1 U10967 ( .ip1(\ANSWER/mem[3][4][11] ), .ip2(n9658), .s(n9944), .op(
        n2700) );
  mux2_1 U10968 ( .ip1(\ANSWER/mem[3][5][11] ), .ip2(n9658), .s(n9945), .op(
        n2699) );
  mux2_1 U10969 ( .ip1(\ANSWER/mem[3][6][11] ), .ip2(n9659), .s(n9946), .op(
        n2698) );
  mux2_1 U10970 ( .ip1(\ANSWER/mem[3][7][11] ), .ip2(n9659), .s(n9947), .op(
        n2697) );
  mux2_1 U10971 ( .ip1(\ANSWER/mem[3][8][11] ), .ip2(n9659), .s(n9948), .op(
        n2696) );
  mux2_1 U10972 ( .ip1(\ANSWER/mem[3][9][11] ), .ip2(n9659), .s(n9949), .op(
        n2695) );
  mux2_1 U10973 ( .ip1(\ANSWER/mem[4][0][11] ), .ip2(n9659), .s(n9950), .op(
        n2694) );
  mux2_1 U10974 ( .ip1(\ANSWER/mem[4][1][11] ), .ip2(n9659), .s(n9951), .op(
        n2693) );
  mux2_1 U10975 ( .ip1(\ANSWER/mem[4][2][11] ), .ip2(n9659), .s(n9952), .op(
        n2692) );
  mux2_1 U10976 ( .ip1(\ANSWER/mem[4][3][11] ), .ip2(n9660), .s(n9953), .op(
        n2691) );
  mux2_1 U10977 ( .ip1(\ANSWER/mem[4][4][11] ), .ip2(n9660), .s(n9954), .op(
        n2690) );
  mux2_1 U10978 ( .ip1(\ANSWER/mem[4][5][11] ), .ip2(n9660), .s(n9955), .op(
        n2689) );
  mux2_1 U10979 ( .ip1(\ANSWER/mem[4][6][11] ), .ip2(n9660), .s(n9956), .op(
        n2688) );
  mux2_1 U10980 ( .ip1(\ANSWER/mem[4][7][11] ), .ip2(n9660), .s(n9957), .op(
        n2687) );
  mux2_1 U10981 ( .ip1(\ANSWER/mem[4][8][11] ), .ip2(n9660), .s(n9958), .op(
        n2686) );
  mux2_1 U10982 ( .ip1(\ANSWER/mem[4][9][11] ), .ip2(n9660), .s(n9959), .op(
        n2685) );
  mux2_1 U10983 ( .ip1(\ANSWER/mem[5][0][11] ), .ip2(n9660), .s(n9960), .op(
        n2684) );
  mux2_1 U10984 ( .ip1(\ANSWER/mem[5][1][11] ), .ip2(n9660), .s(n9961), .op(
        n2683) );
  mux2_1 U10985 ( .ip1(\ANSWER/mem[5][2][11] ), .ip2(n9660), .s(n9962), .op(
        n2682) );
  mux2_1 U10986 ( .ip1(\ANSWER/mem[5][3][11] ), .ip2(n9659), .s(n9963), .op(
        n2681) );
  mux2_1 U10987 ( .ip1(\ANSWER/mem[5][4][11] ), .ip2(n9660), .s(n9964), .op(
        n2680) );
  mux2_1 U10988 ( .ip1(\ANSWER/mem[5][5][11] ), .ip2(n9659), .s(n9965), .op(
        n2679) );
  mux2_1 U10989 ( .ip1(\ANSWER/mem[5][6][11] ), .ip2(n9659), .s(n9966), .op(
        n2678) );
  mux2_1 U10990 ( .ip1(\ANSWER/mem[5][7][11] ), .ip2(n9659), .s(n9967), .op(
        n2677) );
  mux2_1 U10991 ( .ip1(\ANSWER/mem[5][8][11] ), .ip2(n9659), .s(n9968), .op(
        n2676) );
  mux2_1 U10992 ( .ip1(\ANSWER/mem[5][9][11] ), .ip2(n9659), .s(n9969), .op(
        n2675) );
  mux2_1 U10993 ( .ip1(\ANSWER/mem[6][0][11] ), .ip2(n9659), .s(n9970), .op(
        n2674) );
  mux2_1 U10994 ( .ip1(\ANSWER/mem[6][1][11] ), .ip2(n9659), .s(n9971), .op(
        n2673) );
  mux2_1 U10995 ( .ip1(\ANSWER/mem[6][2][11] ), .ip2(n9659), .s(n9972), .op(
        n2672) );
  mux2_1 U10996 ( .ip1(\ANSWER/mem[6][3][11] ), .ip2(n9659), .s(n9973), .op(
        n2671) );
  mux2_1 U10997 ( .ip1(\ANSWER/mem[6][4][11] ), .ip2(n9659), .s(n9974), .op(
        n2670) );
  mux2_1 U10998 ( .ip1(\ANSWER/mem[6][5][11] ), .ip2(n9659), .s(n9975), .op(
        n2669) );
  mux2_1 U10999 ( .ip1(\ANSWER/mem[6][6][11] ), .ip2(n9659), .s(n9976), .op(
        n2668) );
  mux2_1 U11000 ( .ip1(\ANSWER/mem[6][7][11] ), .ip2(n9659), .s(n9977), .op(
        n2667) );
  mux2_1 U11001 ( .ip1(\ANSWER/mem[6][8][11] ), .ip2(n9659), .s(n9978), .op(
        n2666) );
  mux2_1 U11002 ( .ip1(\ANSWER/mem[6][9][11] ), .ip2(n9659), .s(n9979), .op(
        n2665) );
  mux2_1 U11003 ( .ip1(\ANSWER/mem[7][0][11] ), .ip2(n9659), .s(n9980), .op(
        n2664) );
  mux2_1 U11004 ( .ip1(\ANSWER/mem[7][1][11] ), .ip2(n9659), .s(n9981), .op(
        n2663) );
  buf_1 U11005 ( .ip(n9659), .op(n9660) );
  mux2_1 U11006 ( .ip1(\ANSWER/mem[7][2][11] ), .ip2(n9660), .s(n9983), .op(
        n2662) );
  mux2_1 U11007 ( .ip1(\ANSWER/mem[7][3][11] ), .ip2(n9660), .s(n9984), .op(
        n2661) );
  mux2_1 U11008 ( .ip1(\ANSWER/mem[7][4][11] ), .ip2(n9660), .s(n9985), .op(
        n2660) );
  mux2_1 U11009 ( .ip1(\ANSWER/mem[7][5][11] ), .ip2(n9660), .s(n9986), .op(
        n2659) );
  mux2_1 U11010 ( .ip1(\ANSWER/mem[7][6][11] ), .ip2(n9660), .s(n9987), .op(
        n2658) );
  mux2_1 U11011 ( .ip1(\ANSWER/mem[7][7][11] ), .ip2(n9660), .s(n9988), .op(
        n2657) );
  mux2_1 U11012 ( .ip1(\ANSWER/mem[7][8][11] ), .ip2(n9660), .s(n9989), .op(
        n2656) );
  mux2_1 U11013 ( .ip1(\ANSWER/mem[7][9][11] ), .ip2(n9660), .s(n9990), .op(
        n2655) );
  mux2_1 U11014 ( .ip1(\ANSWER/mem[8][0][11] ), .ip2(n9659), .s(n9991), .op(
        n2654) );
  mux2_1 U11015 ( .ip1(\ANSWER/mem[8][1][11] ), .ip2(n9660), .s(n9992), .op(
        n2653) );
  mux2_1 U11016 ( .ip1(\ANSWER/mem[8][2][11] ), .ip2(n9660), .s(n9993), .op(
        n2652) );
  mux2_1 U11017 ( .ip1(\ANSWER/mem[8][3][11] ), .ip2(n9660), .s(n9994), .op(
        n2651) );
  mux2_1 U11018 ( .ip1(\ANSWER/mem[8][4][11] ), .ip2(n9659), .s(n9996), .op(
        n2650) );
  mux2_1 U11019 ( .ip1(\ANSWER/mem[8][5][11] ), .ip2(n9659), .s(n9997), .op(
        n2649) );
  mux2_1 U11020 ( .ip1(\ANSWER/mem[8][6][11] ), .ip2(n9659), .s(n9998), .op(
        n2648) );
  mux2_1 U11021 ( .ip1(\ANSWER/mem[8][7][11] ), .ip2(n9659), .s(n9999), .op(
        n2647) );
  mux2_1 U11022 ( .ip1(\ANSWER/mem[8][8][11] ), .ip2(n9659), .s(n10000), .op(
        n2646) );
  mux2_1 U11023 ( .ip1(\ANSWER/mem[8][9][11] ), .ip2(n9659), .s(n10001), .op(
        n2645) );
  mux2_1 U11024 ( .ip1(\ANSWER/mem[9][0][11] ), .ip2(n9659), .s(n10002), .op(
        n2644) );
  mux2_1 U11025 ( .ip1(\ANSWER/mem[9][1][11] ), .ip2(n9659), .s(n10003), .op(
        n2643) );
  mux2_1 U11026 ( .ip1(\ANSWER/mem[9][2][11] ), .ip2(n9659), .s(n10004), .op(
        n2642) );
  mux2_1 U11027 ( .ip1(\ANSWER/mem[9][3][11] ), .ip2(n9659), .s(n10005), .op(
        n2641) );
  mux2_1 U11028 ( .ip1(\ANSWER/mem[9][4][11] ), .ip2(n9659), .s(n10006), .op(
        n2640) );
  mux2_1 U11029 ( .ip1(\ANSWER/mem[9][5][11] ), .ip2(n9659), .s(n10007), .op(
        n2639) );
  mux2_1 U11030 ( .ip1(\ANSWER/mem[9][6][11] ), .ip2(n9660), .s(n10008), .op(
        n2638) );
  mux2_1 U11031 ( .ip1(\ANSWER/mem[9][7][11] ), .ip2(n9660), .s(n10009), .op(
        n2637) );
  mux2_1 U11032 ( .ip1(\ANSWER/mem[9][8][11] ), .ip2(n9660), .s(n10010), .op(
        n2636) );
  mux2_1 U11033 ( .ip1(\ANSWER/mem[9][9][11] ), .ip2(n9660), .s(n10011), .op(
        n2635) );
  fulladder U11034 ( .a(n9663), .b(n9662), .ci(n9661), .co(n9777), .s(n9715)
         );
  nand2_1 U11035 ( .ip1(q_w2[11]), .ip2(m2DataIn[9]), .op(n9664) );
  nand2_1 U11036 ( .ip1(n9664), .ip2(n9736), .op(n9665) );
  nor2_1 U11037 ( .ip1(n9792), .ip2(n9791), .op(n9894) );
  nand3_1 U11038 ( .ip1(m2DataIn[9]), .ip2(q_w2[10]), .ip3(n9894), .op(n9752)
         );
  nand2_1 U11039 ( .ip1(n9665), .ip2(n9752), .op(n9753) );
  mux2_1 U11040 ( .ip1(rdata[12]), .ip2(n9754), .s(n9753), .op(n9760) );
  fulladder U11041 ( .a(n9668), .b(n9667), .ci(n9666), .co(n9759), .s(n9639)
         );
  or2_1 U11042 ( .ip1(rdata[11]), .ip2(n9669), .op(n9672) );
  or2_1 U11043 ( .ip1(n9670), .ip2(n9669), .op(n9671) );
  nand2_1 U11044 ( .ip1(n9672), .ip2(n9671), .op(n9758) );
  inv_1 U11045 ( .ip(n9673), .op(n9767) );
  fulladder U11046 ( .a(n9676), .b(n9675), .ci(n9674), .co(n9766), .s(n9644)
         );
  fulladder U11047 ( .a(n9679), .b(n9678), .ci(n9677), .co(n9765), .s(n9637)
         );
  inv_1 U11048 ( .ip(n9680), .op(n9774) );
  fulladder U11049 ( .a(n9683), .b(n9682), .ci(n9681), .co(n9773), .s(n9712)
         );
  fulladder U11050 ( .a(n9686), .b(n9685), .ci(n9684), .co(n9772), .s(n9663)
         );
  nand2_1 U11051 ( .ip1(m2DataIn[12]), .ip2(q_w2[8]), .op(n9744) );
  nor2_1 U11052 ( .ip1(n9694), .ip2(n9744), .op(n9688) );
  or2_1 U11053 ( .ip1(n9687), .ip2(n9688), .op(n9691) );
  or2_1 U11054 ( .ip1(n9689), .ip2(n9688), .op(n9690) );
  nand2_1 U11055 ( .ip1(n9691), .ip2(n9690), .op(n9763) );
  nor2_1 U11056 ( .ip1(n9863), .ip2(n9732), .op(n9697) );
  nand2_1 U11057 ( .ip1(q_w2[9]), .ip2(m2DataIn[11]), .op(n9693) );
  nand2_1 U11058 ( .ip1(m2DataIn[13]), .ip2(q_w2[7]), .op(n9692) );
  nand2_1 U11059 ( .ip1(n9693), .ip2(n9692), .op(n9696) );
  nor3_1 U11060 ( .ip1(n9799), .ip2(n9864), .ip3(n9694), .op(n9734) );
  inv_1 U11061 ( .ip(n9734), .op(n9695) );
  nand2_1 U11062 ( .ip1(n9696), .ip2(n9695), .op(n9731) );
  xor2_1 U11063 ( .ip1(n9697), .ip2(n9731), .op(n9762) );
  fulladder U11064 ( .a(n9700), .b(n9699), .ci(n9698), .co(n9761), .s(n9641)
         );
  nor2_1 U11065 ( .ip1(n9702), .ip2(n9701), .op(n9730) );
  nand2_1 U11066 ( .ip1(m2DataIn[6]), .ip2(q_w2[14]), .op(n9729) );
  nand2_1 U11067 ( .ip1(m2DataIn[8]), .ip2(q_w2[12]), .op(n9728) );
  nor2_1 U11068 ( .ip1(n9704), .ip2(n9703), .op(n9745) );
  nand2_1 U11069 ( .ip1(m2DataIn[7]), .ip2(q_w2[13]), .op(n9743) );
  fulladder U11070 ( .a(n9707), .b(n9706), .ci(n9705), .co(n9746), .s(n9709)
         );
  fulladder U11071 ( .a(n9710), .b(n9709), .ci(n9708), .co(n9769), .s(n9685)
         );
  fulladder U11072 ( .a(n9713), .b(n9712), .ci(n9711), .co(n9721), .s(n9662)
         );
  fulladder U11073 ( .a(n9716), .b(n9715), .ci(n9714), .co(n9775), .s(n9657)
         );
  nor2_1 U11074 ( .ip1(n9907), .ip2(n9717), .op(n9718) );
  buf_1 U11075 ( .ip(n9718), .op(n9719) );
  mux2_1 U11076 ( .ip1(\ANSWER/mem[0][0][12] ), .ip2(n9719), .s(n9910), .op(
        n2634) );
  mux2_1 U11077 ( .ip1(\ANSWER/mem[0][1][12] ), .ip2(n9719), .s(n9911), .op(
        n2633) );
  mux2_1 U11078 ( .ip1(\ANSWER/mem[0][2][12] ), .ip2(n9719), .s(n9912), .op(
        n2632) );
  mux2_1 U11079 ( .ip1(\ANSWER/mem[0][3][12] ), .ip2(n9719), .s(n9913), .op(
        n2631) );
  mux2_1 U11080 ( .ip1(\ANSWER/mem[0][4][12] ), .ip2(n9719), .s(n9914), .op(
        n2630) );
  mux2_1 U11081 ( .ip1(\ANSWER/mem[0][5][12] ), .ip2(n9719), .s(n9915), .op(
        n2629) );
  mux2_1 U11082 ( .ip1(\ANSWER/mem[0][6][12] ), .ip2(n9719), .s(n9916), .op(
        n2628) );
  mux2_1 U11083 ( .ip1(\ANSWER/mem[0][7][12] ), .ip2(n9719), .s(n9917), .op(
        n2627) );
  mux2_1 U11084 ( .ip1(\ANSWER/mem[0][8][12] ), .ip2(n9719), .s(n9918), .op(
        n2626) );
  mux2_1 U11085 ( .ip1(\ANSWER/mem[0][9][12] ), .ip2(n9719), .s(n9919), .op(
        n2625) );
  mux2_1 U11086 ( .ip1(\ANSWER/mem[1][0][12] ), .ip2(n9719), .s(n9920), .op(
        n2624) );
  mux2_1 U11087 ( .ip1(\ANSWER/mem[1][1][12] ), .ip2(n9719), .s(n9921), .op(
        n2623) );
  mux2_1 U11088 ( .ip1(\ANSWER/mem[1][2][12] ), .ip2(n9718), .s(n9922), .op(
        n2622) );
  mux2_1 U11089 ( .ip1(\ANSWER/mem[1][3][12] ), .ip2(n9718), .s(n9923), .op(
        n2621) );
  mux2_1 U11090 ( .ip1(\ANSWER/mem[1][4][12] ), .ip2(n9718), .s(n9924), .op(
        n2620) );
  mux2_1 U11091 ( .ip1(\ANSWER/mem[1][5][12] ), .ip2(n9718), .s(n9925), .op(
        n2619) );
  mux2_1 U11092 ( .ip1(\ANSWER/mem[1][6][12] ), .ip2(n9718), .s(n9926), .op(
        n2618) );
  mux2_1 U11093 ( .ip1(\ANSWER/mem[1][7][12] ), .ip2(n9718), .s(n9927), .op(
        n2617) );
  mux2_1 U11094 ( .ip1(\ANSWER/mem[1][8][12] ), .ip2(n9718), .s(n9928), .op(
        n2616) );
  mux2_1 U11095 ( .ip1(\ANSWER/mem[1][9][12] ), .ip2(n9718), .s(n9929), .op(
        n2615) );
  mux2_1 U11096 ( .ip1(\ANSWER/mem[2][0][12] ), .ip2(n9718), .s(n9930), .op(
        n2614) );
  mux2_1 U11097 ( .ip1(\ANSWER/mem[2][1][12] ), .ip2(n9718), .s(n9931), .op(
        n2613) );
  mux2_1 U11098 ( .ip1(\ANSWER/mem[2][2][12] ), .ip2(n9718), .s(n9932), .op(
        n2612) );
  mux2_1 U11099 ( .ip1(\ANSWER/mem[2][3][12] ), .ip2(n9718), .s(n9933), .op(
        n2611) );
  buf_1 U11100 ( .ip(n9718), .op(n9720) );
  mux2_1 U11101 ( .ip1(\ANSWER/mem[2][4][12] ), .ip2(n9720), .s(n9934), .op(
        n2610) );
  mux2_1 U11102 ( .ip1(\ANSWER/mem[2][5][12] ), .ip2(n9720), .s(n9935), .op(
        n2609) );
  mux2_1 U11103 ( .ip1(\ANSWER/mem[2][6][12] ), .ip2(n9719), .s(n9936), .op(
        n2608) );
  mux2_1 U11104 ( .ip1(\ANSWER/mem[2][7][12] ), .ip2(n9718), .s(n9937), .op(
        n2607) );
  mux2_1 U11105 ( .ip1(\ANSWER/mem[2][8][12] ), .ip2(n9718), .s(n9938), .op(
        n2606) );
  mux2_1 U11106 ( .ip1(\ANSWER/mem[2][9][12] ), .ip2(n9718), .s(n9939), .op(
        n2605) );
  mux2_1 U11107 ( .ip1(\ANSWER/mem[3][0][12] ), .ip2(n9718), .s(n9940), .op(
        n2604) );
  mux2_1 U11108 ( .ip1(\ANSWER/mem[3][1][12] ), .ip2(n9718), .s(n9941), .op(
        n2603) );
  mux2_1 U11109 ( .ip1(\ANSWER/mem[3][2][12] ), .ip2(n9718), .s(n9942), .op(
        n2602) );
  mux2_1 U11110 ( .ip1(\ANSWER/mem[3][3][12] ), .ip2(n9718), .s(n9943), .op(
        n2601) );
  mux2_1 U11111 ( .ip1(\ANSWER/mem[3][4][12] ), .ip2(n9718), .s(n9944), .op(
        n2600) );
  mux2_1 U11112 ( .ip1(\ANSWER/mem[3][5][12] ), .ip2(n9718), .s(n9945), .op(
        n2599) );
  mux2_1 U11113 ( .ip1(\ANSWER/mem[3][6][12] ), .ip2(n9720), .s(n9946), .op(
        n2598) );
  mux2_1 U11114 ( .ip1(\ANSWER/mem[3][7][12] ), .ip2(n9719), .s(n9947), .op(
        n2597) );
  mux2_1 U11115 ( .ip1(\ANSWER/mem[3][8][12] ), .ip2(n9720), .s(n9948), .op(
        n2596) );
  mux2_1 U11116 ( .ip1(\ANSWER/mem[3][9][12] ), .ip2(n9718), .s(n9949), .op(
        n2595) );
  mux2_1 U11117 ( .ip1(\ANSWER/mem[4][0][12] ), .ip2(n9719), .s(n9950), .op(
        n2594) );
  mux2_1 U11118 ( .ip1(\ANSWER/mem[4][1][12] ), .ip2(n9720), .s(n9951), .op(
        n2593) );
  mux2_1 U11119 ( .ip1(\ANSWER/mem[4][2][12] ), .ip2(n9718), .s(n9952), .op(
        n2592) );
  mux2_1 U11120 ( .ip1(\ANSWER/mem[4][3][12] ), .ip2(n9720), .s(n9953), .op(
        n2591) );
  mux2_1 U11121 ( .ip1(\ANSWER/mem[4][4][12] ), .ip2(n9720), .s(n9954), .op(
        n2590) );
  mux2_1 U11122 ( .ip1(\ANSWER/mem[4][5][12] ), .ip2(n9719), .s(n9955), .op(
        n2589) );
  mux2_1 U11123 ( .ip1(\ANSWER/mem[4][6][12] ), .ip2(n9719), .s(n9956), .op(
        n2588) );
  mux2_1 U11124 ( .ip1(\ANSWER/mem[4][7][12] ), .ip2(n9720), .s(n9957), .op(
        n2587) );
  mux2_1 U11125 ( .ip1(\ANSWER/mem[4][8][12] ), .ip2(n9718), .s(n9958), .op(
        n2586) );
  mux2_1 U11126 ( .ip1(\ANSWER/mem[4][9][12] ), .ip2(n9720), .s(n9959), .op(
        n2585) );
  mux2_1 U11127 ( .ip1(\ANSWER/mem[5][0][12] ), .ip2(n9720), .s(n9960), .op(
        n2584) );
  mux2_1 U11128 ( .ip1(\ANSWER/mem[5][1][12] ), .ip2(n9720), .s(n9961), .op(
        n2583) );
  mux2_1 U11129 ( .ip1(\ANSWER/mem[5][2][12] ), .ip2(n9720), .s(n9962), .op(
        n2582) );
  mux2_1 U11130 ( .ip1(\ANSWER/mem[5][3][12] ), .ip2(n9720), .s(n9963), .op(
        n2581) );
  mux2_1 U11131 ( .ip1(\ANSWER/mem[5][4][12] ), .ip2(n9720), .s(n9964), .op(
        n2580) );
  mux2_1 U11132 ( .ip1(\ANSWER/mem[5][5][12] ), .ip2(n9720), .s(n9965), .op(
        n2579) );
  mux2_1 U11133 ( .ip1(\ANSWER/mem[5][6][12] ), .ip2(n9720), .s(n9966), .op(
        n2578) );
  mux2_1 U11134 ( .ip1(\ANSWER/mem[5][7][12] ), .ip2(n9720), .s(n9967), .op(
        n2577) );
  mux2_1 U11135 ( .ip1(\ANSWER/mem[5][8][12] ), .ip2(n9719), .s(n9968), .op(
        n2576) );
  mux2_1 U11136 ( .ip1(\ANSWER/mem[5][9][12] ), .ip2(n9718), .s(n9969), .op(
        n2575) );
  mux2_1 U11137 ( .ip1(\ANSWER/mem[6][0][12] ), .ip2(n9718), .s(n9970), .op(
        n2574) );
  mux2_1 U11138 ( .ip1(\ANSWER/mem[6][1][12] ), .ip2(n9718), .s(n9971), .op(
        n2573) );
  mux2_1 U11139 ( .ip1(\ANSWER/mem[6][2][12] ), .ip2(n9718), .s(n9972), .op(
        n2572) );
  mux2_1 U11140 ( .ip1(\ANSWER/mem[6][3][12] ), .ip2(n9720), .s(n9973), .op(
        n2571) );
  mux2_1 U11141 ( .ip1(\ANSWER/mem[6][4][12] ), .ip2(n9719), .s(n9974), .op(
        n2570) );
  mux2_1 U11142 ( .ip1(\ANSWER/mem[6][5][12] ), .ip2(n9720), .s(n9975), .op(
        n2569) );
  mux2_1 U11143 ( .ip1(\ANSWER/mem[6][6][12] ), .ip2(n9719), .s(n9976), .op(
        n2568) );
  mux2_1 U11144 ( .ip1(\ANSWER/mem[6][7][12] ), .ip2(n9718), .s(n9977), .op(
        n2567) );
  mux2_1 U11145 ( .ip1(\ANSWER/mem[6][8][12] ), .ip2(n9720), .s(n9978), .op(
        n2566) );
  mux2_1 U11146 ( .ip1(\ANSWER/mem[6][9][12] ), .ip2(n9719), .s(n9979), .op(
        n2565) );
  mux2_1 U11147 ( .ip1(\ANSWER/mem[7][0][12] ), .ip2(n9718), .s(n9980), .op(
        n2564) );
  mux2_1 U11148 ( .ip1(\ANSWER/mem[7][1][12] ), .ip2(n9718), .s(n9981), .op(
        n2563) );
  mux2_1 U11149 ( .ip1(\ANSWER/mem[7][2][12] ), .ip2(n9718), .s(n9983), .op(
        n2562) );
  mux2_1 U11150 ( .ip1(\ANSWER/mem[7][3][12] ), .ip2(n9719), .s(n9984), .op(
        n2561) );
  mux2_1 U11151 ( .ip1(\ANSWER/mem[7][4][12] ), .ip2(n9719), .s(n9985), .op(
        n2560) );
  mux2_1 U11152 ( .ip1(\ANSWER/mem[7][5][12] ), .ip2(n9720), .s(n9986), .op(
        n2559) );
  mux2_1 U11153 ( .ip1(\ANSWER/mem[7][6][12] ), .ip2(n9720), .s(n9987), .op(
        n2558) );
  mux2_1 U11154 ( .ip1(\ANSWER/mem[7][7][12] ), .ip2(n9720), .s(n9988), .op(
        n2557) );
  mux2_1 U11155 ( .ip1(\ANSWER/mem[7][8][12] ), .ip2(n9719), .s(n9989), .op(
        n2556) );
  mux2_1 U11156 ( .ip1(\ANSWER/mem[7][9][12] ), .ip2(n9718), .s(n9990), .op(
        n2555) );
  mux2_1 U11157 ( .ip1(\ANSWER/mem[8][0][12] ), .ip2(n9718), .s(n9991), .op(
        n2554) );
  mux2_1 U11158 ( .ip1(\ANSWER/mem[8][1][12] ), .ip2(n9718), .s(n9992), .op(
        n2553) );
  mux2_1 U11159 ( .ip1(\ANSWER/mem[8][2][12] ), .ip2(n9719), .s(n9993), .op(
        n2552) );
  mux2_1 U11160 ( .ip1(\ANSWER/mem[8][3][12] ), .ip2(n9720), .s(n9994), .op(
        n2551) );
  mux2_1 U11161 ( .ip1(\ANSWER/mem[8][4][12] ), .ip2(n9718), .s(n9996), .op(
        n2550) );
  mux2_1 U11162 ( .ip1(\ANSWER/mem[8][5][12] ), .ip2(n9718), .s(n9997), .op(
        n2549) );
  mux2_1 U11163 ( .ip1(\ANSWER/mem[8][6][12] ), .ip2(n9718), .s(n9998), .op(
        n2548) );
  mux2_1 U11164 ( .ip1(\ANSWER/mem[8][7][12] ), .ip2(n9718), .s(n9999), .op(
        n2547) );
  mux2_1 U11165 ( .ip1(\ANSWER/mem[8][8][12] ), .ip2(n9720), .s(n10000), .op(
        n2546) );
  mux2_1 U11166 ( .ip1(\ANSWER/mem[8][9][12] ), .ip2(n9719), .s(n10001), .op(
        n2545) );
  mux2_1 U11167 ( .ip1(\ANSWER/mem[9][0][12] ), .ip2(n9719), .s(n10002), .op(
        n2544) );
  mux2_1 U11168 ( .ip1(\ANSWER/mem[9][1][12] ), .ip2(n9719), .s(n10003), .op(
        n2543) );
  mux2_1 U11169 ( .ip1(\ANSWER/mem[9][2][12] ), .ip2(n9720), .s(n10004), .op(
        n2542) );
  mux2_1 U11170 ( .ip1(\ANSWER/mem[9][3][12] ), .ip2(n9719), .s(n10005), .op(
        n2541) );
  mux2_1 U11171 ( .ip1(\ANSWER/mem[9][4][12] ), .ip2(n9720), .s(n10006), .op(
        n2540) );
  mux2_1 U11172 ( .ip1(\ANSWER/mem[9][5][12] ), .ip2(n9719), .s(n10007), .op(
        n2539) );
  mux2_1 U11173 ( .ip1(\ANSWER/mem[9][6][12] ), .ip2(n9720), .s(n10008), .op(
        n2538) );
  mux2_1 U11174 ( .ip1(\ANSWER/mem[9][7][12] ), .ip2(n9720), .s(n10009), .op(
        n2537) );
  mux2_1 U11175 ( .ip1(\ANSWER/mem[9][8][12] ), .ip2(n9720), .s(n10010), .op(
        n2536) );
  mux2_1 U11176 ( .ip1(\ANSWER/mem[9][9][12] ), .ip2(n9720), .s(n10011), .op(
        n2535) );
  fulladder U11177 ( .a(n9723), .b(n9722), .ci(n9721), .co(n9834), .s(n9776)
         );
  nor2_1 U11178 ( .ip1(n9790), .ip2(n9724), .op(n9805) );
  nor2_1 U11179 ( .ip1(n9725), .ip2(n9816), .op(n9804) );
  nand2_1 U11180 ( .ip1(m2DataIn[15]), .ip2(q_w2[6]), .op(n9803) );
  inv_1 U11181 ( .ip(n9726), .op(n9809) );
  nor2_1 U11182 ( .ip1(n9815), .ip2(n9864), .op(n9787) );
  nor2_1 U11183 ( .ip1(n9817), .ip2(n9789), .op(n9786) );
  nand2_1 U11184 ( .ip1(m2DataIn[6]), .ip2(q_w2[15]), .op(n9785) );
  inv_1 U11185 ( .ip(n9727), .op(n9808) );
  fulladder U11186 ( .a(n9730), .b(n9729), .ci(n9728), .co(n9807), .s(n9748)
         );
  nor3_1 U11187 ( .ip1(n9863), .ip2(n9732), .ip3(n9731), .op(n9733) );
  nor2_1 U11188 ( .ip1(n9734), .ip2(n9733), .op(n9821) );
  nor2_1 U11189 ( .ip1(n9735), .ip2(n9791), .op(n9793) );
  inv_1 U11190 ( .ip(n9736), .op(n9737) );
  nand2_1 U11191 ( .ip1(n9793), .ip2(n9737), .op(n9802) );
  inv_1 U11192 ( .ip(n9802), .op(n9741) );
  or2_1 U11193 ( .ip1(q_w2[10]), .ip2(n9894), .op(n9739) );
  or2_1 U11194 ( .ip1(m2DataIn[11]), .ip2(n9894), .op(n9738) );
  nand2_1 U11195 ( .ip1(n9739), .ip2(n9738), .op(n9740) );
  nor2_1 U11196 ( .ip1(n9741), .ip2(n9740), .op(n9800) );
  mux2_1 U11197 ( .ip1(n9742), .ip2(rdata[13]), .s(n9800), .op(n9820) );
  fulladder U11198 ( .a(n9745), .b(n9744), .ci(n9743), .co(n9819), .s(n9747)
         );
  fulladder U11199 ( .a(n9748), .b(n9747), .ci(n9746), .co(n9829), .s(n9770)
         );
  inv_1 U11200 ( .ip(n9749), .op(n9827) );
  nand2_1 U11201 ( .ip1(q_w2[7]), .ip2(m2DataIn[14]), .op(n9751) );
  nor2_1 U11202 ( .ip1(n9799), .ip2(n9788), .op(n9750) );
  xor2_1 U11203 ( .ip1(n9751), .ip2(n9750), .op(n9810) );
  inv_1 U11204 ( .ip(n9810), .op(n9757) );
  inv_1 U11205 ( .ip(n9752), .op(n9756) );
  nor2_1 U11206 ( .ip1(n9754), .ip2(n9753), .op(n9755) );
  nor2_1 U11207 ( .ip1(n9756), .ip2(n9755), .op(n9811) );
  mux2_1 U11208 ( .ip1(n9757), .ip2(n9810), .s(n9811), .op(n9824) );
  fulladder U11209 ( .a(n9760), .b(n9759), .ci(n9758), .co(n9823), .s(n9673)
         );
  fulladder U11210 ( .a(n9763), .b(n9762), .ci(n9761), .co(n9822), .s(n9771)
         );
  inv_1 U11211 ( .ip(n9764), .op(n9826) );
  fulladder U11212 ( .a(n9767), .b(n9766), .ci(n9765), .co(n9825), .s(n9680)
         );
  inv_1 U11213 ( .ip(n9768), .op(n9784) );
  fulladder U11214 ( .a(n9771), .b(n9770), .ci(n9769), .co(n9783), .s(n9722)
         );
  fulladder U11215 ( .a(n9774), .b(n9773), .ci(n9772), .co(n9782), .s(n9723)
         );
  fulladder U11216 ( .a(n9777), .b(n9776), .ci(n9775), .co(n9832), .s(n9717)
         );
  nor2_1 U11217 ( .ip1(n9907), .ip2(n9778), .op(n9780) );
  buf_1 U11218 ( .ip(n9780), .op(n9779) );
  mux2_1 U11219 ( .ip1(\ANSWER/mem[0][0][13] ), .ip2(n9779), .s(n9910), .op(
        n2534) );
  mux2_1 U11220 ( .ip1(\ANSWER/mem[0][1][13] ), .ip2(n9779), .s(n9911), .op(
        n2533) );
  mux2_1 U11221 ( .ip1(\ANSWER/mem[0][2][13] ), .ip2(n9779), .s(n9912), .op(
        n2532) );
  mux2_1 U11222 ( .ip1(\ANSWER/mem[0][3][13] ), .ip2(n9779), .s(n9913), .op(
        n2531) );
  mux2_1 U11223 ( .ip1(\ANSWER/mem[0][4][13] ), .ip2(n9779), .s(n9914), .op(
        n2530) );
  mux2_1 U11224 ( .ip1(\ANSWER/mem[0][5][13] ), .ip2(n9779), .s(n9915), .op(
        n2529) );
  mux2_1 U11225 ( .ip1(\ANSWER/mem[0][6][13] ), .ip2(n9779), .s(n9916), .op(
        n2528) );
  mux2_1 U11226 ( .ip1(\ANSWER/mem[0][7][13] ), .ip2(n9779), .s(n9917), .op(
        n2527) );
  mux2_1 U11227 ( .ip1(\ANSWER/mem[0][8][13] ), .ip2(n9779), .s(n9918), .op(
        n2526) );
  mux2_1 U11228 ( .ip1(\ANSWER/mem[0][9][13] ), .ip2(n9779), .s(n9919), .op(
        n2525) );
  mux2_1 U11229 ( .ip1(\ANSWER/mem[1][0][13] ), .ip2(n9779), .s(n9920), .op(
        n2524) );
  mux2_1 U11230 ( .ip1(\ANSWER/mem[1][1][13] ), .ip2(n9779), .s(n9921), .op(
        n2523) );
  mux2_1 U11231 ( .ip1(\ANSWER/mem[1][2][13] ), .ip2(n9779), .s(n9922), .op(
        n2522) );
  mux2_1 U11232 ( .ip1(\ANSWER/mem[1][3][13] ), .ip2(n9779), .s(n9923), .op(
        n2521) );
  mux2_1 U11233 ( .ip1(\ANSWER/mem[1][4][13] ), .ip2(n9779), .s(n9924), .op(
        n2520) );
  mux2_1 U11234 ( .ip1(\ANSWER/mem[1][5][13] ), .ip2(n9779), .s(n9925), .op(
        n2519) );
  mux2_1 U11235 ( .ip1(\ANSWER/mem[1][6][13] ), .ip2(n9779), .s(n9926), .op(
        n2518) );
  mux2_1 U11236 ( .ip1(\ANSWER/mem[1][7][13] ), .ip2(n9779), .s(n9927), .op(
        n2517) );
  mux2_1 U11237 ( .ip1(\ANSWER/mem[1][8][13] ), .ip2(n9779), .s(n9928), .op(
        n2516) );
  mux2_1 U11238 ( .ip1(\ANSWER/mem[1][9][13] ), .ip2(n9779), .s(n9929), .op(
        n2515) );
  mux2_1 U11239 ( .ip1(\ANSWER/mem[2][0][13] ), .ip2(n9779), .s(n9930), .op(
        n2514) );
  mux2_1 U11240 ( .ip1(\ANSWER/mem[2][1][13] ), .ip2(n9779), .s(n9931), .op(
        n2513) );
  mux2_1 U11241 ( .ip1(\ANSWER/mem[2][2][13] ), .ip2(n9779), .s(n9932), .op(
        n2512) );
  mux2_1 U11242 ( .ip1(\ANSWER/mem[2][3][13] ), .ip2(n9779), .s(n9933), .op(
        n2511) );
  mux2_1 U11243 ( .ip1(\ANSWER/mem[2][4][13] ), .ip2(n9779), .s(n9934), .op(
        n2510) );
  mux2_1 U11244 ( .ip1(\ANSWER/mem[2][5][13] ), .ip2(n9779), .s(n9935), .op(
        n2509) );
  mux2_1 U11245 ( .ip1(\ANSWER/mem[2][6][13] ), .ip2(n9779), .s(n9936), .op(
        n2508) );
  mux2_1 U11246 ( .ip1(\ANSWER/mem[2][7][13] ), .ip2(n9779), .s(n9937), .op(
        n2507) );
  mux2_1 U11247 ( .ip1(\ANSWER/mem[2][8][13] ), .ip2(n9779), .s(n9938), .op(
        n2506) );
  mux2_1 U11248 ( .ip1(\ANSWER/mem[2][9][13] ), .ip2(n9779), .s(n9939), .op(
        n2505) );
  mux2_1 U11249 ( .ip1(\ANSWER/mem[3][0][13] ), .ip2(n9779), .s(n9940), .op(
        n2504) );
  mux2_1 U11250 ( .ip1(\ANSWER/mem[3][1][13] ), .ip2(n9779), .s(n9941), .op(
        n2503) );
  mux2_1 U11251 ( .ip1(\ANSWER/mem[3][2][13] ), .ip2(n9779), .s(n9942), .op(
        n2502) );
  mux2_1 U11252 ( .ip1(\ANSWER/mem[3][3][13] ), .ip2(n9779), .s(n9943), .op(
        n2501) );
  mux2_1 U11253 ( .ip1(\ANSWER/mem[3][4][13] ), .ip2(n9779), .s(n9944), .op(
        n2500) );
  mux2_1 U11254 ( .ip1(\ANSWER/mem[3][5][13] ), .ip2(n9779), .s(n9945), .op(
        n2499) );
  mux2_1 U11255 ( .ip1(\ANSWER/mem[3][6][13] ), .ip2(n9780), .s(n9946), .op(
        n2498) );
  mux2_1 U11256 ( .ip1(\ANSWER/mem[3][7][13] ), .ip2(n9780), .s(n9947), .op(
        n2497) );
  mux2_1 U11257 ( .ip1(\ANSWER/mem[3][8][13] ), .ip2(n9780), .s(n9948), .op(
        n2496) );
  mux2_1 U11258 ( .ip1(\ANSWER/mem[3][9][13] ), .ip2(n9780), .s(n9949), .op(
        n2495) );
  mux2_1 U11259 ( .ip1(\ANSWER/mem[4][0][13] ), .ip2(n9780), .s(n9950), .op(
        n2494) );
  mux2_1 U11260 ( .ip1(\ANSWER/mem[4][1][13] ), .ip2(n9780), .s(n9951), .op(
        n2493) );
  mux2_1 U11261 ( .ip1(\ANSWER/mem[4][2][13] ), .ip2(n9780), .s(n9952), .op(
        n2492) );
  mux2_1 U11262 ( .ip1(\ANSWER/mem[4][3][13] ), .ip2(n9781), .s(n9953), .op(
        n2491) );
  mux2_1 U11263 ( .ip1(\ANSWER/mem[4][4][13] ), .ip2(n9781), .s(n9954), .op(
        n2490) );
  mux2_1 U11264 ( .ip1(\ANSWER/mem[4][5][13] ), .ip2(n9781), .s(n9955), .op(
        n2489) );
  mux2_1 U11265 ( .ip1(\ANSWER/mem[4][6][13] ), .ip2(n9781), .s(n9956), .op(
        n2488) );
  mux2_1 U11266 ( .ip1(\ANSWER/mem[4][7][13] ), .ip2(n9781), .s(n9957), .op(
        n2487) );
  mux2_1 U11267 ( .ip1(\ANSWER/mem[4][8][13] ), .ip2(n9781), .s(n9958), .op(
        n2486) );
  mux2_1 U11268 ( .ip1(\ANSWER/mem[4][9][13] ), .ip2(n9781), .s(n9959), .op(
        n2485) );
  mux2_1 U11269 ( .ip1(\ANSWER/mem[5][0][13] ), .ip2(n9781), .s(n9960), .op(
        n2484) );
  mux2_1 U11270 ( .ip1(\ANSWER/mem[5][1][13] ), .ip2(n9781), .s(n9961), .op(
        n2483) );
  mux2_1 U11271 ( .ip1(\ANSWER/mem[5][2][13] ), .ip2(n9781), .s(n9962), .op(
        n2482) );
  mux2_1 U11272 ( .ip1(\ANSWER/mem[5][3][13] ), .ip2(n9780), .s(n9963), .op(
        n2481) );
  mux2_1 U11273 ( .ip1(\ANSWER/mem[5][4][13] ), .ip2(n9781), .s(n9964), .op(
        n2480) );
  mux2_1 U11274 ( .ip1(\ANSWER/mem[5][5][13] ), .ip2(n9780), .s(n9965), .op(
        n2479) );
  mux2_1 U11275 ( .ip1(\ANSWER/mem[5][6][13] ), .ip2(n9780), .s(n9966), .op(
        n2478) );
  mux2_1 U11276 ( .ip1(\ANSWER/mem[5][7][13] ), .ip2(n9780), .s(n9967), .op(
        n2477) );
  mux2_1 U11277 ( .ip1(\ANSWER/mem[5][8][13] ), .ip2(n9780), .s(n9968), .op(
        n2476) );
  mux2_1 U11278 ( .ip1(\ANSWER/mem[5][9][13] ), .ip2(n9780), .s(n9969), .op(
        n2475) );
  mux2_1 U11279 ( .ip1(\ANSWER/mem[6][0][13] ), .ip2(n9780), .s(n9970), .op(
        n2474) );
  mux2_1 U11280 ( .ip1(\ANSWER/mem[6][1][13] ), .ip2(n9780), .s(n9971), .op(
        n2473) );
  mux2_1 U11281 ( .ip1(\ANSWER/mem[6][2][13] ), .ip2(n9780), .s(n9972), .op(
        n2472) );
  mux2_1 U11282 ( .ip1(\ANSWER/mem[6][3][13] ), .ip2(n9780), .s(n9973), .op(
        n2471) );
  mux2_1 U11283 ( .ip1(\ANSWER/mem[6][4][13] ), .ip2(n9780), .s(n9974), .op(
        n2470) );
  mux2_1 U11284 ( .ip1(\ANSWER/mem[6][5][13] ), .ip2(n9780), .s(n9975), .op(
        n2469) );
  mux2_1 U11285 ( .ip1(\ANSWER/mem[6][6][13] ), .ip2(n9780), .s(n9976), .op(
        n2468) );
  mux2_1 U11286 ( .ip1(\ANSWER/mem[6][7][13] ), .ip2(n9780), .s(n9977), .op(
        n2467) );
  mux2_1 U11287 ( .ip1(\ANSWER/mem[6][8][13] ), .ip2(n9780), .s(n9978), .op(
        n2466) );
  mux2_1 U11288 ( .ip1(\ANSWER/mem[6][9][13] ), .ip2(n9780), .s(n9979), .op(
        n2465) );
  mux2_1 U11289 ( .ip1(\ANSWER/mem[7][0][13] ), .ip2(n9780), .s(n9980), .op(
        n2464) );
  mux2_1 U11290 ( .ip1(\ANSWER/mem[7][1][13] ), .ip2(n9780), .s(n9981), .op(
        n2463) );
  buf_1 U11291 ( .ip(n9780), .op(n9781) );
  mux2_1 U11292 ( .ip1(\ANSWER/mem[7][2][13] ), .ip2(n9781), .s(n9983), .op(
        n2462) );
  mux2_1 U11293 ( .ip1(\ANSWER/mem[7][3][13] ), .ip2(n9781), .s(n9984), .op(
        n2461) );
  mux2_1 U11294 ( .ip1(\ANSWER/mem[7][4][13] ), .ip2(n9781), .s(n9985), .op(
        n2460) );
  mux2_1 U11295 ( .ip1(\ANSWER/mem[7][5][13] ), .ip2(n9781), .s(n9986), .op(
        n2459) );
  mux2_1 U11296 ( .ip1(\ANSWER/mem[7][6][13] ), .ip2(n9781), .s(n9987), .op(
        n2458) );
  mux2_1 U11297 ( .ip1(\ANSWER/mem[7][7][13] ), .ip2(n9781), .s(n9988), .op(
        n2457) );
  mux2_1 U11298 ( .ip1(\ANSWER/mem[7][8][13] ), .ip2(n9781), .s(n9989), .op(
        n2456) );
  mux2_1 U11299 ( .ip1(\ANSWER/mem[7][9][13] ), .ip2(n9781), .s(n9990), .op(
        n2455) );
  mux2_1 U11300 ( .ip1(\ANSWER/mem[8][0][13] ), .ip2(n9780), .s(n9991), .op(
        n2454) );
  mux2_1 U11301 ( .ip1(\ANSWER/mem[8][1][13] ), .ip2(n9781), .s(n9992), .op(
        n2453) );
  mux2_1 U11302 ( .ip1(\ANSWER/mem[8][2][13] ), .ip2(n9781), .s(n9993), .op(
        n2452) );
  mux2_1 U11303 ( .ip1(\ANSWER/mem[8][3][13] ), .ip2(n9781), .s(n9994), .op(
        n2451) );
  mux2_1 U11304 ( .ip1(\ANSWER/mem[8][4][13] ), .ip2(n9780), .s(n9996), .op(
        n2450) );
  mux2_1 U11305 ( .ip1(\ANSWER/mem[8][5][13] ), .ip2(n9780), .s(n9997), .op(
        n2449) );
  mux2_1 U11306 ( .ip1(\ANSWER/mem[8][6][13] ), .ip2(n9780), .s(n9998), .op(
        n2448) );
  mux2_1 U11307 ( .ip1(\ANSWER/mem[8][7][13] ), .ip2(n9780), .s(n9999), .op(
        n2447) );
  mux2_1 U11308 ( .ip1(\ANSWER/mem[8][8][13] ), .ip2(n9780), .s(n10000), .op(
        n2446) );
  mux2_1 U11309 ( .ip1(\ANSWER/mem[8][9][13] ), .ip2(n9780), .s(n10001), .op(
        n2445) );
  mux2_1 U11310 ( .ip1(\ANSWER/mem[9][0][13] ), .ip2(n9780), .s(n10002), .op(
        n2444) );
  mux2_1 U11311 ( .ip1(\ANSWER/mem[9][1][13] ), .ip2(n9780), .s(n10003), .op(
        n2443) );
  mux2_1 U11312 ( .ip1(\ANSWER/mem[9][2][13] ), .ip2(n9780), .s(n10004), .op(
        n2442) );
  mux2_1 U11313 ( .ip1(\ANSWER/mem[9][3][13] ), .ip2(n9780), .s(n10005), .op(
        n2441) );
  mux2_1 U11314 ( .ip1(\ANSWER/mem[9][4][13] ), .ip2(n9780), .s(n10006), .op(
        n2440) );
  mux2_1 U11315 ( .ip1(\ANSWER/mem[9][5][13] ), .ip2(n9780), .s(n10007), .op(
        n2439) );
  mux2_1 U11316 ( .ip1(\ANSWER/mem[9][6][13] ), .ip2(n9781), .s(n10008), .op(
        n2438) );
  mux2_1 U11317 ( .ip1(\ANSWER/mem[9][7][13] ), .ip2(n9781), .s(n10009), .op(
        n2437) );
  mux2_1 U11318 ( .ip1(\ANSWER/mem[9][8][13] ), .ip2(n9781), .s(n10010), .op(
        n2436) );
  mux2_1 U11319 ( .ip1(\ANSWER/mem[9][9][13] ), .ip2(n9781), .s(n10011), .op(
        n2435) );
  fulladder U11320 ( .a(n9784), .b(n9783), .ci(n9782), .co(n9871), .s(n9833)
         );
  fulladder U11321 ( .a(n9787), .b(n9786), .ci(n9785), .co(n9841), .s(n9727)
         );
  nor2_1 U11322 ( .ip1(n9863), .ip2(n9788), .op(n9844) );
  nor2_1 U11323 ( .ip1(n9790), .ip2(n9789), .op(n9843) );
  nand2_1 U11324 ( .ip1(m2DataIn[7]), .ip2(q_w2[15]), .op(n9842) );
  nor3_1 U11325 ( .ip1(n9792), .ip2(n9791), .ip3(n9898), .op(n9796) );
  or2_1 U11326 ( .ip1(q_w2[12]), .ip2(n9793), .op(n9795) );
  or2_1 U11327 ( .ip1(m2DataIn[10]), .ip2(n9793), .op(n9794) );
  nand2_1 U11328 ( .ip1(n9795), .ip2(n9794), .op(n9896) );
  nor2_1 U11329 ( .ip1(n9796), .ip2(n9896), .op(n9797) );
  mux2_1 U11330 ( .ip1(rdata[14]), .ip2(n9895), .s(n9797), .op(n9839) );
  inv_1 U11331 ( .ip(n9798), .op(n9852) );
  nor2_1 U11332 ( .ip1(n9799), .ip2(n9864), .op(n9889) );
  nand2_1 U11333 ( .ip1(rdata[13]), .ip2(n9800), .op(n9801) );
  nand2_1 U11334 ( .ip1(n9802), .ip2(n9801), .op(n9888) );
  fulladder U11335 ( .a(n9805), .b(n9804), .ci(n9803), .co(n9887), .s(n9726)
         );
  inv_1 U11336 ( .ip(n9806), .op(n9851) );
  fulladder U11337 ( .a(n9809), .b(n9808), .ci(n9807), .co(n9850), .s(n9831)
         );
  and3_1 U11338 ( .ip1(m2DataIn[13]), .ip2(q_w2[7]), .ip3(n9844), .op(n9813)
         );
  nor2_1 U11339 ( .ip1(n9811), .ip2(n9810), .op(n9812) );
  nor2_1 U11340 ( .ip1(n9813), .ip2(n9812), .op(n9882) );
  nor2_1 U11341 ( .ip1(n9815), .ip2(n9814), .op(n9879) );
  nor2_1 U11342 ( .ip1(n9817), .ip2(n9816), .op(n9878) );
  nand2_1 U11343 ( .ip1(m2DataIn[15]), .ip2(q_w2[7]), .op(n9877) );
  inv_1 U11344 ( .ip(n9818), .op(n9881) );
  fulladder U11345 ( .a(n9821), .b(n9820), .ci(n9819), .co(n9880), .s(n9830)
         );
  fulladder U11346 ( .a(n9824), .b(n9823), .ci(n9822), .co(n9847), .s(n9764)
         );
  fulladder U11347 ( .a(n9827), .b(n9826), .ci(n9825), .co(n9828), .s(n9768)
         );
  inv_1 U11348 ( .ip(n9828), .op(n9873) );
  fulladder U11349 ( .a(n9831), .b(n9830), .ci(n9829), .co(n9872), .s(n9749)
         );
  fulladder U11350 ( .a(n9834), .b(n9833), .ci(n9832), .co(n9869), .s(n9778)
         );
  nor2_1 U11351 ( .ip1(n9907), .ip2(n9835), .op(n9837) );
  buf_1 U11352 ( .ip(n9837), .op(n9836) );
  mux2_1 U11353 ( .ip1(\ANSWER/mem[0][0][14] ), .ip2(n9836), .s(n9910), .op(
        n2434) );
  mux2_1 U11354 ( .ip1(\ANSWER/mem[0][1][14] ), .ip2(n9836), .s(n9911), .op(
        n2433) );
  mux2_1 U11355 ( .ip1(\ANSWER/mem[0][2][14] ), .ip2(n9836), .s(n9912), .op(
        n2432) );
  mux2_1 U11356 ( .ip1(\ANSWER/mem[0][3][14] ), .ip2(n9836), .s(n9913), .op(
        n2431) );
  mux2_1 U11357 ( .ip1(\ANSWER/mem[0][4][14] ), .ip2(n9836), .s(n9914), .op(
        n2430) );
  mux2_1 U11358 ( .ip1(\ANSWER/mem[0][5][14] ), .ip2(n9836), .s(n9915), .op(
        n2429) );
  mux2_1 U11359 ( .ip1(\ANSWER/mem[0][6][14] ), .ip2(n9836), .s(n9916), .op(
        n2428) );
  mux2_1 U11360 ( .ip1(\ANSWER/mem[0][7][14] ), .ip2(n9836), .s(n9917), .op(
        n2427) );
  mux2_1 U11361 ( .ip1(\ANSWER/mem[0][8][14] ), .ip2(n9836), .s(n9918), .op(
        n2426) );
  mux2_1 U11362 ( .ip1(\ANSWER/mem[0][9][14] ), .ip2(n9836), .s(n9919), .op(
        n2425) );
  mux2_1 U11363 ( .ip1(\ANSWER/mem[1][0][14] ), .ip2(n9836), .s(n9920), .op(
        n2424) );
  mux2_1 U11364 ( .ip1(\ANSWER/mem[1][1][14] ), .ip2(n9836), .s(n9921), .op(
        n2423) );
  mux2_1 U11365 ( .ip1(\ANSWER/mem[1][2][14] ), .ip2(n9836), .s(n9922), .op(
        n2422) );
  mux2_1 U11366 ( .ip1(\ANSWER/mem[1][3][14] ), .ip2(n9836), .s(n9923), .op(
        n2421) );
  mux2_1 U11367 ( .ip1(\ANSWER/mem[1][4][14] ), .ip2(n9836), .s(n9924), .op(
        n2420) );
  mux2_1 U11368 ( .ip1(\ANSWER/mem[1][5][14] ), .ip2(n9836), .s(n9925), .op(
        n2419) );
  mux2_1 U11369 ( .ip1(\ANSWER/mem[1][6][14] ), .ip2(n9836), .s(n9926), .op(
        n2418) );
  mux2_1 U11370 ( .ip1(\ANSWER/mem[1][7][14] ), .ip2(n9836), .s(n9927), .op(
        n2417) );
  mux2_1 U11371 ( .ip1(\ANSWER/mem[1][8][14] ), .ip2(n9836), .s(n9928), .op(
        n2416) );
  mux2_1 U11372 ( .ip1(\ANSWER/mem[1][9][14] ), .ip2(n9836), .s(n9929), .op(
        n2415) );
  mux2_1 U11373 ( .ip1(\ANSWER/mem[2][0][14] ), .ip2(n9836), .s(n9930), .op(
        n2414) );
  mux2_1 U11374 ( .ip1(\ANSWER/mem[2][1][14] ), .ip2(n9836), .s(n9931), .op(
        n2413) );
  mux2_1 U11375 ( .ip1(\ANSWER/mem[2][2][14] ), .ip2(n9836), .s(n9932), .op(
        n2412) );
  mux2_1 U11376 ( .ip1(\ANSWER/mem[2][3][14] ), .ip2(n9836), .s(n9933), .op(
        n2411) );
  mux2_1 U11377 ( .ip1(\ANSWER/mem[2][4][14] ), .ip2(n9836), .s(n9934), .op(
        n2410) );
  mux2_1 U11378 ( .ip1(\ANSWER/mem[2][5][14] ), .ip2(n9836), .s(n9935), .op(
        n2409) );
  mux2_1 U11379 ( .ip1(\ANSWER/mem[2][6][14] ), .ip2(n9836), .s(n9936), .op(
        n2408) );
  mux2_1 U11380 ( .ip1(\ANSWER/mem[2][7][14] ), .ip2(n9836), .s(n9937), .op(
        n2407) );
  mux2_1 U11381 ( .ip1(\ANSWER/mem[2][8][14] ), .ip2(n9836), .s(n9938), .op(
        n2406) );
  mux2_1 U11382 ( .ip1(\ANSWER/mem[2][9][14] ), .ip2(n9836), .s(n9939), .op(
        n2405) );
  mux2_1 U11383 ( .ip1(\ANSWER/mem[3][0][14] ), .ip2(n9836), .s(n9940), .op(
        n2404) );
  mux2_1 U11384 ( .ip1(\ANSWER/mem[3][1][14] ), .ip2(n9836), .s(n9941), .op(
        n2403) );
  mux2_1 U11385 ( .ip1(\ANSWER/mem[3][2][14] ), .ip2(n9836), .s(n9942), .op(
        n2402) );
  mux2_1 U11386 ( .ip1(\ANSWER/mem[3][3][14] ), .ip2(n9836), .s(n9943), .op(
        n2401) );
  mux2_1 U11387 ( .ip1(\ANSWER/mem[3][4][14] ), .ip2(n9836), .s(n9944), .op(
        n2400) );
  mux2_1 U11388 ( .ip1(\ANSWER/mem[3][5][14] ), .ip2(n9836), .s(n9945), .op(
        n2399) );
  mux2_1 U11389 ( .ip1(\ANSWER/mem[3][6][14] ), .ip2(n9837), .s(n9946), .op(
        n2398) );
  mux2_1 U11390 ( .ip1(\ANSWER/mem[3][7][14] ), .ip2(n9837), .s(n9947), .op(
        n2397) );
  mux2_1 U11391 ( .ip1(\ANSWER/mem[3][8][14] ), .ip2(n9837), .s(n9948), .op(
        n2396) );
  mux2_1 U11392 ( .ip1(\ANSWER/mem[3][9][14] ), .ip2(n9837), .s(n9949), .op(
        n2395) );
  mux2_1 U11393 ( .ip1(\ANSWER/mem[4][0][14] ), .ip2(n9837), .s(n9950), .op(
        n2394) );
  mux2_1 U11394 ( .ip1(\ANSWER/mem[4][1][14] ), .ip2(n9837), .s(n9951), .op(
        n2393) );
  mux2_1 U11395 ( .ip1(\ANSWER/mem[4][2][14] ), .ip2(n9837), .s(n9952), .op(
        n2392) );
  mux2_1 U11396 ( .ip1(\ANSWER/mem[4][3][14] ), .ip2(n9838), .s(n9953), .op(
        n2391) );
  mux2_1 U11397 ( .ip1(\ANSWER/mem[4][4][14] ), .ip2(n9838), .s(n9954), .op(
        n2390) );
  mux2_1 U11398 ( .ip1(\ANSWER/mem[4][5][14] ), .ip2(n9838), .s(n9955), .op(
        n2389) );
  mux2_1 U11399 ( .ip1(\ANSWER/mem[4][6][14] ), .ip2(n9838), .s(n9956), .op(
        n2388) );
  mux2_1 U11400 ( .ip1(\ANSWER/mem[4][7][14] ), .ip2(n9838), .s(n9957), .op(
        n2387) );
  mux2_1 U11401 ( .ip1(\ANSWER/mem[4][8][14] ), .ip2(n9838), .s(n9958), .op(
        n2386) );
  mux2_1 U11402 ( .ip1(\ANSWER/mem[4][9][14] ), .ip2(n9838), .s(n9959), .op(
        n2385) );
  mux2_1 U11403 ( .ip1(\ANSWER/mem[5][0][14] ), .ip2(n9838), .s(n9960), .op(
        n2384) );
  mux2_1 U11404 ( .ip1(\ANSWER/mem[5][1][14] ), .ip2(n9838), .s(n9961), .op(
        n2383) );
  mux2_1 U11405 ( .ip1(\ANSWER/mem[5][2][14] ), .ip2(n9838), .s(n9962), .op(
        n2382) );
  mux2_1 U11406 ( .ip1(\ANSWER/mem[5][3][14] ), .ip2(n9837), .s(n9963), .op(
        n2381) );
  mux2_1 U11407 ( .ip1(\ANSWER/mem[5][4][14] ), .ip2(n9838), .s(n9964), .op(
        n2380) );
  mux2_1 U11408 ( .ip1(\ANSWER/mem[5][5][14] ), .ip2(n9837), .s(n9965), .op(
        n2379) );
  mux2_1 U11409 ( .ip1(\ANSWER/mem[5][6][14] ), .ip2(n9837), .s(n9966), .op(
        n2378) );
  mux2_1 U11410 ( .ip1(\ANSWER/mem[5][7][14] ), .ip2(n9837), .s(n9967), .op(
        n2377) );
  mux2_1 U11411 ( .ip1(\ANSWER/mem[5][8][14] ), .ip2(n9837), .s(n9968), .op(
        n2376) );
  mux2_1 U11412 ( .ip1(\ANSWER/mem[5][9][14] ), .ip2(n9837), .s(n9969), .op(
        n2375) );
  mux2_1 U11413 ( .ip1(\ANSWER/mem[6][0][14] ), .ip2(n9837), .s(n9970), .op(
        n2374) );
  mux2_1 U11414 ( .ip1(\ANSWER/mem[6][1][14] ), .ip2(n9837), .s(n9971), .op(
        n2373) );
  mux2_1 U11415 ( .ip1(\ANSWER/mem[6][2][14] ), .ip2(n9837), .s(n9972), .op(
        n2372) );
  mux2_1 U11416 ( .ip1(\ANSWER/mem[6][3][14] ), .ip2(n9837), .s(n9973), .op(
        n2371) );
  mux2_1 U11417 ( .ip1(\ANSWER/mem[6][4][14] ), .ip2(n9837), .s(n9974), .op(
        n2370) );
  mux2_1 U11418 ( .ip1(\ANSWER/mem[6][5][14] ), .ip2(n9837), .s(n9975), .op(
        n2369) );
  mux2_1 U11419 ( .ip1(\ANSWER/mem[6][6][14] ), .ip2(n9837), .s(n9976), .op(
        n2368) );
  mux2_1 U11420 ( .ip1(\ANSWER/mem[6][7][14] ), .ip2(n9837), .s(n9977), .op(
        n2367) );
  mux2_1 U11421 ( .ip1(\ANSWER/mem[6][8][14] ), .ip2(n9837), .s(n9978), .op(
        n2366) );
  mux2_1 U11422 ( .ip1(\ANSWER/mem[6][9][14] ), .ip2(n9837), .s(n9979), .op(
        n2365) );
  mux2_1 U11423 ( .ip1(\ANSWER/mem[7][0][14] ), .ip2(n9837), .s(n9980), .op(
        n2364) );
  mux2_1 U11424 ( .ip1(\ANSWER/mem[7][1][14] ), .ip2(n9837), .s(n9981), .op(
        n2363) );
  buf_1 U11425 ( .ip(n9837), .op(n9838) );
  mux2_1 U11426 ( .ip1(\ANSWER/mem[7][2][14] ), .ip2(n9838), .s(n9983), .op(
        n2362) );
  mux2_1 U11427 ( .ip1(\ANSWER/mem[7][3][14] ), .ip2(n9838), .s(n9984), .op(
        n2361) );
  mux2_1 U11428 ( .ip1(\ANSWER/mem[7][4][14] ), .ip2(n9838), .s(n9985), .op(
        n2360) );
  mux2_1 U11429 ( .ip1(\ANSWER/mem[7][5][14] ), .ip2(n9838), .s(n9986), .op(
        n2359) );
  mux2_1 U11430 ( .ip1(\ANSWER/mem[7][6][14] ), .ip2(n9838), .s(n9987), .op(
        n2358) );
  mux2_1 U11431 ( .ip1(\ANSWER/mem[7][7][14] ), .ip2(n9838), .s(n9988), .op(
        n2357) );
  mux2_1 U11432 ( .ip1(\ANSWER/mem[7][8][14] ), .ip2(n9838), .s(n9989), .op(
        n2356) );
  mux2_1 U11433 ( .ip1(\ANSWER/mem[7][9][14] ), .ip2(n9838), .s(n9990), .op(
        n2355) );
  mux2_1 U11434 ( .ip1(\ANSWER/mem[8][0][14] ), .ip2(n9837), .s(n9991), .op(
        n2354) );
  mux2_1 U11435 ( .ip1(\ANSWER/mem[8][1][14] ), .ip2(n9838), .s(n9992), .op(
        n2353) );
  mux2_1 U11436 ( .ip1(\ANSWER/mem[8][2][14] ), .ip2(n9838), .s(n9993), .op(
        n2352) );
  mux2_1 U11437 ( .ip1(\ANSWER/mem[8][3][14] ), .ip2(n9838), .s(n9994), .op(
        n2351) );
  mux2_1 U11438 ( .ip1(\ANSWER/mem[8][4][14] ), .ip2(n9837), .s(n9996), .op(
        n2350) );
  mux2_1 U11439 ( .ip1(\ANSWER/mem[8][5][14] ), .ip2(n9837), .s(n9997), .op(
        n2349) );
  mux2_1 U11440 ( .ip1(\ANSWER/mem[8][6][14] ), .ip2(n9837), .s(n9998), .op(
        n2348) );
  mux2_1 U11441 ( .ip1(\ANSWER/mem[8][7][14] ), .ip2(n9837), .s(n9999), .op(
        n2347) );
  mux2_1 U11442 ( .ip1(\ANSWER/mem[8][8][14] ), .ip2(n9837), .s(n10000), .op(
        n2346) );
  mux2_1 U11443 ( .ip1(\ANSWER/mem[8][9][14] ), .ip2(n9837), .s(n10001), .op(
        n2345) );
  mux2_1 U11444 ( .ip1(\ANSWER/mem[9][0][14] ), .ip2(n9837), .s(n10002), .op(
        n2344) );
  mux2_1 U11445 ( .ip1(\ANSWER/mem[9][1][14] ), .ip2(n9837), .s(n10003), .op(
        n2343) );
  mux2_1 U11446 ( .ip1(\ANSWER/mem[9][2][14] ), .ip2(n9837), .s(n10004), .op(
        n2342) );
  mux2_1 U11447 ( .ip1(\ANSWER/mem[9][3][14] ), .ip2(n9837), .s(n10005), .op(
        n2341) );
  mux2_1 U11448 ( .ip1(\ANSWER/mem[9][4][14] ), .ip2(n9837), .s(n10006), .op(
        n2340) );
  mux2_1 U11449 ( .ip1(\ANSWER/mem[9][5][14] ), .ip2(n9837), .s(n10007), .op(
        n2339) );
  mux2_1 U11450 ( .ip1(\ANSWER/mem[9][6][14] ), .ip2(n9838), .s(n10008), .op(
        n2338) );
  mux2_1 U11451 ( .ip1(\ANSWER/mem[9][7][14] ), .ip2(n9838), .s(n10009), .op(
        n2337) );
  mux2_1 U11452 ( .ip1(\ANSWER/mem[9][8][14] ), .ip2(n9838), .s(n10010), .op(
        n2336) );
  mux2_1 U11453 ( .ip1(\ANSWER/mem[9][9][14] ), .ip2(n9838), .s(n10011), .op(
        n2335) );
  fulladder U11454 ( .a(n9841), .b(n9840), .ci(n9839), .co(n9846), .s(n9798)
         );
  fulladder U11455 ( .a(n9844), .b(n9843), .ci(n9842), .co(n9845), .s(n9840)
         );
  xor2_1 U11456 ( .ip1(n9846), .ip2(n9845), .op(n9856) );
  fulladder U11457 ( .a(n9849), .b(n9848), .ci(n9847), .co(n9854), .s(n9874)
         );
  fulladder U11458 ( .a(n9852), .b(n9851), .ci(n9850), .co(n9853), .s(n9849)
         );
  xor2_1 U11459 ( .ip1(n9854), .ip2(n9853), .op(n9855) );
  xor2_1 U11460 ( .ip1(n9856), .ip2(n9855), .op(n9860) );
  nand2_1 U11461 ( .ip1(q_w2[15]), .ip2(m2DataIn[8]), .op(n9858) );
  nand2_1 U11462 ( .ip1(q_w2[8]), .ip2(m2DataIn[15]), .op(n9857) );
  xor2_1 U11463 ( .ip1(n9858), .ip2(n9857), .op(n9859) );
  xor2_1 U11464 ( .ip1(n9860), .ip2(n9859), .op(n9861) );
  xor2_1 U11465 ( .ip1(n9862), .ip2(n9861), .op(n9909) );
  nor2_1 U11466 ( .ip1(n9864), .ip2(n9863), .op(n9866) );
  nand2_1 U11467 ( .ip1(q_w2[11]), .ip2(m2DataIn[12]), .op(n9865) );
  xor2_1 U11468 ( .ip1(n9866), .ip2(n9865), .op(n9905) );
  nand2_1 U11469 ( .ip1(q_w2[10]), .ip2(m2DataIn[13]), .op(n9868) );
  nand2_1 U11470 ( .ip1(q_w2[13]), .ip2(m2DataIn[10]), .op(n9867) );
  xor2_1 U11471 ( .ip1(n9868), .ip2(n9867), .op(n9903) );
  fulladder U11472 ( .a(n9871), .b(n9870), .ci(n9869), .co(n9876), .s(n9835)
         );
  fulladder U11473 ( .a(n9874), .b(n9873), .ci(n9872), .co(n9875), .s(n9870)
         );
  xor2_1 U11474 ( .ip1(n9876), .ip2(n9875), .op(n9886) );
  fulladder U11475 ( .a(n9879), .b(n9878), .ci(n9877), .co(n9884), .s(n9818)
         );
  fulladder U11476 ( .a(n9882), .b(n9881), .ci(n9880), .co(n9883), .s(n9848)
         );
  xor2_1 U11477 ( .ip1(n9884), .ip2(n9883), .op(n9885) );
  xor2_1 U11478 ( .ip1(n9886), .ip2(n9885), .op(n9893) );
  inv_1 U11479 ( .ip(rdata[15]), .op(n9891) );
  fulladder U11480 ( .a(n9889), .b(n9888), .ci(n9887), .co(n9890), .s(n9806)
         );
  mux2_1 U11481 ( .ip1(n9891), .ip2(rdata[15]), .s(n9890), .op(n9892) );
  xor2_1 U11482 ( .ip1(n9893), .ip2(n9892), .op(n9901) );
  nor2_1 U11483 ( .ip1(n9894), .ip2(n9898), .op(n9899) );
  nor2_1 U11484 ( .ip1(n9896), .ip2(n9895), .op(n9897) );
  mux2_1 U11485 ( .ip1(n9899), .ip2(n9898), .s(n9897), .op(n9900) );
  xor2_1 U11486 ( .ip1(n9901), .ip2(n9900), .op(n9902) );
  xor2_1 U11487 ( .ip1(n9903), .ip2(n9902), .op(n9904) );
  xor2_1 U11488 ( .ip1(n9905), .ip2(n9904), .op(n9908) );
  nor2_1 U11489 ( .ip1(n9909), .ip2(n9908), .op(n9906) );
  not_ab_or_c_or_d U11490 ( .ip1(n9909), .ip2(n9908), .ip3(n9907), .ip4(n9906), 
        .op(n9982) );
  buf_1 U11491 ( .ip(n9982), .op(n10012) );
  mux2_1 U11492 ( .ip1(\ANSWER/mem[0][0][15] ), .ip2(n10012), .s(n9910), .op(
        n2334) );
  mux2_1 U11493 ( .ip1(\ANSWER/mem[0][1][15] ), .ip2(n10012), .s(n9911), .op(
        n2333) );
  mux2_1 U11494 ( .ip1(\ANSWER/mem[0][2][15] ), .ip2(n10012), .s(n9912), .op(
        n2332) );
  mux2_1 U11495 ( .ip1(\ANSWER/mem[0][3][15] ), .ip2(n10012), .s(n9913), .op(
        n2331) );
  mux2_1 U11496 ( .ip1(\ANSWER/mem[0][4][15] ), .ip2(n10012), .s(n9914), .op(
        n2330) );
  mux2_1 U11497 ( .ip1(\ANSWER/mem[0][5][15] ), .ip2(n10012), .s(n9915), .op(
        n2329) );
  mux2_1 U11498 ( .ip1(\ANSWER/mem[0][6][15] ), .ip2(n10012), .s(n9916), .op(
        n2328) );
  mux2_1 U11499 ( .ip1(\ANSWER/mem[0][7][15] ), .ip2(n10012), .s(n9917), .op(
        n2327) );
  mux2_1 U11500 ( .ip1(\ANSWER/mem[0][8][15] ), .ip2(n10012), .s(n9918), .op(
        n2326) );
  mux2_1 U11501 ( .ip1(\ANSWER/mem[0][9][15] ), .ip2(n10012), .s(n9919), .op(
        n2325) );
  mux2_1 U11502 ( .ip1(\ANSWER/mem[1][0][15] ), .ip2(n10012), .s(n9920), .op(
        n2324) );
  mux2_1 U11503 ( .ip1(\ANSWER/mem[1][1][15] ), .ip2(n10012), .s(n9921), .op(
        n2323) );
  mux2_1 U11504 ( .ip1(\ANSWER/mem[1][2][15] ), .ip2(n10012), .s(n9922), .op(
        n2322) );
  mux2_1 U11505 ( .ip1(\ANSWER/mem[1][3][15] ), .ip2(n10012), .s(n9923), .op(
        n2321) );
  mux2_1 U11506 ( .ip1(\ANSWER/mem[1][4][15] ), .ip2(n10012), .s(n9924), .op(
        n2320) );
  mux2_1 U11507 ( .ip1(\ANSWER/mem[1][5][15] ), .ip2(n10012), .s(n9925), .op(
        n2319) );
  mux2_1 U11508 ( .ip1(\ANSWER/mem[1][6][15] ), .ip2(n9982), .s(n9926), .op(
        n2318) );
  mux2_1 U11509 ( .ip1(\ANSWER/mem[1][7][15] ), .ip2(n9982), .s(n9927), .op(
        n2317) );
  mux2_1 U11510 ( .ip1(\ANSWER/mem[1][8][15] ), .ip2(n10012), .s(n9928), .op(
        n2316) );
  mux2_1 U11511 ( .ip1(\ANSWER/mem[1][9][15] ), .ip2(n10012), .s(n9929), .op(
        n2315) );
  mux2_1 U11512 ( .ip1(\ANSWER/mem[2][0][15] ), .ip2(n10012), .s(n9930), .op(
        n2314) );
  mux2_1 U11513 ( .ip1(\ANSWER/mem[2][1][15] ), .ip2(n10012), .s(n9931), .op(
        n2313) );
  mux2_1 U11514 ( .ip1(\ANSWER/mem[2][2][15] ), .ip2(n10012), .s(n9932), .op(
        n2312) );
  mux2_1 U11515 ( .ip1(\ANSWER/mem[2][3][15] ), .ip2(n9982), .s(n9933), .op(
        n2311) );
  mux2_1 U11516 ( .ip1(\ANSWER/mem[2][4][15] ), .ip2(n9982), .s(n9934), .op(
        n2310) );
  mux2_1 U11517 ( .ip1(\ANSWER/mem[2][5][15] ), .ip2(n9982), .s(n9935), .op(
        n2309) );
  mux2_1 U11518 ( .ip1(\ANSWER/mem[2][6][15] ), .ip2(n9982), .s(n9936), .op(
        n2308) );
  mux2_1 U11519 ( .ip1(\ANSWER/mem[2][7][15] ), .ip2(n9982), .s(n9937), .op(
        n2307) );
  mux2_1 U11520 ( .ip1(\ANSWER/mem[2][8][15] ), .ip2(n9982), .s(n9938), .op(
        n2306) );
  mux2_1 U11521 ( .ip1(\ANSWER/mem[2][9][15] ), .ip2(n9982), .s(n9939), .op(
        n2305) );
  mux2_1 U11522 ( .ip1(\ANSWER/mem[3][0][15] ), .ip2(n9982), .s(n9940), .op(
        n2304) );
  mux2_1 U11523 ( .ip1(\ANSWER/mem[3][1][15] ), .ip2(n9982), .s(n9941), .op(
        n2303) );
  mux2_1 U11524 ( .ip1(\ANSWER/mem[3][2][15] ), .ip2(n9982), .s(n9942), .op(
        n2302) );
  mux2_1 U11525 ( .ip1(\ANSWER/mem[3][3][15] ), .ip2(n9982), .s(n9943), .op(
        n2301) );
  mux2_1 U11526 ( .ip1(\ANSWER/mem[3][4][15] ), .ip2(n9982), .s(n9944), .op(
        n2300) );
  mux2_1 U11527 ( .ip1(\ANSWER/mem[3][5][15] ), .ip2(n9982), .s(n9945), .op(
        n2299) );
  buf_1 U11528 ( .ip(n9982), .op(n9995) );
  mux2_1 U11529 ( .ip1(\ANSWER/mem[3][6][15] ), .ip2(n9995), .s(n9946), .op(
        n2298) );
  mux2_1 U11530 ( .ip1(\ANSWER/mem[3][7][15] ), .ip2(n9982), .s(n9947), .op(
        n2297) );
  mux2_1 U11531 ( .ip1(\ANSWER/mem[3][8][15] ), .ip2(n9995), .s(n9948), .op(
        n2296) );
  mux2_1 U11532 ( .ip1(\ANSWER/mem[3][9][15] ), .ip2(n9995), .s(n9949), .op(
        n2295) );
  mux2_1 U11533 ( .ip1(\ANSWER/mem[4][0][15] ), .ip2(n9995), .s(n9950), .op(
        n2294) );
  mux2_1 U11534 ( .ip1(\ANSWER/mem[4][1][15] ), .ip2(n9995), .s(n9951), .op(
        n2293) );
  mux2_1 U11535 ( .ip1(\ANSWER/mem[4][2][15] ), .ip2(n9995), .s(n9952), .op(
        n2292) );
  mux2_1 U11536 ( .ip1(\ANSWER/mem[4][3][15] ), .ip2(n9982), .s(n9953), .op(
        n2291) );
  mux2_1 U11537 ( .ip1(\ANSWER/mem[4][4][15] ), .ip2(n9982), .s(n9954), .op(
        n2290) );
  mux2_1 U11538 ( .ip1(\ANSWER/mem[4][5][15] ), .ip2(n9982), .s(n9955), .op(
        n2289) );
  mux2_1 U11539 ( .ip1(\ANSWER/mem[4][6][15] ), .ip2(n9995), .s(n9956), .op(
        n2288) );
  mux2_1 U11540 ( .ip1(\ANSWER/mem[4][7][15] ), .ip2(n9995), .s(n9957), .op(
        n2287) );
  mux2_1 U11541 ( .ip1(\ANSWER/mem[4][8][15] ), .ip2(n9982), .s(n9958), .op(
        n2286) );
  mux2_1 U11542 ( .ip1(\ANSWER/mem[4][9][15] ), .ip2(n9982), .s(n9959), .op(
        n2285) );
  mux2_1 U11543 ( .ip1(\ANSWER/mem[5][0][15] ), .ip2(n9982), .s(n9960), .op(
        n2284) );
  mux2_1 U11544 ( .ip1(\ANSWER/mem[5][1][15] ), .ip2(n9982), .s(n9961), .op(
        n2283) );
  mux2_1 U11545 ( .ip1(\ANSWER/mem[5][2][15] ), .ip2(n9982), .s(n9962), .op(
        n2282) );
  mux2_1 U11546 ( .ip1(\ANSWER/mem[5][3][15] ), .ip2(n9995), .s(n9963), .op(
        n2281) );
  mux2_1 U11547 ( .ip1(\ANSWER/mem[5][4][15] ), .ip2(n9982), .s(n9964), .op(
        n2280) );
  mux2_1 U11548 ( .ip1(\ANSWER/mem[5][5][15] ), .ip2(n9982), .s(n9965), .op(
        n2279) );
  mux2_1 U11549 ( .ip1(\ANSWER/mem[5][6][15] ), .ip2(n9982), .s(n9966), .op(
        n2278) );
  mux2_1 U11550 ( .ip1(\ANSWER/mem[5][7][15] ), .ip2(n9982), .s(n9967), .op(
        n2277) );
  mux2_1 U11551 ( .ip1(\ANSWER/mem[5][8][15] ), .ip2(n9982), .s(n9968), .op(
        n2276) );
  mux2_1 U11552 ( .ip1(\ANSWER/mem[5][9][15] ), .ip2(n9982), .s(n9969), .op(
        n2275) );
  mux2_1 U11553 ( .ip1(\ANSWER/mem[6][0][15] ), .ip2(n9982), .s(n9970), .op(
        n2274) );
  mux2_1 U11554 ( .ip1(\ANSWER/mem[6][1][15] ), .ip2(n9982), .s(n9971), .op(
        n2273) );
  mux2_1 U11555 ( .ip1(\ANSWER/mem[6][2][15] ), .ip2(n9982), .s(n9972), .op(
        n2272) );
  mux2_1 U11556 ( .ip1(\ANSWER/mem[6][3][15] ), .ip2(n9995), .s(n9973), .op(
        n2271) );
  mux2_1 U11557 ( .ip1(\ANSWER/mem[6][4][15] ), .ip2(n9995), .s(n9974), .op(
        n2270) );
  mux2_1 U11558 ( .ip1(\ANSWER/mem[6][5][15] ), .ip2(n9995), .s(n9975), .op(
        n2269) );
  mux2_1 U11559 ( .ip1(\ANSWER/mem[6][6][15] ), .ip2(n9995), .s(n9976), .op(
        n2268) );
  mux2_1 U11560 ( .ip1(\ANSWER/mem[6][7][15] ), .ip2(n9982), .s(n9977), .op(
        n2267) );
  mux2_1 U11561 ( .ip1(\ANSWER/mem[6][8][15] ), .ip2(n9982), .s(n9978), .op(
        n2266) );
  mux2_1 U11562 ( .ip1(\ANSWER/mem[6][9][15] ), .ip2(n9982), .s(n9979), .op(
        n2265) );
  mux2_1 U11563 ( .ip1(\ANSWER/mem[7][0][15] ), .ip2(n9982), .s(n9980), .op(
        n2264) );
  mux2_1 U11564 ( .ip1(\ANSWER/mem[7][1][15] ), .ip2(n9982), .s(n9981), .op(
        n2263) );
  mux2_1 U11565 ( .ip1(\ANSWER/mem[7][2][15] ), .ip2(n9995), .s(n9983), .op(
        n2262) );
  mux2_1 U11566 ( .ip1(\ANSWER/mem[7][3][15] ), .ip2(n9995), .s(n9984), .op(
        n2261) );
  mux2_1 U11567 ( .ip1(\ANSWER/mem[7][4][15] ), .ip2(n9995), .s(n9985), .op(
        n2260) );
  mux2_1 U11568 ( .ip1(\ANSWER/mem[7][5][15] ), .ip2(n9995), .s(n9986), .op(
        n2259) );
  mux2_1 U11569 ( .ip1(\ANSWER/mem[7][6][15] ), .ip2(n9995), .s(n9987), .op(
        n2258) );
  mux2_1 U11570 ( .ip1(\ANSWER/mem[7][7][15] ), .ip2(n9995), .s(n9988), .op(
        n2257) );
  mux2_1 U11571 ( .ip1(\ANSWER/mem[7][8][15] ), .ip2(n9995), .s(n9989), .op(
        n2256) );
  mux2_1 U11572 ( .ip1(\ANSWER/mem[7][9][15] ), .ip2(n9995), .s(n9990), .op(
        n2255) );
  mux2_1 U11573 ( .ip1(\ANSWER/mem[8][0][15] ), .ip2(n9995), .s(n9991), .op(
        n2254) );
  mux2_1 U11574 ( .ip1(\ANSWER/mem[8][1][15] ), .ip2(n9995), .s(n9992), .op(
        n2253) );
  mux2_1 U11575 ( .ip1(\ANSWER/mem[8][2][15] ), .ip2(n9995), .s(n9993), .op(
        n2252) );
  mux2_1 U11576 ( .ip1(\ANSWER/mem[8][3][15] ), .ip2(n9995), .s(n9994), .op(
        n2251) );
  mux2_1 U11577 ( .ip1(\ANSWER/mem[8][4][15] ), .ip2(n9995), .s(n9996), .op(
        n2250) );
  mux2_1 U11578 ( .ip1(\ANSWER/mem[8][5][15] ), .ip2(n10012), .s(n9997), .op(
        n2249) );
  mux2_1 U11579 ( .ip1(\ANSWER/mem[8][6][15] ), .ip2(n9995), .s(n9998), .op(
        n2248) );
  mux2_1 U11580 ( .ip1(\ANSWER/mem[8][7][15] ), .ip2(n10012), .s(n9999), .op(
        n2247) );
  mux2_1 U11581 ( .ip1(\ANSWER/mem[8][8][15] ), .ip2(n9995), .s(n10000), .op(
        n2246) );
  mux2_1 U11582 ( .ip1(\ANSWER/mem[8][9][15] ), .ip2(n10012), .s(n10001), .op(
        n2245) );
  mux2_1 U11583 ( .ip1(\ANSWER/mem[9][0][15] ), .ip2(n9982), .s(n10002), .op(
        n2244) );
  mux2_1 U11584 ( .ip1(\ANSWER/mem[9][1][15] ), .ip2(n9995), .s(n10003), .op(
        n2243) );
  mux2_1 U11585 ( .ip1(\ANSWER/mem[9][2][15] ), .ip2(n10012), .s(n10004), .op(
        n2242) );
  mux2_1 U11586 ( .ip1(\ANSWER/mem[9][3][15] ), .ip2(n9995), .s(n10005), .op(
        n2241) );
  mux2_1 U11587 ( .ip1(\ANSWER/mem[9][4][15] ), .ip2(n10012), .s(n10006), .op(
        n2240) );
  mux2_1 U11588 ( .ip1(\ANSWER/mem[9][5][15] ), .ip2(n9995), .s(n10007), .op(
        n2239) );
  mux2_1 U11589 ( .ip1(\ANSWER/mem[9][6][15] ), .ip2(n10012), .s(n10008), .op(
        n2238) );
  mux2_1 U11590 ( .ip1(\ANSWER/mem[9][7][15] ), .ip2(n10012), .s(n10009), .op(
        n2237) );
  mux2_1 U11591 ( .ip1(\ANSWER/mem[9][8][15] ), .ip2(n10012), .s(n10010), .op(
        n2236) );
  mux2_1 U11592 ( .ip1(\ANSWER/mem[9][9][15] ), .ip2(n10012), .s(n10011), .op(
        n2235) );
  buf_1 U11593 ( .ip(inputSramWe), .op(n10015) );
  buf_1 U11594 ( .ip(n10015), .op(n10013) );
  mux2_1 U11595 ( .ip1(\INPUTSRAM/mem_i[0][0] ), .ip2(pixels[0]), .s(n10013), 
        .op(n2234) );
  mux2_1 U11596 ( .ip1(\INPUTSRAM/mem_i[0][1] ), .ip2(pixels[1]), .s(n10013), 
        .op(n2233) );
  mux2_1 U11597 ( .ip1(\INPUTSRAM/mem_i[0][2] ), .ip2(pixels[2]), .s(n10013), 
        .op(n2232) );
  mux2_1 U11598 ( .ip1(\INPUTSRAM/mem_i[0][3] ), .ip2(pixels[3]), .s(n10013), 
        .op(n2231) );
  mux2_1 U11599 ( .ip1(\INPUTSRAM/mem_i[0][4] ), .ip2(pixels[4]), .s(n10013), 
        .op(n2230) );
  mux2_1 U11600 ( .ip1(\INPUTSRAM/mem_i[0][5] ), .ip2(pixels[5]), .s(n10013), 
        .op(n2229) );
  mux2_1 U11601 ( .ip1(\INPUTSRAM/mem_i[0][6] ), .ip2(pixels[6]), .s(n10013), 
        .op(n2228) );
  mux2_1 U11602 ( .ip1(\INPUTSRAM/mem_i[0][7] ), .ip2(pixels[7]), .s(n10013), 
        .op(n2227) );
  mux2_1 U11603 ( .ip1(\INPUTSRAM/mem_i[0][8] ), .ip2(pixels[8]), .s(n10013), 
        .op(n2226) );
  mux2_1 U11604 ( .ip1(\INPUTSRAM/mem_i[1][0] ), .ip2(pixels[9]), .s(n10013), 
        .op(n2225) );
  mux2_1 U11605 ( .ip1(\INPUTSRAM/mem_i[1][1] ), .ip2(pixels[10]), .s(n10013), 
        .op(n2224) );
  mux2_1 U11606 ( .ip1(\INPUTSRAM/mem_i[1][2] ), .ip2(pixels[11]), .s(n10013), 
        .op(n2223) );
  mux2_1 U11607 ( .ip1(\INPUTSRAM/mem_i[1][3] ), .ip2(pixels[12]), .s(n10013), 
        .op(n2222) );
  buf_1 U11608 ( .ip(n10015), .op(n10014) );
  mux2_1 U11609 ( .ip1(\INPUTSRAM/mem_i[1][4] ), .ip2(pixels[13]), .s(n10014), 
        .op(n2221) );
  mux2_1 U11610 ( .ip1(\INPUTSRAM/mem_i[1][5] ), .ip2(pixels[14]), .s(n10014), 
        .op(n2220) );
  mux2_1 U11611 ( .ip1(\INPUTSRAM/mem_i[1][6] ), .ip2(pixels[15]), .s(n10014), 
        .op(n2219) );
  mux2_1 U11612 ( .ip1(\INPUTSRAM/mem_i[1][7] ), .ip2(pixels[16]), .s(n10014), 
        .op(n2218) );
  mux2_1 U11613 ( .ip1(\INPUTSRAM/mem_i[1][8] ), .ip2(pixels[17]), .s(n10014), 
        .op(n2217) );
  mux2_1 U11614 ( .ip1(\INPUTSRAM/mem_i[2][0] ), .ip2(pixels[18]), .s(n10014), 
        .op(n2216) );
  mux2_1 U11615 ( .ip1(\INPUTSRAM/mem_i[2][1] ), .ip2(pixels[19]), .s(n10014), 
        .op(n2215) );
  mux2_1 U11616 ( .ip1(\INPUTSRAM/mem_i[2][2] ), .ip2(pixels[20]), .s(n10014), 
        .op(n2214) );
  mux2_1 U11617 ( .ip1(\INPUTSRAM/mem_i[2][3] ), .ip2(pixels[21]), .s(n10014), 
        .op(n2213) );
  mux2_1 U11618 ( .ip1(\INPUTSRAM/mem_i[2][4] ), .ip2(pixels[22]), .s(n10014), 
        .op(n2212) );
  mux2_1 U11619 ( .ip1(\INPUTSRAM/mem_i[2][5] ), .ip2(pixels[23]), .s(n10014), 
        .op(n2211) );
  mux2_1 U11620 ( .ip1(\INPUTSRAM/mem_i[2][6] ), .ip2(pixels[24]), .s(n10014), 
        .op(n2210) );
  mux2_1 U11621 ( .ip1(\INPUTSRAM/mem_i[2][7] ), .ip2(pixels[25]), .s(n10014), 
        .op(n2209) );
  mux2_1 U11622 ( .ip1(\INPUTSRAM/mem_i[2][8] ), .ip2(pixels[26]), .s(n10015), 
        .op(n2208) );
  mux2_1 U11623 ( .ip1(\INPUTSRAM/mem_i[3][0] ), .ip2(pixels[27]), .s(
        inputSramWe), .op(n2207) );
  buf_1 U11624 ( .ip(n10015), .op(n10016) );
  mux2_1 U11625 ( .ip1(\INPUTSRAM/mem_i[3][1] ), .ip2(pixels[28]), .s(n10016), 
        .op(n2206) );
  mux2_1 U11626 ( .ip1(\INPUTSRAM/mem_i[3][2] ), .ip2(pixels[29]), .s(n10013), 
        .op(n2205) );
  mux2_1 U11627 ( .ip1(\INPUTSRAM/mem_i[3][3] ), .ip2(pixels[30]), .s(n10014), 
        .op(n2204) );
  mux2_1 U11628 ( .ip1(\INPUTSRAM/mem_i[3][4] ), .ip2(pixels[31]), .s(n10015), 
        .op(n2203) );
  mux2_1 U11629 ( .ip1(\INPUTSRAM/mem_i[3][5] ), .ip2(pixels[32]), .s(
        inputSramWe), .op(n2202) );
  mux2_1 U11630 ( .ip1(\INPUTSRAM/mem_i[3][6] ), .ip2(pixels[33]), .s(n10016), 
        .op(n2201) );
  mux2_1 U11631 ( .ip1(\INPUTSRAM/mem_i[3][7] ), .ip2(pixels[34]), .s(n10013), 
        .op(n2200) );
  mux2_1 U11632 ( .ip1(\INPUTSRAM/mem_i[3][8] ), .ip2(pixels[35]), .s(n10014), 
        .op(n2199) );
  mux2_1 U11633 ( .ip1(\INPUTSRAM/mem_i[4][0] ), .ip2(pixels[36]), .s(n10015), 
        .op(n2198) );
  mux2_1 U11634 ( .ip1(\INPUTSRAM/mem_i[4][1] ), .ip2(pixels[37]), .s(
        inputSramWe), .op(n2197) );
  mux2_1 U11635 ( .ip1(\INPUTSRAM/mem_i[4][2] ), .ip2(pixels[38]), .s(n10016), 
        .op(n2196) );
  mux2_1 U11636 ( .ip1(\INPUTSRAM/mem_i[4][3] ), .ip2(pixels[39]), .s(n10015), 
        .op(n2195) );
  mux2_1 U11637 ( .ip1(\INPUTSRAM/mem_i[4][4] ), .ip2(pixels[40]), .s(n10015), 
        .op(n2194) );
  mux2_1 U11638 ( .ip1(\INPUTSRAM/mem_i[4][5] ), .ip2(pixels[41]), .s(n10015), 
        .op(n2193) );
  mux2_1 U11639 ( .ip1(\INPUTSRAM/mem_i[4][6] ), .ip2(pixels[42]), .s(n10015), 
        .op(n2192) );
  mux2_1 U11640 ( .ip1(\INPUTSRAM/mem_i[4][7] ), .ip2(pixels[43]), .s(n10016), 
        .op(n2191) );
  mux2_1 U11641 ( .ip1(\INPUTSRAM/mem_i[4][8] ), .ip2(pixels[44]), .s(n10013), 
        .op(n2190) );
  mux2_1 U11642 ( .ip1(\INPUTSRAM/mem_i[5][0] ), .ip2(pixels[45]), .s(n10014), 
        .op(n2189) );
  mux2_1 U11643 ( .ip1(\INPUTSRAM/mem_i[5][1] ), .ip2(pixels[46]), .s(n10015), 
        .op(n2188) );
  mux2_1 U11644 ( .ip1(\INPUTSRAM/mem_i[5][2] ), .ip2(pixels[47]), .s(n10015), 
        .op(n2187) );
  mux2_1 U11645 ( .ip1(\INPUTSRAM/mem_i[5][3] ), .ip2(pixels[48]), .s(
        inputSramWe), .op(n2186) );
  mux2_1 U11646 ( .ip1(\INPUTSRAM/mem_i[5][4] ), .ip2(pixels[49]), .s(n10016), 
        .op(n2185) );
  mux2_1 U11647 ( .ip1(\INPUTSRAM/mem_i[5][5] ), .ip2(pixels[50]), .s(n10013), 
        .op(n2184) );
  mux2_1 U11648 ( .ip1(\INPUTSRAM/mem_i[5][6] ), .ip2(pixels[51]), .s(n10014), 
        .op(n2183) );
  mux2_1 U11649 ( .ip1(\INPUTSRAM/mem_i[5][7] ), .ip2(pixels[52]), .s(n10015), 
        .op(n2182) );
  mux2_1 U11650 ( .ip1(\INPUTSRAM/mem_i[5][8] ), .ip2(pixels[53]), .s(n10015), 
        .op(n2181) );
  mux2_1 U11651 ( .ip1(\INPUTSRAM/mem_i[6][0] ), .ip2(pixels[54]), .s(n10015), 
        .op(n2180) );
  mux2_1 U11652 ( .ip1(\INPUTSRAM/mem_i[6][1] ), .ip2(pixels[55]), .s(
        inputSramWe), .op(n2179) );
  mux2_1 U11653 ( .ip1(\INPUTSRAM/mem_i[6][2] ), .ip2(pixels[56]), .s(n10015), 
        .op(n2178) );
  mux2_1 U11654 ( .ip1(\INPUTSRAM/mem_i[6][3] ), .ip2(pixels[57]), .s(
        inputSramWe), .op(n2177) );
  mux2_1 U11655 ( .ip1(\INPUTSRAM/mem_i[6][4] ), .ip2(pixels[58]), .s(n10016), 
        .op(n2176) );
  mux2_1 U11656 ( .ip1(\INPUTSRAM/mem_i[6][5] ), .ip2(pixels[59]), .s(n10013), 
        .op(n2175) );
  mux2_1 U11657 ( .ip1(\INPUTSRAM/mem_i[6][6] ), .ip2(pixels[60]), .s(n10014), 
        .op(n2174) );
  mux2_1 U11658 ( .ip1(\INPUTSRAM/mem_i[6][7] ), .ip2(pixels[61]), .s(n10015), 
        .op(n2173) );
  mux2_1 U11659 ( .ip1(\INPUTSRAM/mem_i[6][8] ), .ip2(pixels[62]), .s(n10015), 
        .op(n2172) );
  mux2_1 U11660 ( .ip1(\INPUTSRAM/mem_i[7][0] ), .ip2(pixels[63]), .s(n10015), 
        .op(n2171) );
  mux2_1 U11661 ( .ip1(\INPUTSRAM/mem_i[7][1] ), .ip2(pixels[64]), .s(
        inputSramWe), .op(n2170) );
  mux2_1 U11662 ( .ip1(\INPUTSRAM/mem_i[7][2] ), .ip2(pixels[65]), .s(
        inputSramWe), .op(n2169) );
  mux2_1 U11663 ( .ip1(\INPUTSRAM/mem_i[7][3] ), .ip2(pixels[66]), .s(
        inputSramWe), .op(n2168) );
  mux2_1 U11664 ( .ip1(\INPUTSRAM/mem_i[7][4] ), .ip2(pixels[67]), .s(
        inputSramWe), .op(n2167) );
  mux2_1 U11665 ( .ip1(\INPUTSRAM/mem_i[7][5] ), .ip2(pixels[68]), .s(
        inputSramWe), .op(n2166) );
  mux2_1 U11666 ( .ip1(\INPUTSRAM/mem_i[7][6] ), .ip2(pixels[69]), .s(
        inputSramWe), .op(n2165) );
  mux2_1 U11667 ( .ip1(\INPUTSRAM/mem_i[7][7] ), .ip2(pixels[70]), .s(
        inputSramWe), .op(n2164) );
  mux2_1 U11668 ( .ip1(\INPUTSRAM/mem_i[7][8] ), .ip2(pixels[71]), .s(
        inputSramWe), .op(n2163) );
  mux2_1 U11669 ( .ip1(\INPUTSRAM/mem_i[8][0] ), .ip2(pixels[72]), .s(
        inputSramWe), .op(n2162) );
  mux2_1 U11670 ( .ip1(\INPUTSRAM/mem_i[8][1] ), .ip2(pixels[73]), .s(
        inputSramWe), .op(n2161) );
  mux2_1 U11671 ( .ip1(\INPUTSRAM/mem_i[8][2] ), .ip2(pixels[74]), .s(
        inputSramWe), .op(n2160) );
  mux2_1 U11672 ( .ip1(\INPUTSRAM/mem_i[8][3] ), .ip2(pixels[75]), .s(n10015), 
        .op(n2159) );
  mux2_1 U11673 ( .ip1(\INPUTSRAM/mem_i[8][4] ), .ip2(pixels[76]), .s(
        inputSramWe), .op(n2158) );
  mux2_1 U11674 ( .ip1(\INPUTSRAM/mem_i[8][5] ), .ip2(pixels[77]), .s(n10016), 
        .op(n2157) );
  mux2_1 U11675 ( .ip1(\INPUTSRAM/mem_i[8][6] ), .ip2(pixels[78]), .s(n10016), 
        .op(n2156) );
  mux2_1 U11676 ( .ip1(\INPUTSRAM/mem_i[8][7] ), .ip2(pixels[79]), .s(n10016), 
        .op(n2155) );
  mux2_1 U11677 ( .ip1(\INPUTSRAM/mem_i[8][8] ), .ip2(pixels[80]), .s(n10016), 
        .op(n2154) );
  mux2_1 U11678 ( .ip1(\INPUTSRAM/mem_i[9][0] ), .ip2(pixels[81]), .s(n10016), 
        .op(n2153) );
  mux2_1 U11679 ( .ip1(\INPUTSRAM/mem_i[9][1] ), .ip2(pixels[82]), .s(n10016), 
        .op(n2152) );
  mux2_1 U11680 ( .ip1(\INPUTSRAM/mem_i[9][2] ), .ip2(pixels[83]), .s(n10016), 
        .op(n2151) );
  mux2_1 U11681 ( .ip1(\INPUTSRAM/mem_i[9][3] ), .ip2(pixels[84]), .s(n10016), 
        .op(n2150) );
  mux2_1 U11682 ( .ip1(\INPUTSRAM/mem_i[9][4] ), .ip2(pixels[85]), .s(n10016), 
        .op(n2149) );
  mux2_1 U11683 ( .ip1(\INPUTSRAM/mem_i[9][5] ), .ip2(pixels[86]), .s(n10016), 
        .op(n2148) );
  mux2_1 U11684 ( .ip1(\INPUTSRAM/mem_i[9][6] ), .ip2(pixels[87]), .s(n10016), 
        .op(n2147) );
  mux2_1 U11685 ( .ip1(\INPUTSRAM/mem_i[9][7] ), .ip2(pixels[88]), .s(n10016), 
        .op(n2146) );
  mux2_1 U11686 ( .ip1(\INPUTSRAM/mem_i[9][8] ), .ip2(pixels[89]), .s(n10016), 
        .op(n2145) );
  inv_1 U11687 ( .ip(n10017), .op(n10478) );
  nand2_1 U11688 ( .ip1(column[8]), .ip2(n10478), .op(n10022) );
  nand2_1 U11689 ( .ip1(n10053), .ip2(n10435), .op(n10432) );
  nand2_1 U11690 ( .ip1(\ROUTEDATA/regData [8]), .ip2(n10432), .op(n10021) );
  inv_1 U11691 ( .ip(n10018), .op(n10434) );
  nand2_1 U11692 ( .ip1(n10434), .ip2(n10019), .op(n10058) );
  inv_1 U11693 ( .ip(n10058), .op(n10054) );
  nand2_1 U11694 ( .ip1(n10054), .ip2(n10435), .op(n10020) );
  nand3_1 U11695 ( .ip1(n10022), .ip2(n10021), .ip3(n10020), .op(n2128) );
  buf_1 U11696 ( .ip(n10478), .op(n10472) );
  buf_1 U11697 ( .ip(n10472), .op(n10485) );
  or2_1 U11698 ( .ip1(n10485), .ip2(n10023), .op(n10440) );
  nand2_1 U11699 ( .ip1(n10053), .ip2(n10440), .op(n10439) );
  nand2_1 U11700 ( .ip1(\ROUTEDATA/regData [24]), .ip2(n10439), .op(n10027) );
  nand2_1 U11701 ( .ip1(n10485), .ip2(column[24]), .op(n10024) );
  nand2_1 U11702 ( .ip1(n10024), .ip2(n10058), .op(n10025) );
  nand2_1 U11703 ( .ip1(n10025), .ip2(n10440), .op(n10026) );
  nand2_1 U11704 ( .ip1(n10027), .ip2(n10026), .op(n2127) );
  nand2_1 U11705 ( .ip1(column[40]), .ip2(n10478), .op(n10031) );
  buf_1 U11706 ( .ip(n10472), .op(n10444) );
  or2_1 U11707 ( .ip1(n10444), .ip2(n10028), .op(n10445) );
  nand2_1 U11708 ( .ip1(n10053), .ip2(n10445), .op(n10446) );
  nand2_1 U11709 ( .ip1(\ROUTEDATA/regData [40]), .ip2(n10446), .op(n10030) );
  nand2_1 U11710 ( .ip1(n10054), .ip2(n10445), .op(n10029) );
  nand3_1 U11711 ( .ip1(n10031), .ip2(n10030), .ip3(n10029), .op(n2126) );
  nand2_1 U11712 ( .ip1(column[56]), .ip2(n10444), .op(n10035) );
  or2_1 U11713 ( .ip1(n10444), .ip2(n10032), .op(n10452) );
  nand2_1 U11714 ( .ip1(n10054), .ip2(n10452), .op(n10034) );
  nand2_1 U11715 ( .ip1(n10053), .ip2(n10452), .op(n10450) );
  nand2_1 U11716 ( .ip1(\ROUTEDATA/regData [56]), .ip2(n10450), .op(n10033) );
  nand3_1 U11717 ( .ip1(n10035), .ip2(n10034), .ip3(n10033), .op(n2125) );
  nand2_1 U11718 ( .ip1(column[72]), .ip2(n10478), .op(n10039) );
  nor2_1 U11719 ( .ip1(n10485), .ip2(n10036), .op(n10412) );
  inv_1 U11720 ( .ip(n10412), .op(n10456) );
  nand2_1 U11721 ( .ip1(n10053), .ip2(n10456), .op(n10457) );
  nand2_1 U11722 ( .ip1(\ROUTEDATA/regData [72]), .ip2(n10457), .op(n10038) );
  nand2_1 U11723 ( .ip1(n10054), .ip2(n10456), .op(n10037) );
  nand3_1 U11724 ( .ip1(n10039), .ip2(n10038), .ip3(n10037), .op(n2124) );
  nand2_1 U11725 ( .ip1(column[88]), .ip2(n10444), .op(n10043) );
  or2_1 U11726 ( .ip1(n10444), .ip2(n10040), .op(n10461) );
  nand2_1 U11727 ( .ip1(n10053), .ip2(n10461), .op(n10462) );
  nand2_1 U11728 ( .ip1(\ROUTEDATA/regData [88]), .ip2(n10462), .op(n10042) );
  nand2_1 U11729 ( .ip1(n10054), .ip2(n10461), .op(n10041) );
  nand3_1 U11730 ( .ip1(n10043), .ip2(n10042), .ip3(n10041), .op(n2123) );
  nand2_1 U11731 ( .ip1(column[104]), .ip2(n10444), .op(n10047) );
  or2_1 U11732 ( .ip1(n10444), .ip2(n10044), .op(n10466) );
  nand2_1 U11733 ( .ip1(n10054), .ip2(n10466), .op(n10046) );
  nand2_1 U11734 ( .ip1(n10053), .ip2(n10466), .op(n10467) );
  nand2_1 U11735 ( .ip1(\ROUTEDATA/regData [104]), .ip2(n10467), .op(n10045)
         );
  nand3_1 U11736 ( .ip1(n10047), .ip2(n10046), .ip3(n10045), .op(n2122) );
  nand2_1 U11737 ( .ip1(column[120]), .ip2(n10478), .op(n10051) );
  or2_1 U11738 ( .ip1(n10485), .ip2(n10048), .op(n10474) );
  nand2_1 U11739 ( .ip1(n10054), .ip2(n10474), .op(n10050) );
  nand2_1 U11740 ( .ip1(n10053), .ip2(n10474), .op(n10471) );
  nand2_1 U11741 ( .ip1(\ROUTEDATA/regData [120]), .ip2(n10471), .op(n10049)
         );
  nand3_1 U11742 ( .ip1(n10051), .ip2(n10050), .ip3(n10049), .op(n2121) );
  nand2_1 U11743 ( .ip1(column[136]), .ip2(n10472), .op(n10057) );
  or2_1 U11744 ( .ip1(n10444), .ip2(n10052), .op(n10480) );
  nand2_1 U11745 ( .ip1(n10053), .ip2(n10480), .op(n10479) );
  nand2_1 U11746 ( .ip1(\ROUTEDATA/regData [136]), .ip2(n10479), .op(n10056)
         );
  nand2_1 U11747 ( .ip1(n10054), .ip2(n10480), .op(n10055) );
  nand3_1 U11748 ( .ip1(n10057), .ip2(n10056), .ip3(n10055), .op(n2120) );
  nand2_1 U11749 ( .ip1(n10485), .ip2(column[152]), .op(n10059) );
  nand2_1 U11750 ( .ip1(n10059), .ip2(n10058), .op(n10060) );
  nor2_1 U11751 ( .ip1(n10485), .ip2(weight2_loadNextRow), .op(n10488) );
  mux2_1 U11752 ( .ip1(n10060), .ip2(\ROUTEDATA/regData [152]), .s(n10488), 
        .op(n2119) );
  nand2_1 U11753 ( .ip1(n10485), .ip2(column[9]), .op(n10062) );
  nand2_1 U11754 ( .ip1(\ROUTEDATA/regData [9]), .ip2(n10432), .op(n10061) );
  nand2_1 U11755 ( .ip1(n10062), .ip2(n10061), .op(n2118) );
  nand2_1 U11756 ( .ip1(n10485), .ip2(column[25]), .op(n10064) );
  nand2_1 U11757 ( .ip1(\ROUTEDATA/regData [25]), .ip2(n10439), .op(n10063) );
  nand2_1 U11758 ( .ip1(n10064), .ip2(n10063), .op(n2117) );
  nand2_1 U11759 ( .ip1(n10485), .ip2(column[41]), .op(n10066) );
  nand2_1 U11760 ( .ip1(\ROUTEDATA/regData [41]), .ip2(n10446), .op(n10065) );
  nand2_1 U11761 ( .ip1(n10066), .ip2(n10065), .op(n2116) );
  nand2_1 U11762 ( .ip1(n10485), .ip2(column[57]), .op(n10068) );
  nand2_1 U11763 ( .ip1(\ROUTEDATA/regData [57]), .ip2(n10450), .op(n10067) );
  nand2_1 U11764 ( .ip1(n10068), .ip2(n10067), .op(n2115) );
  nand2_1 U11765 ( .ip1(n10485), .ip2(column[73]), .op(n10070) );
  nand2_1 U11766 ( .ip1(\ROUTEDATA/regData [73]), .ip2(n10457), .op(n10069) );
  nand2_1 U11767 ( .ip1(n10070), .ip2(n10069), .op(n2114) );
  nand2_1 U11768 ( .ip1(n10485), .ip2(column[89]), .op(n10072) );
  nand2_1 U11769 ( .ip1(\ROUTEDATA/regData [89]), .ip2(n10462), .op(n10071) );
  nand2_1 U11770 ( .ip1(n10072), .ip2(n10071), .op(n2113) );
  nand2_1 U11771 ( .ip1(n10485), .ip2(column[105]), .op(n10074) );
  nand2_1 U11772 ( .ip1(\ROUTEDATA/regData [105]), .ip2(n10467), .op(n10073)
         );
  nand2_1 U11773 ( .ip1(n10074), .ip2(n10073), .op(n2112) );
  nand2_1 U11774 ( .ip1(n10485), .ip2(column[121]), .op(n10076) );
  nand2_1 U11775 ( .ip1(\ROUTEDATA/regData [121]), .ip2(n10471), .op(n10075)
         );
  nand2_1 U11776 ( .ip1(n10076), .ip2(n10075), .op(n2111) );
  nand2_1 U11777 ( .ip1(n10472), .ip2(column[137]), .op(n10078) );
  nand2_1 U11778 ( .ip1(\ROUTEDATA/regData [137]), .ip2(n10479), .op(n10077)
         );
  nand2_1 U11779 ( .ip1(n10078), .ip2(n10077), .op(n2110) );
  nand2_1 U11780 ( .ip1(n10488), .ip2(\ROUTEDATA/regData [153]), .op(n10080)
         );
  nand2_1 U11781 ( .ip1(column[153]), .ip2(n10485), .op(n10079) );
  nand2_1 U11782 ( .ip1(n10080), .ip2(n10079), .op(n2109) );
  nand2_1 U11783 ( .ip1(n10472), .ip2(column[10]), .op(n10082) );
  nand2_1 U11784 ( .ip1(\ROUTEDATA/regData [10]), .ip2(n10432), .op(n10081) );
  nand2_1 U11785 ( .ip1(n10082), .ip2(n10081), .op(n2108) );
  nand2_1 U11786 ( .ip1(n10472), .ip2(column[26]), .op(n10084) );
  nand2_1 U11787 ( .ip1(\ROUTEDATA/regData [26]), .ip2(n10439), .op(n10083) );
  nand2_1 U11788 ( .ip1(n10084), .ip2(n10083), .op(n2107) );
  nand2_1 U11789 ( .ip1(n10472), .ip2(column[42]), .op(n10086) );
  nand2_1 U11790 ( .ip1(\ROUTEDATA/regData [42]), .ip2(n10446), .op(n10085) );
  nand2_1 U11791 ( .ip1(n10086), .ip2(n10085), .op(n2106) );
  nand2_1 U11792 ( .ip1(n10472), .ip2(column[58]), .op(n10088) );
  nand2_1 U11793 ( .ip1(\ROUTEDATA/regData [58]), .ip2(n10450), .op(n10087) );
  nand2_1 U11794 ( .ip1(n10088), .ip2(n10087), .op(n2105) );
  nand2_1 U11795 ( .ip1(n10472), .ip2(column[74]), .op(n10090) );
  nand2_1 U11796 ( .ip1(\ROUTEDATA/regData [74]), .ip2(n10457), .op(n10089) );
  nand2_1 U11797 ( .ip1(n10090), .ip2(n10089), .op(n2104) );
  nand2_1 U11798 ( .ip1(n10472), .ip2(column[90]), .op(n10092) );
  nand2_1 U11799 ( .ip1(\ROUTEDATA/regData [90]), .ip2(n10462), .op(n10091) );
  nand2_1 U11800 ( .ip1(n10092), .ip2(n10091), .op(n2103) );
  nand2_1 U11801 ( .ip1(n10472), .ip2(column[106]), .op(n10094) );
  nand2_1 U11802 ( .ip1(\ROUTEDATA/regData [106]), .ip2(n10467), .op(n10093)
         );
  nand2_1 U11803 ( .ip1(n10094), .ip2(n10093), .op(n2102) );
  nand2_1 U11804 ( .ip1(n10472), .ip2(column[122]), .op(n10096) );
  nand2_1 U11805 ( .ip1(\ROUTEDATA/regData [122]), .ip2(n10471), .op(n10095)
         );
  nand2_1 U11806 ( .ip1(n10096), .ip2(n10095), .op(n2101) );
  nand2_1 U11807 ( .ip1(n10472), .ip2(column[138]), .op(n10098) );
  nand2_1 U11808 ( .ip1(\ROUTEDATA/regData [138]), .ip2(n10479), .op(n10097)
         );
  nand2_1 U11809 ( .ip1(n10098), .ip2(n10097), .op(n2100) );
  nand2_1 U11810 ( .ip1(n10488), .ip2(\ROUTEDATA/regData [154]), .op(n10100)
         );
  nand2_1 U11811 ( .ip1(column[154]), .ip2(n10444), .op(n10099) );
  nand2_1 U11812 ( .ip1(n10100), .ip2(n10099), .op(n2099) );
  nand2_1 U11813 ( .ip1(n10472), .ip2(column[11]), .op(n10102) );
  nand2_1 U11814 ( .ip1(\ROUTEDATA/regData [11]), .ip2(n10432), .op(n10101) );
  nand2_1 U11815 ( .ip1(n10102), .ip2(n10101), .op(n2098) );
  nand2_1 U11816 ( .ip1(n10472), .ip2(column[27]), .op(n10104) );
  nand2_1 U11817 ( .ip1(\ROUTEDATA/regData [27]), .ip2(n10439), .op(n10103) );
  nand2_1 U11818 ( .ip1(n10104), .ip2(n10103), .op(n2097) );
  nand2_1 U11819 ( .ip1(n10472), .ip2(column[43]), .op(n10106) );
  nand2_1 U11820 ( .ip1(\ROUTEDATA/regData [43]), .ip2(n10446), .op(n10105) );
  nand2_1 U11821 ( .ip1(n10106), .ip2(n10105), .op(n2096) );
  nand2_1 U11822 ( .ip1(n10485), .ip2(column[59]), .op(n10108) );
  nand2_1 U11823 ( .ip1(\ROUTEDATA/regData [59]), .ip2(n10450), .op(n10107) );
  nand2_1 U11824 ( .ip1(n10108), .ip2(n10107), .op(n2095) );
  nand2_1 U11825 ( .ip1(n10478), .ip2(column[75]), .op(n10110) );
  nand2_1 U11826 ( .ip1(\ROUTEDATA/regData [75]), .ip2(n10457), .op(n10109) );
  nand2_1 U11827 ( .ip1(n10110), .ip2(n10109), .op(n2094) );
  nand2_1 U11828 ( .ip1(n10478), .ip2(column[91]), .op(n10112) );
  nand2_1 U11829 ( .ip1(\ROUTEDATA/regData [91]), .ip2(n10462), .op(n10111) );
  nand2_1 U11830 ( .ip1(n10112), .ip2(n10111), .op(n2093) );
  nand2_1 U11831 ( .ip1(n10478), .ip2(column[107]), .op(n10114) );
  nand2_1 U11832 ( .ip1(\ROUTEDATA/regData [107]), .ip2(n10467), .op(n10113)
         );
  nand2_1 U11833 ( .ip1(n10114), .ip2(n10113), .op(n2092) );
  nand2_1 U11834 ( .ip1(n10472), .ip2(column[123]), .op(n10116) );
  nand2_1 U11835 ( .ip1(\ROUTEDATA/regData [123]), .ip2(n10471), .op(n10115)
         );
  nand2_1 U11836 ( .ip1(n10116), .ip2(n10115), .op(n2091) );
  nand2_1 U11837 ( .ip1(n10478), .ip2(column[139]), .op(n10118) );
  nand2_1 U11838 ( .ip1(\ROUTEDATA/regData [139]), .ip2(n10479), .op(n10117)
         );
  nand2_1 U11839 ( .ip1(n10118), .ip2(n10117), .op(n2090) );
  nand2_1 U11840 ( .ip1(n10488), .ip2(\ROUTEDATA/regData [155]), .op(n10120)
         );
  nand2_1 U11841 ( .ip1(column[155]), .ip2(n10478), .op(n10119) );
  nand2_1 U11842 ( .ip1(n10120), .ip2(n10119), .op(n2089) );
  nand2_1 U11843 ( .ip1(n10485), .ip2(column[12]), .op(n10122) );
  nand2_1 U11844 ( .ip1(\ROUTEDATA/regData [12]), .ip2(n10432), .op(n10121) );
  nand2_1 U11845 ( .ip1(n10122), .ip2(n10121), .op(n2088) );
  nand2_1 U11846 ( .ip1(n10478), .ip2(column[28]), .op(n10124) );
  nand2_1 U11847 ( .ip1(\ROUTEDATA/regData [28]), .ip2(n10439), .op(n10123) );
  nand2_1 U11848 ( .ip1(n10124), .ip2(n10123), .op(n2087) );
  nand2_1 U11849 ( .ip1(n10472), .ip2(column[44]), .op(n10126) );
  nand2_1 U11850 ( .ip1(\ROUTEDATA/regData [44]), .ip2(n10446), .op(n10125) );
  nand2_1 U11851 ( .ip1(n10126), .ip2(n10125), .op(n2086) );
  nand2_1 U11852 ( .ip1(n10478), .ip2(column[60]), .op(n10128) );
  nand2_1 U11853 ( .ip1(\ROUTEDATA/regData [60]), .ip2(n10450), .op(n10127) );
  nand2_1 U11854 ( .ip1(n10128), .ip2(n10127), .op(n2085) );
  nand2_1 U11855 ( .ip1(n10478), .ip2(column[76]), .op(n10130) );
  nand2_1 U11856 ( .ip1(\ROUTEDATA/regData [76]), .ip2(n10457), .op(n10129) );
  nand2_1 U11857 ( .ip1(n10130), .ip2(n10129), .op(n2084) );
  nand2_1 U11858 ( .ip1(column[92]), .ip2(n10478), .op(n10132) );
  nand2_1 U11859 ( .ip1(\ROUTEDATA/regData [92]), .ip2(n10462), .op(n10131) );
  nand2_1 U11860 ( .ip1(n10132), .ip2(n10131), .op(n2083) );
  nand2_1 U11861 ( .ip1(n10485), .ip2(column[108]), .op(n10134) );
  nand2_1 U11862 ( .ip1(\ROUTEDATA/regData [108]), .ip2(n10467), .op(n10133)
         );
  nand2_1 U11863 ( .ip1(n10134), .ip2(n10133), .op(n2082) );
  nand2_1 U11864 ( .ip1(n10478), .ip2(column[124]), .op(n10136) );
  nand2_1 U11865 ( .ip1(\ROUTEDATA/regData [124]), .ip2(n10471), .op(n10135)
         );
  nand2_1 U11866 ( .ip1(n10136), .ip2(n10135), .op(n2081) );
  nand2_1 U11867 ( .ip1(n10478), .ip2(column[140]), .op(n10138) );
  nand2_1 U11868 ( .ip1(\ROUTEDATA/regData [140]), .ip2(n10479), .op(n10137)
         );
  nand2_1 U11869 ( .ip1(n10138), .ip2(n10137), .op(n2080) );
  nand2_1 U11870 ( .ip1(n10488), .ip2(\ROUTEDATA/regData [156]), .op(n10140)
         );
  nand2_1 U11871 ( .ip1(column[156]), .ip2(n10478), .op(n10139) );
  nand2_1 U11872 ( .ip1(n10140), .ip2(n10139), .op(n2079) );
  nand2_1 U11873 ( .ip1(n10478), .ip2(column[13]), .op(n10142) );
  nand2_1 U11874 ( .ip1(\ROUTEDATA/regData [13]), .ip2(n10432), .op(n10141) );
  nand2_1 U11875 ( .ip1(n10142), .ip2(n10141), .op(n2078) );
  nand2_1 U11876 ( .ip1(n10444), .ip2(column[29]), .op(n10144) );
  nand2_1 U11877 ( .ip1(\ROUTEDATA/regData [29]), .ip2(n10439), .op(n10143) );
  nand2_1 U11878 ( .ip1(n10144), .ip2(n10143), .op(n2077) );
  nand2_1 U11879 ( .ip1(n10444), .ip2(column[45]), .op(n10146) );
  nand2_1 U11880 ( .ip1(\ROUTEDATA/regData [45]), .ip2(n10446), .op(n10145) );
  nand2_1 U11881 ( .ip1(n10146), .ip2(n10145), .op(n2076) );
  nand2_1 U11882 ( .ip1(n10478), .ip2(column[61]), .op(n10148) );
  nand2_1 U11883 ( .ip1(\ROUTEDATA/regData [61]), .ip2(n10450), .op(n10147) );
  nand2_1 U11884 ( .ip1(n10148), .ip2(n10147), .op(n2075) );
  nand2_1 U11885 ( .ip1(n10444), .ip2(column[77]), .op(n10150) );
  nand2_1 U11886 ( .ip1(\ROUTEDATA/regData [77]), .ip2(n10457), .op(n10149) );
  nand2_1 U11887 ( .ip1(n10150), .ip2(n10149), .op(n2074) );
  nand2_1 U11888 ( .ip1(n10485), .ip2(column[93]), .op(n10152) );
  nand2_1 U11889 ( .ip1(\ROUTEDATA/regData [93]), .ip2(n10462), .op(n10151) );
  nand2_1 U11890 ( .ip1(n10152), .ip2(n10151), .op(n2073) );
  nand2_1 U11891 ( .ip1(n10444), .ip2(column[109]), .op(n10154) );
  nand2_1 U11892 ( .ip1(\ROUTEDATA/regData [109]), .ip2(n10467), .op(n10153)
         );
  nand2_1 U11893 ( .ip1(n10154), .ip2(n10153), .op(n2072) );
  nand2_1 U11894 ( .ip1(n10478), .ip2(column[125]), .op(n10156) );
  nand2_1 U11895 ( .ip1(\ROUTEDATA/regData [125]), .ip2(n10471), .op(n10155)
         );
  nand2_1 U11896 ( .ip1(n10156), .ip2(n10155), .op(n2071) );
  nand2_1 U11897 ( .ip1(n10478), .ip2(column[141]), .op(n10158) );
  nand2_1 U11898 ( .ip1(\ROUTEDATA/regData [141]), .ip2(n10479), .op(n10157)
         );
  nand2_1 U11899 ( .ip1(n10158), .ip2(n10157), .op(n2070) );
  nand2_1 U11900 ( .ip1(n10488), .ip2(\ROUTEDATA/regData [157]), .op(n10160)
         );
  nand2_1 U11901 ( .ip1(column[157]), .ip2(n10444), .op(n10159) );
  nand2_1 U11902 ( .ip1(n10160), .ip2(n10159), .op(n2069) );
  nand2_1 U11903 ( .ip1(n10478), .ip2(column[14]), .op(n10162) );
  nand2_1 U11904 ( .ip1(\ROUTEDATA/regData [14]), .ip2(n10432), .op(n10161) );
  nand2_1 U11905 ( .ip1(n10162), .ip2(n10161), .op(n2068) );
  nand2_1 U11906 ( .ip1(n10444), .ip2(column[30]), .op(n10164) );
  nand2_1 U11907 ( .ip1(\ROUTEDATA/regData [30]), .ip2(n10439), .op(n10163) );
  nand2_1 U11908 ( .ip1(n10164), .ip2(n10163), .op(n2067) );
  nand2_1 U11909 ( .ip1(n10478), .ip2(column[46]), .op(n10166) );
  nand2_1 U11910 ( .ip1(\ROUTEDATA/regData [46]), .ip2(n10446), .op(n10165) );
  nand2_1 U11911 ( .ip1(n10166), .ip2(n10165), .op(n2066) );
  nand2_1 U11912 ( .ip1(n10472), .ip2(column[62]), .op(n10168) );
  nand2_1 U11913 ( .ip1(\ROUTEDATA/regData [62]), .ip2(n10450), .op(n10167) );
  nand2_1 U11914 ( .ip1(n10168), .ip2(n10167), .op(n2065) );
  nand2_1 U11915 ( .ip1(n10485), .ip2(column[78]), .op(n10170) );
  nand2_1 U11916 ( .ip1(\ROUTEDATA/regData [78]), .ip2(n10457), .op(n10169) );
  nand2_1 U11917 ( .ip1(n10170), .ip2(n10169), .op(n2064) );
  nand2_1 U11918 ( .ip1(n10478), .ip2(column[94]), .op(n10172) );
  nand2_1 U11919 ( .ip1(\ROUTEDATA/regData [94]), .ip2(n10462), .op(n10171) );
  nand2_1 U11920 ( .ip1(n10172), .ip2(n10171), .op(n2063) );
  nand2_1 U11921 ( .ip1(n10472), .ip2(column[110]), .op(n10174) );
  nand2_1 U11922 ( .ip1(\ROUTEDATA/regData [110]), .ip2(n10467), .op(n10173)
         );
  nand2_1 U11923 ( .ip1(n10174), .ip2(n10173), .op(n2062) );
  nand2_1 U11924 ( .ip1(n10478), .ip2(column[126]), .op(n10176) );
  nand2_1 U11925 ( .ip1(\ROUTEDATA/regData [126]), .ip2(n10471), .op(n10175)
         );
  nand2_1 U11926 ( .ip1(n10176), .ip2(n10175), .op(n2061) );
  nand2_1 U11927 ( .ip1(n10478), .ip2(column[142]), .op(n10178) );
  nand2_1 U11928 ( .ip1(\ROUTEDATA/regData [142]), .ip2(n10479), .op(n10177)
         );
  nand2_1 U11929 ( .ip1(n10178), .ip2(n10177), .op(n2060) );
  nand2_1 U11930 ( .ip1(n10488), .ip2(\ROUTEDATA/regData [158]), .op(n10180)
         );
  nand2_1 U11931 ( .ip1(column[158]), .ip2(n10472), .op(n10179) );
  nand2_1 U11932 ( .ip1(n10180), .ip2(n10179), .op(n2059) );
  nand2_1 U11933 ( .ip1(n10472), .ip2(column[15]), .op(n10182) );
  nand2_1 U11934 ( .ip1(\ROUTEDATA/regData [15]), .ip2(n10432), .op(n10181) );
  nand2_1 U11935 ( .ip1(n10182), .ip2(n10181), .op(n2058) );
  nand2_1 U11936 ( .ip1(n10472), .ip2(column[31]), .op(n10184) );
  nand2_1 U11937 ( .ip1(\ROUTEDATA/regData [31]), .ip2(n10439), .op(n10183) );
  nand2_1 U11938 ( .ip1(n10184), .ip2(n10183), .op(n2057) );
  nand2_1 U11939 ( .ip1(n10478), .ip2(column[47]), .op(n10186) );
  nand2_1 U11940 ( .ip1(\ROUTEDATA/regData [47]), .ip2(n10446), .op(n10185) );
  nand2_1 U11941 ( .ip1(n10186), .ip2(n10185), .op(n2056) );
  nand2_1 U11942 ( .ip1(n10472), .ip2(column[63]), .op(n10188) );
  nand2_1 U11943 ( .ip1(\ROUTEDATA/regData [63]), .ip2(n10450), .op(n10187) );
  nand2_1 U11944 ( .ip1(n10188), .ip2(n10187), .op(n2055) );
  nand2_1 U11945 ( .ip1(n10478), .ip2(column[79]), .op(n10190) );
  nand2_1 U11946 ( .ip1(\ROUTEDATA/regData [79]), .ip2(n10457), .op(n10189) );
  nand2_1 U11947 ( .ip1(n10190), .ip2(n10189), .op(n2054) );
  nand2_1 U11948 ( .ip1(n10472), .ip2(column[95]), .op(n10192) );
  nand2_1 U11949 ( .ip1(\ROUTEDATA/regData [95]), .ip2(n10462), .op(n10191) );
  nand2_1 U11950 ( .ip1(n10192), .ip2(n10191), .op(n2053) );
  nand2_1 U11951 ( .ip1(n10472), .ip2(column[111]), .op(n10194) );
  nand2_1 U11952 ( .ip1(\ROUTEDATA/regData [111]), .ip2(n10467), .op(n10193)
         );
  nand2_1 U11953 ( .ip1(n10194), .ip2(n10193), .op(n2052) );
  nand2_1 U11954 ( .ip1(n10478), .ip2(column[127]), .op(n10196) );
  nand2_1 U11955 ( .ip1(\ROUTEDATA/regData [127]), .ip2(n10471), .op(n10195)
         );
  nand2_1 U11956 ( .ip1(n10196), .ip2(n10195), .op(n2051) );
  nand2_1 U11957 ( .ip1(n10472), .ip2(column[143]), .op(n10198) );
  nand2_1 U11958 ( .ip1(\ROUTEDATA/regData [143]), .ip2(n10479), .op(n10197)
         );
  nand2_1 U11959 ( .ip1(n10198), .ip2(n10197), .op(n2050) );
  nand2_1 U11960 ( .ip1(n10488), .ip2(\ROUTEDATA/regData [159]), .op(n10200)
         );
  nand2_1 U11961 ( .ip1(column[159]), .ip2(n10478), .op(n10199) );
  nand2_1 U11962 ( .ip1(n10200), .ip2(n10199), .op(n2049) );
  nand2_1 U11963 ( .ip1(n10444), .ip2(column[0]), .op(n10203) );
  nand2_1 U11964 ( .ip1(\ROUTEDATA/regData [0]), .ip2(n10432), .op(n10202) );
  nand2_1 U11965 ( .ip1(\SIGMOID/N64 ), .ip2(n10434), .op(n10229) );
  inv_1 U11966 ( .ip(n10229), .op(n10225) );
  nand2_1 U11967 ( .ip1(n10225), .ip2(n10435), .op(n10201) );
  nand3_1 U11968 ( .ip1(n10203), .ip2(n10202), .ip3(n10201), .op(n2048) );
  nand2_1 U11969 ( .ip1(n10472), .ip2(column[16]), .op(n10206) );
  nand2_1 U11970 ( .ip1(\ROUTEDATA/regData [16]), .ip2(n10439), .op(n10205) );
  nand2_1 U11971 ( .ip1(n10225), .ip2(n10440), .op(n10204) );
  nand3_1 U11972 ( .ip1(n10206), .ip2(n10205), .ip3(n10204), .op(n2047) );
  nand2_1 U11973 ( .ip1(column[32]), .ip2(n10478), .op(n10209) );
  nand2_1 U11974 ( .ip1(n10225), .ip2(n10445), .op(n10208) );
  nand2_1 U11975 ( .ip1(\ROUTEDATA/regData [32]), .ip2(n10446), .op(n10207) );
  nand3_1 U11976 ( .ip1(n10209), .ip2(n10208), .ip3(n10207), .op(n2046) );
  nand2_1 U11977 ( .ip1(column[48]), .ip2(n10478), .op(n10212) );
  nand2_1 U11978 ( .ip1(n10225), .ip2(n10452), .op(n10211) );
  nand2_1 U11979 ( .ip1(\ROUTEDATA/regData [48]), .ip2(n10450), .op(n10210) );
  nand3_1 U11980 ( .ip1(n10212), .ip2(n10211), .ip3(n10210), .op(n2045) );
  nand2_1 U11981 ( .ip1(column[64]), .ip2(n10478), .op(n10215) );
  nand2_1 U11982 ( .ip1(n10225), .ip2(n10456), .op(n10214) );
  nand2_1 U11983 ( .ip1(\ROUTEDATA/regData [64]), .ip2(n10457), .op(n10213) );
  nand3_1 U11984 ( .ip1(n10215), .ip2(n10214), .ip3(n10213), .op(n2044) );
  nand2_1 U11985 ( .ip1(column[80]), .ip2(n10444), .op(n10218) );
  nand2_1 U11986 ( .ip1(\ROUTEDATA/regData [80]), .ip2(n10462), .op(n10217) );
  nand2_1 U11987 ( .ip1(n10225), .ip2(n10461), .op(n10216) );
  nand3_1 U11988 ( .ip1(n10218), .ip2(n10217), .ip3(n10216), .op(n2043) );
  nand2_1 U11989 ( .ip1(column[96]), .ip2(n10472), .op(n10221) );
  nand2_1 U11990 ( .ip1(\ROUTEDATA/regData [96]), .ip2(n10467), .op(n10220) );
  nand2_1 U11991 ( .ip1(n10225), .ip2(n10466), .op(n10219) );
  nand3_1 U11992 ( .ip1(n10221), .ip2(n10220), .ip3(n10219), .op(n2042) );
  nand2_1 U11993 ( .ip1(column[112]), .ip2(n10485), .op(n10224) );
  nand2_1 U11994 ( .ip1(n10225), .ip2(n10474), .op(n10223) );
  nand2_1 U11995 ( .ip1(\ROUTEDATA/regData [112]), .ip2(n10471), .op(n10222)
         );
  nand3_1 U11996 ( .ip1(n10224), .ip2(n10223), .ip3(n10222), .op(n2041) );
  nand2_1 U11997 ( .ip1(column[128]), .ip2(n10478), .op(n10228) );
  nand2_1 U11998 ( .ip1(\ROUTEDATA/regData [128]), .ip2(n10479), .op(n10227)
         );
  nand2_1 U11999 ( .ip1(n10225), .ip2(n10480), .op(n10226) );
  nand3_1 U12000 ( .ip1(n10228), .ip2(n10227), .ip3(n10226), .op(n2040) );
  nand2_1 U12001 ( .ip1(n10472), .ip2(column[144]), .op(n10230) );
  nand2_1 U12002 ( .ip1(n10230), .ip2(n10229), .op(n10231) );
  mux2_1 U12003 ( .ip1(n10231), .ip2(\ROUTEDATA/regData [144]), .s(n10488), 
        .op(n2039) );
  nand2_1 U12004 ( .ip1(n10485), .ip2(column[1]), .op(n10235) );
  nand2_1 U12005 ( .ip1(\ROUTEDATA/regData [1]), .ip2(n10432), .op(n10234) );
  nand2_1 U12006 ( .ip1(n10434), .ip2(n10232), .op(n10261) );
  inv_1 U12007 ( .ip(n10261), .op(n10257) );
  nand2_1 U12008 ( .ip1(n10257), .ip2(n10435), .op(n10233) );
  nand3_1 U12009 ( .ip1(n10235), .ip2(n10234), .ip3(n10233), .op(n2038) );
  nand2_1 U12010 ( .ip1(n10444), .ip2(column[17]), .op(n10238) );
  nand2_1 U12011 ( .ip1(\ROUTEDATA/regData [17]), .ip2(n10439), .op(n10237) );
  nand2_1 U12012 ( .ip1(n10257), .ip2(n10440), .op(n10236) );
  nand3_1 U12013 ( .ip1(n10238), .ip2(n10237), .ip3(n10236), .op(n2037) );
  nand2_1 U12014 ( .ip1(column[33]), .ip2(n10472), .op(n10241) );
  nand2_1 U12015 ( .ip1(n10257), .ip2(n10445), .op(n10240) );
  nand2_1 U12016 ( .ip1(\ROUTEDATA/regData [33]), .ip2(n10446), .op(n10239) );
  nand3_1 U12017 ( .ip1(n10241), .ip2(n10240), .ip3(n10239), .op(n2036) );
  nand2_1 U12018 ( .ip1(column[49]), .ip2(n10478), .op(n10244) );
  nand2_1 U12019 ( .ip1(\ROUTEDATA/regData [49]), .ip2(n10450), .op(n10243) );
  nand2_1 U12020 ( .ip1(n10257), .ip2(n10452), .op(n10242) );
  nand3_1 U12021 ( .ip1(n10244), .ip2(n10243), .ip3(n10242), .op(n2035) );
  nand2_1 U12022 ( .ip1(column[65]), .ip2(n10485), .op(n10247) );
  nand2_1 U12023 ( .ip1(n10257), .ip2(n10456), .op(n10246) );
  nand2_1 U12024 ( .ip1(\ROUTEDATA/regData [65]), .ip2(n10457), .op(n10245) );
  nand3_1 U12025 ( .ip1(n10247), .ip2(n10246), .ip3(n10245), .op(n2034) );
  nand2_1 U12026 ( .ip1(column[81]), .ip2(n10444), .op(n10250) );
  nand2_1 U12027 ( .ip1(\ROUTEDATA/regData [81]), .ip2(n10462), .op(n10249) );
  nand2_1 U12028 ( .ip1(n10257), .ip2(n10461), .op(n10248) );
  nand3_1 U12029 ( .ip1(n10250), .ip2(n10249), .ip3(n10248), .op(n2033) );
  nand2_1 U12030 ( .ip1(column[97]), .ip2(n10478), .op(n10253) );
  nand2_1 U12031 ( .ip1(\ROUTEDATA/regData [97]), .ip2(n10467), .op(n10252) );
  nand2_1 U12032 ( .ip1(n10257), .ip2(n10466), .op(n10251) );
  nand3_1 U12033 ( .ip1(n10253), .ip2(n10252), .ip3(n10251), .op(n2032) );
  nand2_1 U12034 ( .ip1(column[113]), .ip2(n10444), .op(n10256) );
  nand2_1 U12035 ( .ip1(\ROUTEDATA/regData [113]), .ip2(n10471), .op(n10255)
         );
  nand2_1 U12036 ( .ip1(n10257), .ip2(n10474), .op(n10254) );
  nand3_1 U12037 ( .ip1(n10256), .ip2(n10255), .ip3(n10254), .op(n2031) );
  nand2_1 U12038 ( .ip1(column[129]), .ip2(n10485), .op(n10260) );
  nand2_1 U12039 ( .ip1(\ROUTEDATA/regData [129]), .ip2(n10479), .op(n10259)
         );
  nand2_1 U12040 ( .ip1(n10257), .ip2(n10480), .op(n10258) );
  nand3_1 U12041 ( .ip1(n10260), .ip2(n10259), .ip3(n10258), .op(n2030) );
  nand2_1 U12042 ( .ip1(n10444), .ip2(column[145]), .op(n10262) );
  nand2_1 U12043 ( .ip1(n10262), .ip2(n10261), .op(n10263) );
  mux2_1 U12044 ( .ip1(n10263), .ip2(\ROUTEDATA/regData [145]), .s(n10488), 
        .op(n2029) );
  nand2_1 U12045 ( .ip1(n10485), .ip2(column[2]), .op(n10267) );
  nand2_1 U12046 ( .ip1(\ROUTEDATA/regData [2]), .ip2(n10432), .op(n10266) );
  nand2_1 U12047 ( .ip1(n10434), .ip2(n10264), .op(n10293) );
  inv_1 U12048 ( .ip(n10293), .op(n10289) );
  nand2_1 U12049 ( .ip1(n10289), .ip2(n10435), .op(n10265) );
  nand3_1 U12050 ( .ip1(n10267), .ip2(n10266), .ip3(n10265), .op(n2028) );
  nand2_1 U12051 ( .ip1(n10444), .ip2(column[18]), .op(n10270) );
  nand2_1 U12052 ( .ip1(\ROUTEDATA/regData [18]), .ip2(n10439), .op(n10269) );
  nand2_1 U12053 ( .ip1(n10289), .ip2(n10440), .op(n10268) );
  nand3_1 U12054 ( .ip1(n10270), .ip2(n10269), .ip3(n10268), .op(n2027) );
  nand2_1 U12055 ( .ip1(column[34]), .ip2(n10472), .op(n10273) );
  nand2_1 U12056 ( .ip1(n10289), .ip2(n10445), .op(n10272) );
  nand2_1 U12057 ( .ip1(\ROUTEDATA/regData [34]), .ip2(n10446), .op(n10271) );
  nand3_1 U12058 ( .ip1(n10273), .ip2(n10272), .ip3(n10271), .op(n2026) );
  nand2_1 U12059 ( .ip1(column[50]), .ip2(n10485), .op(n10276) );
  nand2_1 U12060 ( .ip1(\ROUTEDATA/regData [50]), .ip2(n10450), .op(n10275) );
  nand2_1 U12061 ( .ip1(n10289), .ip2(n10452), .op(n10274) );
  nand3_1 U12062 ( .ip1(n10276), .ip2(n10275), .ip3(n10274), .op(n2025) );
  nand2_1 U12063 ( .ip1(column[66]), .ip2(n10444), .op(n10279) );
  nand2_1 U12064 ( .ip1(n10289), .ip2(n10456), .op(n10278) );
  nand2_1 U12065 ( .ip1(\ROUTEDATA/regData [66]), .ip2(n10457), .op(n10277) );
  nand3_1 U12066 ( .ip1(n10279), .ip2(n10278), .ip3(n10277), .op(n2024) );
  nand2_1 U12067 ( .ip1(column[82]), .ip2(n10472), .op(n10282) );
  nand2_1 U12068 ( .ip1(n10289), .ip2(n10461), .op(n10281) );
  nand2_1 U12069 ( .ip1(\ROUTEDATA/regData [82]), .ip2(n10462), .op(n10280) );
  nand3_1 U12070 ( .ip1(n10282), .ip2(n10281), .ip3(n10280), .op(n2023) );
  nand2_1 U12071 ( .ip1(column[98]), .ip2(n10478), .op(n10285) );
  nand2_1 U12072 ( .ip1(n10289), .ip2(n10466), .op(n10284) );
  nand2_1 U12073 ( .ip1(\ROUTEDATA/regData [98]), .ip2(n10467), .op(n10283) );
  nand3_1 U12074 ( .ip1(n10285), .ip2(n10284), .ip3(n10283), .op(n2022) );
  nand2_1 U12075 ( .ip1(column[114]), .ip2(n10444), .op(n10288) );
  nand2_1 U12076 ( .ip1(n10289), .ip2(n10474), .op(n10287) );
  nand2_1 U12077 ( .ip1(\ROUTEDATA/regData [114]), .ip2(n10471), .op(n10286)
         );
  nand3_1 U12078 ( .ip1(n10288), .ip2(n10287), .ip3(n10286), .op(n2021) );
  nand2_1 U12079 ( .ip1(column[130]), .ip2(n10444), .op(n10292) );
  nand2_1 U12080 ( .ip1(n10289), .ip2(n10480), .op(n10291) );
  nand2_1 U12081 ( .ip1(\ROUTEDATA/regData [130]), .ip2(n10479), .op(n10290)
         );
  nand3_1 U12082 ( .ip1(n10292), .ip2(n10291), .ip3(n10290), .op(n2020) );
  nand2_1 U12083 ( .ip1(n10485), .ip2(column[146]), .op(n10294) );
  nand2_1 U12084 ( .ip1(n10294), .ip2(n10293), .op(n10295) );
  mux2_1 U12085 ( .ip1(n10295), .ip2(\ROUTEDATA/regData [146]), .s(n10488), 
        .op(n2019) );
  nand2_1 U12086 ( .ip1(n10485), .ip2(column[3]), .op(n10299) );
  nand2_1 U12087 ( .ip1(\ROUTEDATA/regData [3]), .ip2(n10432), .op(n10298) );
  nand2_1 U12088 ( .ip1(n10434), .ip2(n10296), .op(n10325) );
  inv_1 U12089 ( .ip(n10325), .op(n10321) );
  nand2_1 U12090 ( .ip1(n10321), .ip2(n10435), .op(n10297) );
  nand3_1 U12091 ( .ip1(n10299), .ip2(n10298), .ip3(n10297), .op(n2018) );
  nand2_1 U12092 ( .ip1(n10444), .ip2(column[19]), .op(n10302) );
  nand2_1 U12093 ( .ip1(\ROUTEDATA/regData [19]), .ip2(n10439), .op(n10301) );
  nand2_1 U12094 ( .ip1(n10321), .ip2(n10440), .op(n10300) );
  nand3_1 U12095 ( .ip1(n10302), .ip2(n10301), .ip3(n10300), .op(n2017) );
  nand2_1 U12096 ( .ip1(column[35]), .ip2(n10472), .op(n10305) );
  nand2_1 U12097 ( .ip1(n10321), .ip2(n10445), .op(n10304) );
  nand2_1 U12098 ( .ip1(\ROUTEDATA/regData [35]), .ip2(n10446), .op(n10303) );
  nand3_1 U12099 ( .ip1(n10305), .ip2(n10304), .ip3(n10303), .op(n2016) );
  nand2_1 U12100 ( .ip1(column[51]), .ip2(n10485), .op(n10308) );
  nand2_1 U12101 ( .ip1(\ROUTEDATA/regData [51]), .ip2(n10450), .op(n10307) );
  nand2_1 U12102 ( .ip1(n10321), .ip2(n10452), .op(n10306) );
  nand3_1 U12103 ( .ip1(n10308), .ip2(n10307), .ip3(n10306), .op(n2015) );
  nand2_1 U12104 ( .ip1(column[67]), .ip2(n10485), .op(n10311) );
  nand2_1 U12105 ( .ip1(n10321), .ip2(n10456), .op(n10310) );
  nand2_1 U12106 ( .ip1(\ROUTEDATA/regData [67]), .ip2(n10457), .op(n10309) );
  nand3_1 U12107 ( .ip1(n10311), .ip2(n10310), .ip3(n10309), .op(n2014) );
  nand2_1 U12108 ( .ip1(column[83]), .ip2(n10485), .op(n10314) );
  nand2_1 U12109 ( .ip1(\ROUTEDATA/regData [83]), .ip2(n10462), .op(n10313) );
  nand2_1 U12110 ( .ip1(n10321), .ip2(n10461), .op(n10312) );
  nand3_1 U12111 ( .ip1(n10314), .ip2(n10313), .ip3(n10312), .op(n2013) );
  nand2_1 U12112 ( .ip1(column[99]), .ip2(n10444), .op(n10317) );
  nand2_1 U12113 ( .ip1(n10321), .ip2(n10466), .op(n10316) );
  nand2_1 U12114 ( .ip1(\ROUTEDATA/regData [99]), .ip2(n10467), .op(n10315) );
  nand3_1 U12115 ( .ip1(n10317), .ip2(n10316), .ip3(n10315), .op(n2012) );
  nand2_1 U12116 ( .ip1(column[115]), .ip2(n10478), .op(n10320) );
  nand2_1 U12117 ( .ip1(n10321), .ip2(n10474), .op(n10319) );
  nand2_1 U12118 ( .ip1(\ROUTEDATA/regData [115]), .ip2(n10471), .op(n10318)
         );
  nand3_1 U12119 ( .ip1(n10320), .ip2(n10319), .ip3(n10318), .op(n2011) );
  nand2_1 U12120 ( .ip1(column[131]), .ip2(n10444), .op(n10324) );
  nand2_1 U12121 ( .ip1(n10321), .ip2(n10480), .op(n10323) );
  nand2_1 U12122 ( .ip1(\ROUTEDATA/regData [131]), .ip2(n10479), .op(n10322)
         );
  nand3_1 U12123 ( .ip1(n10324), .ip2(n10323), .ip3(n10322), .op(n2010) );
  nand2_1 U12124 ( .ip1(n10485), .ip2(column[147]), .op(n10326) );
  nand2_1 U12125 ( .ip1(n10326), .ip2(n10325), .op(n10327) );
  mux2_1 U12126 ( .ip1(n10327), .ip2(\ROUTEDATA/regData [147]), .s(n10488), 
        .op(n2009) );
  nand2_1 U12127 ( .ip1(n10472), .ip2(column[4]), .op(n10331) );
  nand2_1 U12128 ( .ip1(\ROUTEDATA/regData [4]), .ip2(n10432), .op(n10330) );
  and2_1 U12129 ( .ip1(n10434), .ip2(n10328), .op(n10356) );
  nand2_1 U12130 ( .ip1(n10356), .ip2(n10435), .op(n10329) );
  nand3_1 U12131 ( .ip1(n10331), .ip2(n10330), .ip3(n10329), .op(n2008) );
  nand2_1 U12132 ( .ip1(column[20]), .ip2(n10478), .op(n10334) );
  nand2_1 U12133 ( .ip1(\ROUTEDATA/regData [20]), .ip2(n10439), .op(n10333) );
  nand2_1 U12134 ( .ip1(n10356), .ip2(n10440), .op(n10332) );
  nand3_1 U12135 ( .ip1(n10334), .ip2(n10333), .ip3(n10332), .op(n2007) );
  nand2_1 U12136 ( .ip1(column[36]), .ip2(n10478), .op(n10337) );
  nand2_1 U12137 ( .ip1(\ROUTEDATA/regData [36]), .ip2(n10446), .op(n10336) );
  nand2_1 U12138 ( .ip1(n10356), .ip2(n10445), .op(n10335) );
  nand3_1 U12139 ( .ip1(n10337), .ip2(n10336), .ip3(n10335), .op(n2006) );
  nand2_1 U12140 ( .ip1(column[52]), .ip2(n10478), .op(n10340) );
  nand2_1 U12141 ( .ip1(n10356), .ip2(n10452), .op(n10339) );
  nand2_1 U12142 ( .ip1(\ROUTEDATA/regData [52]), .ip2(n10450), .op(n10338) );
  nand3_1 U12143 ( .ip1(n10340), .ip2(n10339), .ip3(n10338), .op(n2005) );
  nand2_1 U12144 ( .ip1(column[68]), .ip2(n10444), .op(n10343) );
  nand2_1 U12145 ( .ip1(n10356), .ip2(n10456), .op(n10342) );
  nand2_1 U12146 ( .ip1(\ROUTEDATA/regData [68]), .ip2(n10457), .op(n10341) );
  nand3_1 U12147 ( .ip1(n10343), .ip2(n10342), .ip3(n10341), .op(n2004) );
  nand2_1 U12148 ( .ip1(column[84]), .ip2(n10478), .op(n10346) );
  nand2_1 U12149 ( .ip1(\ROUTEDATA/regData [84]), .ip2(n10462), .op(n10345) );
  nand2_1 U12150 ( .ip1(n10356), .ip2(n10461), .op(n10344) );
  nand3_1 U12151 ( .ip1(n10346), .ip2(n10345), .ip3(n10344), .op(n2003) );
  nand2_1 U12152 ( .ip1(column[100]), .ip2(n10485), .op(n10349) );
  nand2_1 U12153 ( .ip1(n10356), .ip2(n10466), .op(n10348) );
  nand2_1 U12154 ( .ip1(\ROUTEDATA/regData [100]), .ip2(n10467), .op(n10347)
         );
  nand3_1 U12155 ( .ip1(n10349), .ip2(n10348), .ip3(n10347), .op(n2002) );
  nand2_1 U12156 ( .ip1(column[116]), .ip2(n10485), .op(n10352) );
  nand2_1 U12157 ( .ip1(\ROUTEDATA/regData [116]), .ip2(n10471), .op(n10351)
         );
  nand2_1 U12158 ( .ip1(n10356), .ip2(n10474), .op(n10350) );
  nand3_1 U12159 ( .ip1(n10352), .ip2(n10351), .ip3(n10350), .op(n2001) );
  nand2_1 U12160 ( .ip1(column[132]), .ip2(n10444), .op(n10355) );
  nand2_1 U12161 ( .ip1(\ROUTEDATA/regData [132]), .ip2(n10479), .op(n10354)
         );
  nand2_1 U12162 ( .ip1(n10356), .ip2(n10480), .op(n10353) );
  nand3_1 U12163 ( .ip1(n10355), .ip2(n10354), .ip3(n10353), .op(n2000) );
  inv_1 U12164 ( .ip(n10488), .op(n10428) );
  nand2_1 U12165 ( .ip1(n10428), .ip2(n10356), .op(n10359) );
  nand2_1 U12166 ( .ip1(n10485), .ip2(column[148]), .op(n10358) );
  nand2_1 U12167 ( .ip1(n10488), .ip2(\ROUTEDATA/regData [148]), .op(n10357)
         );
  nand3_1 U12168 ( .ip1(n10359), .ip2(n10358), .ip3(n10357), .op(n1999) );
  nand2_1 U12169 ( .ip1(column[5]), .ip2(n10444), .op(n10363) );
  and2_1 U12170 ( .ip1(n10434), .ip2(n10360), .op(n10390) );
  nand2_1 U12171 ( .ip1(n10390), .ip2(n10435), .op(n10362) );
  nand2_1 U12172 ( .ip1(\ROUTEDATA/regData [5]), .ip2(n10432), .op(n10361) );
  nand3_1 U12173 ( .ip1(n10363), .ip2(n10362), .ip3(n10361), .op(n1998) );
  nand2_1 U12174 ( .ip1(column[21]), .ip2(n10472), .op(n10366) );
  nand2_1 U12175 ( .ip1(\ROUTEDATA/regData [21]), .ip2(n10439), .op(n10365) );
  nand2_1 U12176 ( .ip1(n10390), .ip2(n10440), .op(n10364) );
  nand3_1 U12177 ( .ip1(n10366), .ip2(n10365), .ip3(n10364), .op(n1997) );
  nand2_1 U12178 ( .ip1(column[37]), .ip2(n10478), .op(n10369) );
  nand2_1 U12179 ( .ip1(n10390), .ip2(n10445), .op(n10368) );
  nand2_1 U12180 ( .ip1(\ROUTEDATA/regData [37]), .ip2(n10446), .op(n10367) );
  nand3_1 U12181 ( .ip1(n10369), .ip2(n10368), .ip3(n10367), .op(n1996) );
  nand2_1 U12182 ( .ip1(column[53]), .ip2(n10485), .op(n10372) );
  nand2_1 U12183 ( .ip1(n10390), .ip2(n10452), .op(n10371) );
  nand2_1 U12184 ( .ip1(\ROUTEDATA/regData [53]), .ip2(n10450), .op(n10370) );
  nand3_1 U12185 ( .ip1(n10372), .ip2(n10371), .ip3(n10370), .op(n1995) );
  nand2_1 U12186 ( .ip1(\ROUTEDATA/regData [69]), .ip2(n10457), .op(n10377) );
  or2_1 U12187 ( .ip1(n10444), .ip2(n10390), .op(n10374) );
  or2_1 U12188 ( .ip1(column[69]), .ip2(n10390), .op(n10373) );
  nand2_1 U12189 ( .ip1(n10374), .ip2(n10373), .op(n10375) );
  or2_1 U12190 ( .ip1(n10412), .ip2(n10375), .op(n10376) );
  nand2_1 U12191 ( .ip1(n10377), .ip2(n10376), .op(n1994) );
  nand2_1 U12192 ( .ip1(column[85]), .ip2(n10444), .op(n10380) );
  nand2_1 U12193 ( .ip1(n10390), .ip2(n10461), .op(n10379) );
  nand2_1 U12194 ( .ip1(\ROUTEDATA/regData [85]), .ip2(n10462), .op(n10378) );
  nand3_1 U12195 ( .ip1(n10380), .ip2(n10379), .ip3(n10378), .op(n1993) );
  nand2_1 U12196 ( .ip1(column[101]), .ip2(n10485), .op(n10383) );
  nand2_1 U12197 ( .ip1(\ROUTEDATA/regData [101]), .ip2(n10467), .op(n10382)
         );
  nand2_1 U12198 ( .ip1(n10390), .ip2(n10466), .op(n10381) );
  nand3_1 U12199 ( .ip1(n10383), .ip2(n10382), .ip3(n10381), .op(n1992) );
  nand2_1 U12200 ( .ip1(column[117]), .ip2(n10444), .op(n10386) );
  nand2_1 U12201 ( .ip1(\ROUTEDATA/regData [117]), .ip2(n10471), .op(n10385)
         );
  nand2_1 U12202 ( .ip1(n10390), .ip2(n10474), .op(n10384) );
  nand3_1 U12203 ( .ip1(n10386), .ip2(n10385), .ip3(n10384), .op(n1991) );
  nand2_1 U12204 ( .ip1(column[133]), .ip2(n10472), .op(n10389) );
  nand2_1 U12205 ( .ip1(n10390), .ip2(n10480), .op(n10388) );
  nand2_1 U12206 ( .ip1(\ROUTEDATA/regData [133]), .ip2(n10479), .op(n10387)
         );
  nand3_1 U12207 ( .ip1(n10389), .ip2(n10388), .ip3(n10387), .op(n1990) );
  nand2_1 U12208 ( .ip1(n10428), .ip2(n10390), .op(n10393) );
  nand2_1 U12209 ( .ip1(n10444), .ip2(column[149]), .op(n10392) );
  nand2_1 U12210 ( .ip1(n10488), .ip2(\ROUTEDATA/regData [149]), .op(n10391)
         );
  nand3_1 U12211 ( .ip1(n10393), .ip2(n10392), .ip3(n10391), .op(n1989) );
  nand2_1 U12212 ( .ip1(column[6]), .ip2(n10472), .op(n10397) );
  nand2_1 U12213 ( .ip1(\ROUTEDATA/regData [6]), .ip2(n10432), .op(n10396) );
  nand2_1 U12214 ( .ip1(n10394), .ip2(n10434), .op(n10401) );
  inv_1 U12215 ( .ip(n10401), .op(n10427) );
  nand2_1 U12216 ( .ip1(n10427), .ip2(n10435), .op(n10395) );
  nand3_1 U12217 ( .ip1(n10397), .ip2(n10396), .ip3(n10395), .op(n1988) );
  nand2_1 U12218 ( .ip1(column[22]), .ip2(n10444), .op(n10400) );
  nand2_1 U12219 ( .ip1(\ROUTEDATA/regData [22]), .ip2(n10439), .op(n10399) );
  nand2_1 U12220 ( .ip1(n10427), .ip2(n10440), .op(n10398) );
  nand3_1 U12221 ( .ip1(n10400), .ip2(n10399), .ip3(n10398), .op(n1987) );
  nand2_1 U12222 ( .ip1(\ROUTEDATA/regData [38]), .ip2(n10446), .op(n10405) );
  nand2_1 U12223 ( .ip1(n10472), .ip2(column[38]), .op(n10402) );
  nand2_1 U12224 ( .ip1(n10402), .ip2(n10401), .op(n10403) );
  nand2_1 U12225 ( .ip1(n10403), .ip2(n10445), .op(n10404) );
  nand2_1 U12226 ( .ip1(n10405), .ip2(n10404), .op(n1986) );
  nand2_1 U12227 ( .ip1(column[54]), .ip2(n10444), .op(n10408) );
  nand2_1 U12228 ( .ip1(\ROUTEDATA/regData [54]), .ip2(n10450), .op(n10407) );
  nand2_1 U12229 ( .ip1(n10427), .ip2(n10452), .op(n10406) );
  nand3_1 U12230 ( .ip1(n10408), .ip2(n10407), .ip3(n10406), .op(n1985) );
  nand2_1 U12231 ( .ip1(\ROUTEDATA/regData [70]), .ip2(n10457), .op(n10414) );
  or2_1 U12232 ( .ip1(n10444), .ip2(n10427), .op(n10410) );
  or2_1 U12233 ( .ip1(column[70]), .ip2(n10427), .op(n10409) );
  nand2_1 U12234 ( .ip1(n10410), .ip2(n10409), .op(n10411) );
  or2_1 U12235 ( .ip1(n10412), .ip2(n10411), .op(n10413) );
  nand2_1 U12236 ( .ip1(n10414), .ip2(n10413), .op(n1984) );
  nand2_1 U12237 ( .ip1(column[86]), .ip2(n10444), .op(n10417) );
  nand2_1 U12238 ( .ip1(n10427), .ip2(n10461), .op(n10416) );
  nand2_1 U12239 ( .ip1(\ROUTEDATA/regData [86]), .ip2(n10462), .op(n10415) );
  nand3_1 U12240 ( .ip1(n10417), .ip2(n10416), .ip3(n10415), .op(n1983) );
  nand2_1 U12241 ( .ip1(column[102]), .ip2(n10472), .op(n10420) );
  nand2_1 U12242 ( .ip1(n10427), .ip2(n10466), .op(n10419) );
  nand2_1 U12243 ( .ip1(\ROUTEDATA/regData [102]), .ip2(n10467), .op(n10418)
         );
  nand3_1 U12244 ( .ip1(n10420), .ip2(n10419), .ip3(n10418), .op(n1982) );
  nand2_1 U12245 ( .ip1(column[118]), .ip2(n10472), .op(n10423) );
  nand2_1 U12246 ( .ip1(n10427), .ip2(n10474), .op(n10422) );
  nand2_1 U12247 ( .ip1(\ROUTEDATA/regData [118]), .ip2(n10471), .op(n10421)
         );
  nand3_1 U12248 ( .ip1(n10423), .ip2(n10422), .ip3(n10421), .op(n1981) );
  nand2_1 U12249 ( .ip1(column[134]), .ip2(n10472), .op(n10426) );
  nand2_1 U12250 ( .ip1(\ROUTEDATA/regData [134]), .ip2(n10479), .op(n10425)
         );
  nand2_1 U12251 ( .ip1(n10427), .ip2(n10480), .op(n10424) );
  nand3_1 U12252 ( .ip1(n10426), .ip2(n10425), .ip3(n10424), .op(n1980) );
  nand2_1 U12253 ( .ip1(n10428), .ip2(n10427), .op(n10431) );
  nand2_1 U12254 ( .ip1(n10444), .ip2(column[150]), .op(n10430) );
  nand2_1 U12255 ( .ip1(n10488), .ip2(\ROUTEDATA/regData [150]), .op(n10429)
         );
  nand3_1 U12256 ( .ip1(n10431), .ip2(n10430), .ip3(n10429), .op(n1979) );
  nand2_1 U12257 ( .ip1(column[7]), .ip2(n10444), .op(n10438) );
  nand2_1 U12258 ( .ip1(\ROUTEDATA/regData [7]), .ip2(n10432), .op(n10437) );
  nand2_1 U12259 ( .ip1(n10434), .ip2(n10433), .op(n10486) );
  inv_1 U12260 ( .ip(n10486), .op(n10481) );
  nand2_1 U12261 ( .ip1(n10481), .ip2(n10435), .op(n10436) );
  nand3_1 U12262 ( .ip1(n10438), .ip2(n10437), .ip3(n10436), .op(n1978) );
  nand2_1 U12263 ( .ip1(column[23]), .ip2(n10444), .op(n10443) );
  nand2_1 U12264 ( .ip1(\ROUTEDATA/regData [23]), .ip2(n10439), .op(n10442) );
  nand2_1 U12265 ( .ip1(n10481), .ip2(n10440), .op(n10441) );
  nand3_1 U12266 ( .ip1(n10443), .ip2(n10442), .ip3(n10441), .op(n1977) );
  nand2_1 U12267 ( .ip1(column[39]), .ip2(n10444), .op(n10449) );
  nand2_1 U12268 ( .ip1(n10481), .ip2(n10445), .op(n10448) );
  nand2_1 U12269 ( .ip1(\ROUTEDATA/regData [39]), .ip2(n10446), .op(n10447) );
  nand3_1 U12270 ( .ip1(n10449), .ip2(n10448), .ip3(n10447), .op(n1976) );
  nand2_1 U12271 ( .ip1(\ROUTEDATA/regData [55]), .ip2(n10450), .op(n10455) );
  nand2_1 U12272 ( .ip1(n10472), .ip2(column[55]), .op(n10451) );
  nand2_1 U12273 ( .ip1(n10451), .ip2(n10486), .op(n10453) );
  nand2_1 U12274 ( .ip1(n10453), .ip2(n10452), .op(n10454) );
  nand2_1 U12275 ( .ip1(n10455), .ip2(n10454), .op(n1975) );
  nand2_1 U12276 ( .ip1(column[71]), .ip2(n10472), .op(n10460) );
  nand2_1 U12277 ( .ip1(n10481), .ip2(n10456), .op(n10459) );
  nand2_1 U12278 ( .ip1(\ROUTEDATA/regData [71]), .ip2(n10457), .op(n10458) );
  nand3_1 U12279 ( .ip1(n10460), .ip2(n10459), .ip3(n10458), .op(n1974) );
  nand2_1 U12280 ( .ip1(column[87]), .ip2(n10478), .op(n10465) );
  nand2_1 U12281 ( .ip1(n10481), .ip2(n10461), .op(n10464) );
  nand2_1 U12282 ( .ip1(\ROUTEDATA/regData [87]), .ip2(n10462), .op(n10463) );
  nand3_1 U12283 ( .ip1(n10465), .ip2(n10464), .ip3(n10463), .op(n1973) );
  nand2_1 U12284 ( .ip1(column[103]), .ip2(n10472), .op(n10470) );
  nand2_1 U12285 ( .ip1(n10481), .ip2(n10466), .op(n10469) );
  nand2_1 U12286 ( .ip1(\ROUTEDATA/regData [103]), .ip2(n10467), .op(n10468)
         );
  nand3_1 U12287 ( .ip1(n10470), .ip2(n10469), .ip3(n10468), .op(n1972) );
  nand2_1 U12288 ( .ip1(\ROUTEDATA/regData [119]), .ip2(n10471), .op(n10477)
         );
  nand2_1 U12289 ( .ip1(n10472), .ip2(column[119]), .op(n10473) );
  nand2_1 U12290 ( .ip1(n10473), .ip2(n10486), .op(n10475) );
  nand2_1 U12291 ( .ip1(n10475), .ip2(n10474), .op(n10476) );
  nand2_1 U12292 ( .ip1(n10477), .ip2(n10476), .op(n1971) );
  nand2_1 U12293 ( .ip1(column[135]), .ip2(n10478), .op(n10484) );
  nand2_1 U12294 ( .ip1(\ROUTEDATA/regData [135]), .ip2(n10479), .op(n10483)
         );
  nand2_1 U12295 ( .ip1(n10481), .ip2(n10480), .op(n10482) );
  nand3_1 U12296 ( .ip1(n10484), .ip2(n10483), .ip3(n10482), .op(n1970) );
  nand2_1 U12297 ( .ip1(n10485), .ip2(column[151]), .op(n10487) );
  nand2_1 U12298 ( .ip1(n10487), .ip2(n10486), .op(n10489) );
  mux2_1 U12299 ( .ip1(n10489), .ip2(\ROUTEDATA/regData [151]), .s(n10488), 
        .op(n1969) );
  mux2_1 U12300 ( .ip1(\ANSWER/mem[0][2][0] ), .ip2(\ANSWER/mem[1][2][0] ), 
        .s(n11506), .op(n10491) );
  mux2_1 U12301 ( .ip1(\ANSWER/mem[2][2][0] ), .ip2(\ANSWER/mem[3][2][0] ), 
        .s(n8833), .op(n10490) );
  mux2_1 U12302 ( .ip1(n10491), .ip2(n10490), .s(n11868), .op(n10495) );
  mux2_1 U12303 ( .ip1(\ANSWER/mem[4][2][0] ), .ip2(\ANSWER/mem[5][2][0] ), 
        .s(n10583), .op(n10493) );
  inv_1 U12304 ( .ip(n12109), .op(n10588) );
  buf_1 U12305 ( .ip(n10588), .op(n10583) );
  mux2_1 U12306 ( .ip1(\ANSWER/mem[6][2][0] ), .ip2(\ANSWER/mem[7][2][0] ), 
        .s(n10583), .op(n10492) );
  mux2_1 U12307 ( .ip1(n10493), .ip2(n10492), .s(n11976), .op(n10494) );
  mux2_1 U12308 ( .ip1(n10495), .ip2(n10494), .s(n11454), .op(n10497) );
  mux2_1 U12309 ( .ip1(\ANSWER/mem[8][2][0] ), .ip2(\ANSWER/mem[9][2][0] ), 
        .s(n10583), .op(n10496) );
  mux2_1 U12310 ( .ip1(n10497), .ip2(n10496), .s(n11336), .op(n10498) );
  nand2_1 U12311 ( .ip1(n12147), .ip2(n10498), .op(n10570) );
  mux2_1 U12312 ( .ip1(\ANSWER/mem[0][1][0] ), .ip2(\ANSWER/mem[1][1][0] ), 
        .s(n12085), .op(n10500) );
  mux2_1 U12313 ( .ip1(\ANSWER/mem[2][1][0] ), .ip2(\ANSWER/mem[3][1][0] ), 
        .s(n11546), .op(n10499) );
  mux2_1 U12314 ( .ip1(n10500), .ip2(n10499), .s(n11868), .op(n10504) );
  mux2_1 U12315 ( .ip1(\ANSWER/mem[4][1][0] ), .ip2(\ANSWER/mem[5][1][0] ), 
        .s(n10816), .op(n10502) );
  mux2_1 U12316 ( .ip1(\ANSWER/mem[6][1][0] ), .ip2(\ANSWER/mem[7][1][0] ), 
        .s(n11070), .op(n10501) );
  mux2_1 U12317 ( .ip1(n10502), .ip2(n10501), .s(n11976), .op(n10503) );
  mux2_1 U12318 ( .ip1(n10504), .ip2(n10503), .s(n11454), .op(n10506) );
  mux2_1 U12319 ( .ip1(\ANSWER/mem[8][1][0] ), .ip2(\ANSWER/mem[9][1][0] ), 
        .s(n11070), .op(n10505) );
  mux2_1 U12320 ( .ip1(n10506), .ip2(n10505), .s(n11336), .op(n10558) );
  mux2_1 U12321 ( .ip1(\ANSWER/mem[0][3][0] ), .ip2(\ANSWER/mem[1][3][0] ), 
        .s(n10583), .op(n10508) );
  mux2_1 U12322 ( .ip1(\ANSWER/mem[2][3][0] ), .ip2(\ANSWER/mem[3][3][0] ), 
        .s(n10583), .op(n10507) );
  mux2_1 U12323 ( .ip1(n10508), .ip2(n10507), .s(n11008), .op(n10512) );
  mux2_1 U12324 ( .ip1(\ANSWER/mem[4][3][0] ), .ip2(\ANSWER/mem[5][3][0] ), 
        .s(n10583), .op(n10510) );
  mux2_1 U12325 ( .ip1(\ANSWER/mem[6][3][0] ), .ip2(\ANSWER/mem[7][3][0] ), 
        .s(n10583), .op(n10509) );
  mux2_1 U12326 ( .ip1(n10510), .ip2(n10509), .s(n11224), .op(n10511) );
  mux2_1 U12327 ( .ip1(n10512), .ip2(n10511), .s(n11454), .op(n10514) );
  mux2_1 U12328 ( .ip1(\ANSWER/mem[8][3][0] ), .ip2(\ANSWER/mem[9][3][0] ), 
        .s(n10583), .op(n10513) );
  mux2_1 U12329 ( .ip1(n10514), .ip2(n10513), .s(n11336), .op(n10515) );
  and2_1 U12330 ( .ip1(n12137), .ip2(n10515), .op(n10557) );
  mux2_1 U12331 ( .ip1(\ANSWER/mem[0][5][0] ), .ip2(\ANSWER/mem[1][5][0] ), 
        .s(n10583), .op(n10517) );
  mux2_1 U12332 ( .ip1(\ANSWER/mem[2][5][0] ), .ip2(\ANSWER/mem[3][5][0] ), 
        .s(n10588), .op(n10516) );
  mux2_1 U12333 ( .ip1(n10517), .ip2(n10516), .s(n11868), .op(n10521) );
  mux2_1 U12334 ( .ip1(\ANSWER/mem[4][5][0] ), .ip2(\ANSWER/mem[5][5][0] ), 
        .s(n10588), .op(n10519) );
  mux2_1 U12335 ( .ip1(\ANSWER/mem[6][5][0] ), .ip2(\ANSWER/mem[7][5][0] ), 
        .s(n10588), .op(n10518) );
  mux2_1 U12336 ( .ip1(n10519), .ip2(n10518), .s(n11976), .op(n10520) );
  mux2_1 U12337 ( .ip1(n10521), .ip2(n10520), .s(n11454), .op(n10523) );
  mux2_1 U12338 ( .ip1(\ANSWER/mem[8][5][0] ), .ip2(\ANSWER/mem[9][5][0] ), 
        .s(n10588), .op(n10522) );
  mux2_1 U12339 ( .ip1(n10523), .ip2(n10522), .s(n11336), .op(n10524) );
  nand2_1 U12340 ( .ip1(n12127), .ip2(n10524), .op(n10555) );
  mux2_1 U12341 ( .ip1(\ANSWER/mem[0][7][0] ), .ip2(\ANSWER/mem[1][7][0] ), 
        .s(n10588), .op(n10526) );
  mux2_1 U12342 ( .ip1(\ANSWER/mem[2][7][0] ), .ip2(\ANSWER/mem[3][7][0] ), 
        .s(n10588), .op(n10525) );
  mux2_1 U12343 ( .ip1(n10526), .ip2(n10525), .s(n11008), .op(n10530) );
  mux2_1 U12344 ( .ip1(\ANSWER/mem[4][7][0] ), .ip2(\ANSWER/mem[5][7][0] ), 
        .s(n10588), .op(n10528) );
  mux2_1 U12345 ( .ip1(\ANSWER/mem[6][7][0] ), .ip2(\ANSWER/mem[7][7][0] ), 
        .s(n10588), .op(n10527) );
  mux2_1 U12346 ( .ip1(n10528), .ip2(n10527), .s(n11868), .op(n10529) );
  mux2_1 U12347 ( .ip1(n10530), .ip2(n10529), .s(n11454), .op(n10532) );
  mux2_1 U12348 ( .ip1(\ANSWER/mem[8][7][0] ), .ip2(\ANSWER/mem[9][7][0] ), 
        .s(n10583), .op(n10531) );
  mux2_1 U12349 ( .ip1(n10532), .ip2(n10531), .s(n11336), .op(n10533) );
  nand2_1 U12350 ( .ip1(n12186), .ip2(n10533), .op(n10554) );
  mux2_1 U12351 ( .ip1(\ANSWER/mem[0][0][0] ), .ip2(\ANSWER/mem[1][0][0] ), 
        .s(n11164), .op(n10535) );
  mux2_1 U12352 ( .ip1(\ANSWER/mem[2][0][0] ), .ip2(\ANSWER/mem[3][0][0] ), 
        .s(n11437), .op(n10534) );
  mux2_1 U12353 ( .ip1(n10535), .ip2(n10534), .s(n11008), .op(n10539) );
  mux2_1 U12354 ( .ip1(\ANSWER/mem[4][0][0] ), .ip2(\ANSWER/mem[5][0][0] ), 
        .s(n11070), .op(n10537) );
  mux2_1 U12355 ( .ip1(\ANSWER/mem[6][0][0] ), .ip2(\ANSWER/mem[7][0][0] ), 
        .s(n11758), .op(n10536) );
  mux2_1 U12356 ( .ip1(n10537), .ip2(n10536), .s(n11868), .op(n10538) );
  mux2_1 U12357 ( .ip1(n10539), .ip2(n10538), .s(n11454), .op(n10541) );
  mux2_1 U12358 ( .ip1(\ANSWER/mem[8][0][0] ), .ip2(\ANSWER/mem[9][0][0] ), 
        .s(n11164), .op(n10540) );
  mux2_1 U12359 ( .ip1(n10541), .ip2(n10540), .s(n11336), .op(n10542) );
  nand2_1 U12360 ( .ip1(n12108), .ip2(n10542), .op(n10553) );
  mux2_1 U12361 ( .ip1(\ANSWER/mem[0][4][0] ), .ip2(\ANSWER/mem[1][4][0] ), 
        .s(n10583), .op(n10544) );
  mux2_1 U12362 ( .ip1(\ANSWER/mem[2][4][0] ), .ip2(\ANSWER/mem[3][4][0] ), 
        .s(n10583), .op(n10543) );
  mux2_1 U12363 ( .ip1(n10544), .ip2(n10543), .s(n11868), .op(n10548) );
  mux2_1 U12364 ( .ip1(\ANSWER/mem[4][4][0] ), .ip2(\ANSWER/mem[5][4][0] ), 
        .s(n10583), .op(n10546) );
  mux2_1 U12365 ( .ip1(\ANSWER/mem[6][4][0] ), .ip2(\ANSWER/mem[7][4][0] ), 
        .s(n10583), .op(n10545) );
  mux2_1 U12366 ( .ip1(n10546), .ip2(n10545), .s(n11224), .op(n10547) );
  mux2_1 U12367 ( .ip1(n10548), .ip2(n10547), .s(n11454), .op(n10550) );
  mux2_1 U12368 ( .ip1(\ANSWER/mem[8][4][0] ), .ip2(\ANSWER/mem[9][4][0] ), 
        .s(n10583), .op(n10549) );
  inv_1 U12369 ( .ip(n11996), .op(n11552) );
  mux2_1 U12370 ( .ip1(n10550), .ip2(n10549), .s(n11552), .op(n10551) );
  nand2_1 U12371 ( .ip1(n12176), .ip2(n10551), .op(n10552) );
  nand4_1 U12372 ( .ip1(n10555), .ip2(n10554), .ip3(n10553), .ip4(n10552), 
        .op(n10556) );
  not_ab_or_c_or_d U12373 ( .ip1(n10558), .ip2(n12157), .ip3(n10557), .ip4(
        n10556), .op(n10569) );
  mux2_1 U12374 ( .ip1(\ANSWER/mem[0][6][0] ), .ip2(\ANSWER/mem[1][6][0] ), 
        .s(n10588), .op(n10560) );
  mux2_1 U12375 ( .ip1(\ANSWER/mem[2][6][0] ), .ip2(\ANSWER/mem[3][6][0] ), 
        .s(n10588), .op(n10559) );
  mux2_1 U12376 ( .ip1(n10560), .ip2(n10559), .s(n11224), .op(n10564) );
  mux2_1 U12377 ( .ip1(\ANSWER/mem[4][6][0] ), .ip2(\ANSWER/mem[5][6][0] ), 
        .s(n10588), .op(n10562) );
  mux2_1 U12378 ( .ip1(\ANSWER/mem[6][6][0] ), .ip2(\ANSWER/mem[7][6][0] ), 
        .s(n10588), .op(n10561) );
  mux2_1 U12379 ( .ip1(n10562), .ip2(n10561), .s(n11976), .op(n10563) );
  mux2_1 U12380 ( .ip1(n10564), .ip2(n10563), .s(n11454), .op(n10566) );
  mux2_1 U12381 ( .ip1(\ANSWER/mem[8][6][0] ), .ip2(\ANSWER/mem[9][6][0] ), 
        .s(n10588), .op(n10565) );
  mux2_1 U12382 ( .ip1(n10566), .ip2(n10565), .s(n11336), .op(n10567) );
  nand2_1 U12383 ( .ip1(n12168), .ip2(n10567), .op(n10568) );
  nand3_1 U12384 ( .ip1(n10570), .ip2(n10569), .ip3(n10568), .op(n10571) );
  nand2_1 U12385 ( .ip1(n10571), .ip2(n12190), .op(n10594) );
  mux2_1 U12386 ( .ip1(\ANSWER/mem[0][8][0] ), .ip2(\ANSWER/mem[1][8][0] ), 
        .s(n10583), .op(n10573) );
  mux2_1 U12387 ( .ip1(\ANSWER/mem[2][8][0] ), .ip2(\ANSWER/mem[3][8][0] ), 
        .s(n10588), .op(n10572) );
  mux2_1 U12388 ( .ip1(n10573), .ip2(n10572), .s(n11976), .op(n10577) );
  mux2_1 U12389 ( .ip1(\ANSWER/mem[4][8][0] ), .ip2(\ANSWER/mem[5][8][0] ), 
        .s(n10588), .op(n10575) );
  mux2_1 U12390 ( .ip1(\ANSWER/mem[6][8][0] ), .ip2(\ANSWER/mem[7][8][0] ), 
        .s(n10588), .op(n10574) );
  mux2_1 U12391 ( .ip1(n10575), .ip2(n10574), .s(n11868), .op(n10576) );
  mux2_1 U12392 ( .ip1(n10577), .ip2(n10576), .s(n11454), .op(n10579) );
  mux2_1 U12393 ( .ip1(\ANSWER/mem[8][8][0] ), .ip2(\ANSWER/mem[9][8][0] ), 
        .s(n10588), .op(n10578) );
  mux2_1 U12394 ( .ip1(n10579), .ip2(n10578), .s(n11336), .op(n10580) );
  nand2_1 U12395 ( .ip1(n12201), .ip2(n10580), .op(n10593) );
  mux2_1 U12396 ( .ip1(\ANSWER/mem[0][9][0] ), .ip2(\ANSWER/mem[1][9][0] ), 
        .s(n10588), .op(n10582) );
  mux2_1 U12397 ( .ip1(\ANSWER/mem[2][9][0] ), .ip2(\ANSWER/mem[3][9][0] ), 
        .s(n10588), .op(n10581) );
  mux2_1 U12398 ( .ip1(n10582), .ip2(n10581), .s(n11224), .op(n10587) );
  mux2_1 U12399 ( .ip1(\ANSWER/mem[4][9][0] ), .ip2(\ANSWER/mem[5][9][0] ), 
        .s(n10583), .op(n10585) );
  mux2_1 U12400 ( .ip1(\ANSWER/mem[6][9][0] ), .ip2(\ANSWER/mem[7][9][0] ), 
        .s(n10588), .op(n10584) );
  mux2_1 U12401 ( .ip1(n10585), .ip2(n10584), .s(n11976), .op(n10586) );
  mux2_1 U12402 ( .ip1(n10587), .ip2(n10586), .s(n11454), .op(n10590) );
  mux2_1 U12403 ( .ip1(\ANSWER/mem[8][9][0] ), .ip2(\ANSWER/mem[9][9][0] ), 
        .s(n10588), .op(n10589) );
  mux2_1 U12404 ( .ip1(n10590), .ip2(n10589), .s(n11336), .op(n10591) );
  nand2_1 U12405 ( .ip1(n12215), .ip2(n10591), .op(n10592) );
  nand3_1 U12406 ( .ip1(n10594), .ip2(n10593), .ip3(n10592), .op(\ANSWER/N487 ) );
  buf_1 U12407 ( .ip(n10878), .op(n10816) );
  mux2_1 U12408 ( .ip1(\ANSWER/mem[0][0][1] ), .ip2(\ANSWER/mem[1][0][1] ), 
        .s(n10816), .op(n10596) );
  mux2_1 U12409 ( .ip1(\ANSWER/mem[2][0][1] ), .ip2(\ANSWER/mem[3][0][1] ), 
        .s(n10816), .op(n10595) );
  mux2_1 U12410 ( .ip1(n10596), .ip2(n10595), .s(n11183), .op(n10600) );
  mux2_1 U12411 ( .ip1(\ANSWER/mem[4][0][1] ), .ip2(\ANSWER/mem[5][0][1] ), 
        .s(n10816), .op(n10598) );
  mux2_1 U12412 ( .ip1(\ANSWER/mem[6][0][1] ), .ip2(\ANSWER/mem[7][0][1] ), 
        .s(n10816), .op(n10597) );
  mux2_1 U12413 ( .ip1(n10598), .ip2(n10597), .s(n10968), .op(n10599) );
  mux2_1 U12414 ( .ip1(n10600), .ip2(n10599), .s(n11656), .op(n10602) );
  mux2_1 U12415 ( .ip1(\ANSWER/mem[8][0][1] ), .ip2(\ANSWER/mem[9][0][1] ), 
        .s(n10816), .op(n10601) );
  inv_1 U12416 ( .ip(n11996), .op(n10798) );
  mux2_1 U12417 ( .ip1(n10602), .ip2(n10601), .s(n10798), .op(n10603) );
  nand2_1 U12418 ( .ip1(n10603), .ip2(n12108), .op(n10675) );
  inv_1 U12419 ( .ip(n12109), .op(n10715) );
  mux2_1 U12420 ( .ip1(\ANSWER/mem[0][4][1] ), .ip2(\ANSWER/mem[1][4][1] ), 
        .s(n10715), .op(n10605) );
  mux2_1 U12421 ( .ip1(\ANSWER/mem[2][4][1] ), .ip2(\ANSWER/mem[3][4][1] ), 
        .s(n10715), .op(n10604) );
  mux2_1 U12422 ( .ip1(n10605), .ip2(n10604), .s(n11507), .op(n10609) );
  mux2_1 U12423 ( .ip1(\ANSWER/mem[4][4][1] ), .ip2(\ANSWER/mem[5][4][1] ), 
        .s(n10715), .op(n10607) );
  mux2_1 U12424 ( .ip1(\ANSWER/mem[6][4][1] ), .ip2(\ANSWER/mem[7][4][1] ), 
        .s(n10715), .op(n10606) );
  mux2_1 U12425 ( .ip1(n10607), .ip2(n10606), .s(n11090), .op(n10608) );
  mux2_1 U12426 ( .ip1(n10609), .ip2(n10608), .s(n11656), .op(n10611) );
  mux2_1 U12427 ( .ip1(\ANSWER/mem[8][4][1] ), .ip2(\ANSWER/mem[9][4][1] ), 
        .s(n10715), .op(n10610) );
  mux2_1 U12428 ( .ip1(n10611), .ip2(n10610), .s(n10798), .op(n10663) );
  buf_1 U12429 ( .ip(n10715), .op(n10797) );
  mux2_1 U12430 ( .ip1(\ANSWER/mem[0][7][1] ), .ip2(\ANSWER/mem[1][7][1] ), 
        .s(n10797), .op(n10613) );
  mux2_1 U12431 ( .ip1(\ANSWER/mem[2][7][1] ), .ip2(\ANSWER/mem[3][7][1] ), 
        .s(n10797), .op(n10612) );
  mux2_1 U12432 ( .ip1(n10613), .ip2(n10612), .s(n11090), .op(n10617) );
  mux2_1 U12433 ( .ip1(\ANSWER/mem[4][7][1] ), .ip2(\ANSWER/mem[5][7][1] ), 
        .s(n10797), .op(n10615) );
  mux2_1 U12434 ( .ip1(\ANSWER/mem[6][7][1] ), .ip2(\ANSWER/mem[7][7][1] ), 
        .s(n10797), .op(n10614) );
  mux2_1 U12435 ( .ip1(n10615), .ip2(n10614), .s(n11307), .op(n10616) );
  mux2_1 U12436 ( .ip1(n10617), .ip2(n10616), .s(n11656), .op(n10619) );
  mux2_1 U12437 ( .ip1(\ANSWER/mem[8][7][1] ), .ip2(\ANSWER/mem[9][7][1] ), 
        .s(n10715), .op(n10618) );
  mux2_1 U12438 ( .ip1(n10619), .ip2(n10618), .s(n10798), .op(n10620) );
  and2_1 U12439 ( .ip1(n12186), .ip2(n10620), .op(n10662) );
  mux2_1 U12440 ( .ip1(\ANSWER/mem[0][2][1] ), .ip2(\ANSWER/mem[1][2][1] ), 
        .s(n10816), .op(n10622) );
  mux2_1 U12441 ( .ip1(\ANSWER/mem[2][2][1] ), .ip2(\ANSWER/mem[3][2][1] ), 
        .s(n10816), .op(n10621) );
  mux2_1 U12442 ( .ip1(n10622), .ip2(n10621), .s(n11507), .op(n10626) );
  mux2_1 U12443 ( .ip1(\ANSWER/mem[4][2][1] ), .ip2(\ANSWER/mem[5][2][1] ), 
        .s(n10816), .op(n10624) );
  mux2_1 U12444 ( .ip1(\ANSWER/mem[6][2][1] ), .ip2(\ANSWER/mem[7][2][1] ), 
        .s(n10715), .op(n10623) );
  mux2_1 U12445 ( .ip1(n10624), .ip2(n10623), .s(n11307), .op(n10625) );
  mux2_1 U12446 ( .ip1(n10626), .ip2(n10625), .s(n11656), .op(n10628) );
  mux2_1 U12447 ( .ip1(\ANSWER/mem[8][2][1] ), .ip2(\ANSWER/mem[9][2][1] ), 
        .s(n10715), .op(n10627) );
  mux2_1 U12448 ( .ip1(n10628), .ip2(n10627), .s(n10798), .op(n10629) );
  nand2_1 U12449 ( .ip1(n12147), .ip2(n10629), .op(n10660) );
  mux2_1 U12450 ( .ip1(\ANSWER/mem[0][1][1] ), .ip2(\ANSWER/mem[1][1][1] ), 
        .s(n10816), .op(n10631) );
  mux2_1 U12451 ( .ip1(\ANSWER/mem[2][1][1] ), .ip2(\ANSWER/mem[3][1][1] ), 
        .s(n10816), .op(n10630) );
  mux2_1 U12452 ( .ip1(n10631), .ip2(n10630), .s(n11868), .op(n10635) );
  mux2_1 U12453 ( .ip1(\ANSWER/mem[4][1][1] ), .ip2(\ANSWER/mem[5][1][1] ), 
        .s(n10816), .op(n10633) );
  mux2_1 U12454 ( .ip1(\ANSWER/mem[6][1][1] ), .ip2(\ANSWER/mem[7][1][1] ), 
        .s(n10816), .op(n10632) );
  mux2_1 U12455 ( .ip1(n10633), .ip2(n10632), .s(n11976), .op(n10634) );
  mux2_1 U12456 ( .ip1(n10635), .ip2(n10634), .s(n11656), .op(n10637) );
  mux2_1 U12457 ( .ip1(\ANSWER/mem[8][1][1] ), .ip2(\ANSWER/mem[9][1][1] ), 
        .s(n10816), .op(n10636) );
  mux2_1 U12458 ( .ip1(n10637), .ip2(n10636), .s(n10798), .op(n10638) );
  nand2_1 U12459 ( .ip1(n12157), .ip2(n10638), .op(n10659) );
  mux2_1 U12460 ( .ip1(\ANSWER/mem[0][3][1] ), .ip2(\ANSWER/mem[1][3][1] ), 
        .s(n10715), .op(n10640) );
  mux2_1 U12461 ( .ip1(\ANSWER/mem[2][3][1] ), .ip2(\ANSWER/mem[3][3][1] ), 
        .s(n10715), .op(n10639) );
  mux2_1 U12462 ( .ip1(n10640), .ip2(n10639), .s(n11735), .op(n10644) );
  mux2_1 U12463 ( .ip1(\ANSWER/mem[4][3][1] ), .ip2(\ANSWER/mem[5][3][1] ), 
        .s(n10715), .op(n10642) );
  mux2_1 U12464 ( .ip1(\ANSWER/mem[6][3][1] ), .ip2(\ANSWER/mem[7][3][1] ), 
        .s(n10715), .op(n10641) );
  mux2_1 U12465 ( .ip1(n10642), .ip2(n10641), .s(n11950), .op(n10643) );
  mux2_1 U12466 ( .ip1(n10644), .ip2(n10643), .s(n11656), .op(n10646) );
  mux2_1 U12467 ( .ip1(\ANSWER/mem[8][3][1] ), .ip2(\ANSWER/mem[9][3][1] ), 
        .s(n10715), .op(n10645) );
  mux2_1 U12468 ( .ip1(n10646), .ip2(n10645), .s(n10798), .op(n10647) );
  nand2_1 U12469 ( .ip1(n12137), .ip2(n10647), .op(n10658) );
  mux2_1 U12470 ( .ip1(\ANSWER/mem[0][6][1] ), .ip2(\ANSWER/mem[1][6][1] ), 
        .s(n10797), .op(n10649) );
  mux2_1 U12471 ( .ip1(\ANSWER/mem[2][6][1] ), .ip2(\ANSWER/mem[3][6][1] ), 
        .s(n10797), .op(n10648) );
  mux2_1 U12472 ( .ip1(n10649), .ip2(n10648), .s(n11414), .op(n10653) );
  mux2_1 U12473 ( .ip1(\ANSWER/mem[4][6][1] ), .ip2(\ANSWER/mem[5][6][1] ), 
        .s(n10797), .op(n10651) );
  mux2_1 U12474 ( .ip1(\ANSWER/mem[6][6][1] ), .ip2(\ANSWER/mem[7][6][1] ), 
        .s(n10797), .op(n10650) );
  mux2_1 U12475 ( .ip1(n10651), .ip2(n10650), .s(n11735), .op(n10652) );
  mux2_1 U12476 ( .ip1(n10653), .ip2(n10652), .s(n11656), .op(n10655) );
  mux2_1 U12477 ( .ip1(\ANSWER/mem[8][6][1] ), .ip2(\ANSWER/mem[9][6][1] ), 
        .s(n10797), .op(n10654) );
  mux2_1 U12478 ( .ip1(n10655), .ip2(n10654), .s(n10798), .op(n10656) );
  nand2_1 U12479 ( .ip1(n12168), .ip2(n10656), .op(n10657) );
  nand4_1 U12480 ( .ip1(n10660), .ip2(n10659), .ip3(n10658), .ip4(n10657), 
        .op(n10661) );
  not_ab_or_c_or_d U12481 ( .ip1(n10663), .ip2(n12176), .ip3(n10662), .ip4(
        n10661), .op(n10674) );
  mux2_1 U12482 ( .ip1(\ANSWER/mem[0][5][1] ), .ip2(\ANSWER/mem[1][5][1] ), 
        .s(n10715), .op(n10665) );
  mux2_1 U12483 ( .ip1(\ANSWER/mem[2][5][1] ), .ip2(\ANSWER/mem[3][5][1] ), 
        .s(n10797), .op(n10664) );
  mux2_1 U12484 ( .ip1(n10665), .ip2(n10664), .s(n11868), .op(n10669) );
  mux2_1 U12485 ( .ip1(\ANSWER/mem[4][5][1] ), .ip2(\ANSWER/mem[5][5][1] ), 
        .s(n10797), .op(n10667) );
  mux2_1 U12486 ( .ip1(\ANSWER/mem[6][5][1] ), .ip2(\ANSWER/mem[7][5][1] ), 
        .s(n10797), .op(n10666) );
  mux2_1 U12487 ( .ip1(n10667), .ip2(n10666), .s(n11183), .op(n10668) );
  mux2_1 U12488 ( .ip1(n10669), .ip2(n10668), .s(n11656), .op(n10671) );
  mux2_1 U12489 ( .ip1(\ANSWER/mem[8][5][1] ), .ip2(\ANSWER/mem[9][5][1] ), 
        .s(n10797), .op(n10670) );
  mux2_1 U12490 ( .ip1(n10671), .ip2(n10670), .s(n10798), .op(n10672) );
  nand2_1 U12491 ( .ip1(n12127), .ip2(n10672), .op(n10673) );
  nand3_1 U12492 ( .ip1(n10675), .ip2(n10674), .ip3(n10673), .op(n10676) );
  nand2_1 U12493 ( .ip1(n10676), .ip2(n12190), .op(n10697) );
  mux2_1 U12494 ( .ip1(\ANSWER/mem[0][8][1] ), .ip2(\ANSWER/mem[1][8][1] ), 
        .s(n10715), .op(n10678) );
  mux2_1 U12495 ( .ip1(\ANSWER/mem[2][8][1] ), .ip2(\ANSWER/mem[3][8][1] ), 
        .s(n10797), .op(n10677) );
  mux2_1 U12496 ( .ip1(n10678), .ip2(n10677), .s(n11414), .op(n10682) );
  mux2_1 U12497 ( .ip1(\ANSWER/mem[4][8][1] ), .ip2(\ANSWER/mem[5][8][1] ), 
        .s(n10715), .op(n10680) );
  mux2_1 U12498 ( .ip1(\ANSWER/mem[6][8][1] ), .ip2(\ANSWER/mem[7][8][1] ), 
        .s(n10715), .op(n10679) );
  mux2_1 U12499 ( .ip1(n10680), .ip2(n10679), .s(n11868), .op(n10681) );
  mux2_1 U12500 ( .ip1(n10682), .ip2(n10681), .s(n11656), .op(n10684) );
  mux2_1 U12501 ( .ip1(\ANSWER/mem[8][8][1] ), .ip2(\ANSWER/mem[9][8][1] ), 
        .s(n10715), .op(n10683) );
  mux2_1 U12502 ( .ip1(n10684), .ip2(n10683), .s(n10798), .op(n10685) );
  nand2_1 U12503 ( .ip1(n12201), .ip2(n10685), .op(n10696) );
  mux2_1 U12504 ( .ip1(\ANSWER/mem[0][9][1] ), .ip2(\ANSWER/mem[1][9][1] ), 
        .s(n10797), .op(n10687) );
  mux2_1 U12505 ( .ip1(\ANSWER/mem[2][9][1] ), .ip2(\ANSWER/mem[3][9][1] ), 
        .s(n10797), .op(n10686) );
  mux2_1 U12506 ( .ip1(n10687), .ip2(n10686), .s(n11950), .op(n10691) );
  mux2_1 U12507 ( .ip1(\ANSWER/mem[4][9][1] ), .ip2(\ANSWER/mem[5][9][1] ), 
        .s(n10715), .op(n10689) );
  mux2_1 U12508 ( .ip1(\ANSWER/mem[6][9][1] ), .ip2(\ANSWER/mem[7][9][1] ), 
        .s(n10715), .op(n10688) );
  mux2_1 U12509 ( .ip1(n10689), .ip2(n10688), .s(n11224), .op(n10690) );
  mux2_1 U12510 ( .ip1(n10691), .ip2(n10690), .s(n11656), .op(n10693) );
  mux2_1 U12511 ( .ip1(\ANSWER/mem[8][9][1] ), .ip2(\ANSWER/mem[9][9][1] ), 
        .s(n10715), .op(n10692) );
  mux2_1 U12512 ( .ip1(n10693), .ip2(n10692), .s(n10798), .op(n10694) );
  nand2_1 U12513 ( .ip1(n12215), .ip2(n10694), .op(n10695) );
  nand3_1 U12514 ( .ip1(n10697), .ip2(n10696), .ip3(n10695), .op(\ANSWER/N486 ) );
  mux2_1 U12515 ( .ip1(\ANSWER/mem[0][3][2] ), .ip2(\ANSWER/mem[1][3][2] ), 
        .s(n10878), .op(n10699) );
  mux2_1 U12516 ( .ip1(\ANSWER/mem[2][3][2] ), .ip2(\ANSWER/mem[3][3][2] ), 
        .s(n10878), .op(n10698) );
  mux2_1 U12517 ( .ip1(n10699), .ip2(n10698), .s(n11090), .op(n10703) );
  mux2_1 U12518 ( .ip1(\ANSWER/mem[4][3][2] ), .ip2(\ANSWER/mem[5][3][2] ), 
        .s(n10878), .op(n10701) );
  mux2_1 U12519 ( .ip1(\ANSWER/mem[6][3][2] ), .ip2(\ANSWER/mem[7][3][2] ), 
        .s(n10878), .op(n10700) );
  mux2_1 U12520 ( .ip1(n10701), .ip2(n10700), .s(n10968), .op(n10702) );
  mux2_1 U12521 ( .ip1(n10703), .ip2(n10702), .s(n11937), .op(n10705) );
  buf_1 U12522 ( .ip(n10715), .op(n10821) );
  mux2_1 U12523 ( .ip1(\ANSWER/mem[8][3][2] ), .ip2(\ANSWER/mem[9][3][2] ), 
        .s(n10821), .op(n10704) );
  mux2_1 U12524 ( .ip1(n10705), .ip2(n10704), .s(n10798), .op(n10706) );
  nand2_1 U12525 ( .ip1(n12137), .ip2(n10706), .op(n10779) );
  mux2_1 U12526 ( .ip1(\ANSWER/mem[0][0][2] ), .ip2(\ANSWER/mem[1][0][2] ), 
        .s(n10821), .op(n10708) );
  mux2_1 U12527 ( .ip1(\ANSWER/mem[2][0][2] ), .ip2(\ANSWER/mem[3][0][2] ), 
        .s(n10821), .op(n10707) );
  mux2_1 U12528 ( .ip1(n10708), .ip2(n10707), .s(n11414), .op(n10712) );
  mux2_1 U12529 ( .ip1(\ANSWER/mem[4][0][2] ), .ip2(\ANSWER/mem[5][0][2] ), 
        .s(n10821), .op(n10710) );
  mux2_1 U12530 ( .ip1(\ANSWER/mem[6][0][2] ), .ip2(\ANSWER/mem[7][0][2] ), 
        .s(n10821), .op(n10709) );
  mux2_1 U12531 ( .ip1(n10710), .ip2(n10709), .s(n10968), .op(n10711) );
  mux2_1 U12532 ( .ip1(n10712), .ip2(n10711), .s(n11937), .op(n10714) );
  mux2_1 U12533 ( .ip1(\ANSWER/mem[8][0][2] ), .ip2(\ANSWER/mem[9][0][2] ), 
        .s(n10821), .op(n10713) );
  mux2_1 U12534 ( .ip1(n10714), .ip2(n10713), .s(n10798), .op(n10767) );
  mux2_1 U12535 ( .ip1(\ANSWER/mem[0][5][2] ), .ip2(\ANSWER/mem[1][5][2] ), 
        .s(n10821), .op(n10717) );
  buf_1 U12536 ( .ip(n10715), .op(n10792) );
  mux2_1 U12537 ( .ip1(\ANSWER/mem[2][5][2] ), .ip2(\ANSWER/mem[3][5][2] ), 
        .s(n10792), .op(n10716) );
  mux2_1 U12538 ( .ip1(n10717), .ip2(n10716), .s(n12062), .op(n10721) );
  mux2_1 U12539 ( .ip1(\ANSWER/mem[4][5][2] ), .ip2(\ANSWER/mem[5][5][2] ), 
        .s(n10792), .op(n10719) );
  mux2_1 U12540 ( .ip1(\ANSWER/mem[6][5][2] ), .ip2(\ANSWER/mem[7][5][2] ), 
        .s(n10792), .op(n10718) );
  mux2_1 U12541 ( .ip1(n10719), .ip2(n10718), .s(n11307), .op(n10720) );
  mux2_1 U12542 ( .ip1(n10721), .ip2(n10720), .s(n11937), .op(n10723) );
  mux2_1 U12543 ( .ip1(\ANSWER/mem[8][5][2] ), .ip2(\ANSWER/mem[9][5][2] ), 
        .s(n10792), .op(n10722) );
  mux2_1 U12544 ( .ip1(n10723), .ip2(n10722), .s(n10798), .op(n10724) );
  and2_1 U12545 ( .ip1(n12127), .ip2(n10724), .op(n10766) );
  mux2_1 U12546 ( .ip1(\ANSWER/mem[0][6][2] ), .ip2(\ANSWER/mem[1][6][2] ), 
        .s(n10792), .op(n10726) );
  mux2_1 U12547 ( .ip1(\ANSWER/mem[2][6][2] ), .ip2(\ANSWER/mem[3][6][2] ), 
        .s(n10792), .op(n10725) );
  mux2_1 U12548 ( .ip1(n10726), .ip2(n10725), .s(n10968), .op(n10730) );
  mux2_1 U12549 ( .ip1(\ANSWER/mem[4][6][2] ), .ip2(\ANSWER/mem[5][6][2] ), 
        .s(n10792), .op(n10728) );
  mux2_1 U12550 ( .ip1(\ANSWER/mem[6][6][2] ), .ip2(\ANSWER/mem[7][6][2] ), 
        .s(n10792), .op(n10727) );
  mux2_1 U12551 ( .ip1(n10728), .ip2(n10727), .s(n11414), .op(n10729) );
  mux2_1 U12552 ( .ip1(n10730), .ip2(n10729), .s(n11937), .op(n10732) );
  mux2_1 U12553 ( .ip1(\ANSWER/mem[8][6][2] ), .ip2(\ANSWER/mem[9][6][2] ), 
        .s(n10792), .op(n10731) );
  mux2_1 U12554 ( .ip1(n10732), .ip2(n10731), .s(n10798), .op(n10733) );
  nand2_1 U12555 ( .ip1(n12168), .ip2(n10733), .op(n10764) );
  mux2_1 U12556 ( .ip1(\ANSWER/mem[0][7][2] ), .ip2(\ANSWER/mem[1][7][2] ), 
        .s(n10792), .op(n10735) );
  mux2_1 U12557 ( .ip1(\ANSWER/mem[2][7][2] ), .ip2(\ANSWER/mem[3][7][2] ), 
        .s(n10792), .op(n10734) );
  mux2_1 U12558 ( .ip1(n10735), .ip2(n10734), .s(n11414), .op(n10739) );
  mux2_1 U12559 ( .ip1(\ANSWER/mem[4][7][2] ), .ip2(\ANSWER/mem[5][7][2] ), 
        .s(n10792), .op(n10737) );
  mux2_1 U12560 ( .ip1(\ANSWER/mem[6][7][2] ), .ip2(\ANSWER/mem[7][7][2] ), 
        .s(n10792), .op(n10736) );
  mux2_1 U12561 ( .ip1(n10737), .ip2(n10736), .s(n11950), .op(n10738) );
  mux2_1 U12562 ( .ip1(n10739), .ip2(n10738), .s(n11937), .op(n10741) );
  mux2_1 U12563 ( .ip1(\ANSWER/mem[8][7][2] ), .ip2(\ANSWER/mem[9][7][2] ), 
        .s(n10821), .op(n10740) );
  mux2_1 U12564 ( .ip1(n10741), .ip2(n10740), .s(n10798), .op(n10742) );
  nand2_1 U12565 ( .ip1(n12186), .ip2(n10742), .op(n10763) );
  mux2_1 U12566 ( .ip1(\ANSWER/mem[0][2][2] ), .ip2(\ANSWER/mem[1][2][2] ), 
        .s(n10821), .op(n10744) );
  mux2_1 U12567 ( .ip1(\ANSWER/mem[2][2][2] ), .ip2(\ANSWER/mem[3][2][2] ), 
        .s(n10821), .op(n10743) );
  mux2_1 U12568 ( .ip1(n10744), .ip2(n10743), .s(n11842), .op(n10748) );
  mux2_1 U12569 ( .ip1(\ANSWER/mem[4][2][2] ), .ip2(\ANSWER/mem[5][2][2] ), 
        .s(n10821), .op(n10746) );
  mux2_1 U12570 ( .ip1(\ANSWER/mem[6][2][2] ), .ip2(\ANSWER/mem[7][2][2] ), 
        .s(n10821), .op(n10745) );
  mux2_1 U12571 ( .ip1(n10746), .ip2(n10745), .s(n11950), .op(n10747) );
  mux2_1 U12572 ( .ip1(n10748), .ip2(n10747), .s(n11937), .op(n10750) );
  mux2_1 U12573 ( .ip1(\ANSWER/mem[8][2][2] ), .ip2(\ANSWER/mem[9][2][2] ), 
        .s(n10797), .op(n10749) );
  mux2_1 U12574 ( .ip1(n10750), .ip2(n10749), .s(n10798), .op(n10751) );
  nand2_1 U12575 ( .ip1(n12147), .ip2(n10751), .op(n10762) );
  mux2_1 U12576 ( .ip1(\ANSWER/mem[0][1][2] ), .ip2(\ANSWER/mem[1][1][2] ), 
        .s(n10821), .op(n10753) );
  mux2_1 U12577 ( .ip1(\ANSWER/mem[2][1][2] ), .ip2(\ANSWER/mem[3][1][2] ), 
        .s(n10821), .op(n10752) );
  mux2_1 U12578 ( .ip1(n10753), .ip2(n10752), .s(n11735), .op(n10757) );
  mux2_1 U12579 ( .ip1(\ANSWER/mem[4][1][2] ), .ip2(\ANSWER/mem[5][1][2] ), 
        .s(n10821), .op(n10755) );
  mux2_1 U12580 ( .ip1(\ANSWER/mem[6][1][2] ), .ip2(\ANSWER/mem[7][1][2] ), 
        .s(n10821), .op(n10754) );
  mux2_1 U12581 ( .ip1(n10755), .ip2(n10754), .s(n11735), .op(n10756) );
  mux2_1 U12582 ( .ip1(n10757), .ip2(n10756), .s(n11937), .op(n10759) );
  mux2_1 U12583 ( .ip1(\ANSWER/mem[8][1][2] ), .ip2(\ANSWER/mem[9][1][2] ), 
        .s(n10821), .op(n10758) );
  mux2_1 U12584 ( .ip1(n10759), .ip2(n10758), .s(n10798), .op(n10760) );
  nand2_1 U12585 ( .ip1(n12157), .ip2(n10760), .op(n10761) );
  nand4_1 U12586 ( .ip1(n10764), .ip2(n10763), .ip3(n10762), .ip4(n10761), 
        .op(n10765) );
  not_ab_or_c_or_d U12587 ( .ip1(n12108), .ip2(n10767), .ip3(n10766), .ip4(
        n10765), .op(n10778) );
  mux2_1 U12588 ( .ip1(\ANSWER/mem[0][4][2] ), .ip2(\ANSWER/mem[1][4][2] ), 
        .s(n10878), .op(n10769) );
  mux2_1 U12589 ( .ip1(\ANSWER/mem[2][4][2] ), .ip2(\ANSWER/mem[3][4][2] ), 
        .s(n10878), .op(n10768) );
  mux2_1 U12590 ( .ip1(n10769), .ip2(n10768), .s(n11224), .op(n10773) );
  mux2_1 U12591 ( .ip1(\ANSWER/mem[4][4][2] ), .ip2(\ANSWER/mem[5][4][2] ), 
        .s(n10878), .op(n10771) );
  mux2_1 U12592 ( .ip1(\ANSWER/mem[6][4][2] ), .ip2(\ANSWER/mem[7][4][2] ), 
        .s(n10878), .op(n10770) );
  mux2_1 U12593 ( .ip1(n10771), .ip2(n10770), .s(n12158), .op(n10772) );
  mux2_1 U12594 ( .ip1(n10773), .ip2(n10772), .s(n11937), .op(n10775) );
  inv_1 U12595 ( .ip(n12109), .op(n10906) );
  buf_1 U12596 ( .ip(n10906), .op(n10899) );
  mux2_1 U12597 ( .ip1(\ANSWER/mem[8][4][2] ), .ip2(\ANSWER/mem[9][4][2] ), 
        .s(n10899), .op(n10774) );
  mux2_1 U12598 ( .ip1(n10775), .ip2(n10774), .s(n10798), .op(n10776) );
  nand2_1 U12599 ( .ip1(n12176), .ip2(n10776), .op(n10777) );
  nand3_1 U12600 ( .ip1(n10779), .ip2(n10778), .ip3(n10777), .op(n10780) );
  nand2_1 U12601 ( .ip1(n10780), .ip2(n12190), .op(n10804) );
  mux2_1 U12602 ( .ip1(\ANSWER/mem[0][9][2] ), .ip2(\ANSWER/mem[1][9][2] ), 
        .s(n10878), .op(n10782) );
  mux2_1 U12603 ( .ip1(\ANSWER/mem[2][9][2] ), .ip2(\ANSWER/mem[3][9][2] ), 
        .s(n10878), .op(n10781) );
  mux2_1 U12604 ( .ip1(n10782), .ip2(n10781), .s(n11842), .op(n10786) );
  mux2_1 U12605 ( .ip1(\ANSWER/mem[4][9][2] ), .ip2(\ANSWER/mem[5][9][2] ), 
        .s(n10792), .op(n10784) );
  mux2_1 U12606 ( .ip1(\ANSWER/mem[6][9][2] ), .ip2(\ANSWER/mem[7][9][2] ), 
        .s(n10878), .op(n10783) );
  mux2_1 U12607 ( .ip1(n10784), .ip2(n10783), .s(n11976), .op(n10785) );
  mux2_1 U12608 ( .ip1(n10786), .ip2(n10785), .s(n11937), .op(n10788) );
  mux2_1 U12609 ( .ip1(\ANSWER/mem[8][9][2] ), .ip2(\ANSWER/mem[9][9][2] ), 
        .s(n10899), .op(n10787) );
  mux2_1 U12610 ( .ip1(n10788), .ip2(n10787), .s(n10798), .op(n10789) );
  nand2_1 U12611 ( .ip1(n12215), .ip2(n10789), .op(n10803) );
  mux2_1 U12612 ( .ip1(\ANSWER/mem[0][8][2] ), .ip2(\ANSWER/mem[1][8][2] ), 
        .s(n10878), .op(n10791) );
  mux2_1 U12613 ( .ip1(\ANSWER/mem[2][8][2] ), .ip2(\ANSWER/mem[3][8][2] ), 
        .s(n10878), .op(n10790) );
  mux2_1 U12614 ( .ip1(n10791), .ip2(n10790), .s(n12158), .op(n10796) );
  mux2_1 U12615 ( .ip1(\ANSWER/mem[4][8][2] ), .ip2(\ANSWER/mem[5][8][2] ), 
        .s(n10792), .op(n10794) );
  mux2_1 U12616 ( .ip1(\ANSWER/mem[6][8][2] ), .ip2(\ANSWER/mem[7][8][2] ), 
        .s(n10792), .op(n10793) );
  mux2_1 U12617 ( .ip1(n10794), .ip2(n10793), .s(n11868), .op(n10795) );
  mux2_1 U12618 ( .ip1(n10796), .ip2(n10795), .s(n11937), .op(n10800) );
  mux2_1 U12619 ( .ip1(\ANSWER/mem[8][8][2] ), .ip2(\ANSWER/mem[9][8][2] ), 
        .s(n10797), .op(n10799) );
  mux2_1 U12620 ( .ip1(n10800), .ip2(n10799), .s(n10798), .op(n10801) );
  nand2_1 U12621 ( .ip1(n12201), .ip2(n10801), .op(n10802) );
  nand3_1 U12622 ( .ip1(n10804), .ip2(n10803), .ip3(n10802), .op(\ANSWER/N485 ) );
  mux2_1 U12623 ( .ip1(\ANSWER/mem[0][0][3] ), .ip2(\ANSWER/mem[1][0][3] ), 
        .s(n10878), .op(n10806) );
  mux2_1 U12624 ( .ip1(\ANSWER/mem[2][0][3] ), .ip2(\ANSWER/mem[3][0][3] ), 
        .s(n10878), .op(n10805) );
  mux2_1 U12625 ( .ip1(n10806), .ip2(n10805), .s(n12158), .op(n10810) );
  mux2_1 U12626 ( .ip1(\ANSWER/mem[4][0][3] ), .ip2(\ANSWER/mem[5][0][3] ), 
        .s(n10878), .op(n10808) );
  mux2_1 U12627 ( .ip1(\ANSWER/mem[6][0][3] ), .ip2(\ANSWER/mem[7][0][3] ), 
        .s(n10878), .op(n10807) );
  mux2_1 U12628 ( .ip1(n10808), .ip2(n10807), .s(n11008), .op(n10809) );
  mux2_1 U12629 ( .ip1(n10810), .ip2(n10809), .s(n8821), .op(n10812) );
  mux2_1 U12630 ( .ip1(\ANSWER/mem[8][0][3] ), .ip2(\ANSWER/mem[9][0][3] ), 
        .s(n10878), .op(n10811) );
  inv_1 U12631 ( .ip(n11996), .op(n11188) );
  mux2_1 U12632 ( .ip1(n10812), .ip2(n10811), .s(n11188), .op(n10813) );
  nand2_1 U12633 ( .ip1(n12108), .ip2(n10813), .op(n10888) );
  mux2_1 U12634 ( .ip1(\ANSWER/mem[0][1][3] ), .ip2(\ANSWER/mem[1][1][3] ), 
        .s(n10816), .op(n10815) );
  mux2_1 U12635 ( .ip1(\ANSWER/mem[2][1][3] ), .ip2(\ANSWER/mem[3][1][3] ), 
        .s(n10816), .op(n10814) );
  mux2_1 U12636 ( .ip1(n10815), .ip2(n10814), .s(n11507), .op(n10820) );
  mux2_1 U12637 ( .ip1(\ANSWER/mem[4][1][3] ), .ip2(\ANSWER/mem[5][1][3] ), 
        .s(n10816), .op(n10818) );
  mux2_1 U12638 ( .ip1(\ANSWER/mem[6][1][3] ), .ip2(\ANSWER/mem[7][1][3] ), 
        .s(n10899), .op(n10817) );
  mux2_1 U12639 ( .ip1(n10818), .ip2(n10817), .s(n11008), .op(n10819) );
  mux2_1 U12640 ( .ip1(n10820), .ip2(n10819), .s(n8821), .op(n10823) );
  mux2_1 U12641 ( .ip1(\ANSWER/mem[8][1][3] ), .ip2(\ANSWER/mem[9][1][3] ), 
        .s(n10821), .op(n10822) );
  mux2_1 U12642 ( .ip1(n10823), .ip2(n10822), .s(n11188), .op(n10875) );
  mux2_1 U12643 ( .ip1(\ANSWER/mem[0][3][3] ), .ip2(\ANSWER/mem[1][3][3] ), 
        .s(n10906), .op(n10825) );
  mux2_1 U12644 ( .ip1(\ANSWER/mem[2][3][3] ), .ip2(\ANSWER/mem[3][3][3] ), 
        .s(n10906), .op(n10824) );
  mux2_1 U12645 ( .ip1(n10825), .ip2(n10824), .s(n11008), .op(n10829) );
  mux2_1 U12646 ( .ip1(\ANSWER/mem[4][3][3] ), .ip2(\ANSWER/mem[5][3][3] ), 
        .s(n10906), .op(n10827) );
  mux2_1 U12647 ( .ip1(\ANSWER/mem[6][3][3] ), .ip2(\ANSWER/mem[7][3][3] ), 
        .s(n10906), .op(n10826) );
  mux2_1 U12648 ( .ip1(n10827), .ip2(n10826), .s(n11307), .op(n10828) );
  mux2_1 U12649 ( .ip1(n10829), .ip2(n10828), .s(n8821), .op(n10831) );
  mux2_1 U12650 ( .ip1(\ANSWER/mem[8][3][3] ), .ip2(\ANSWER/mem[9][3][3] ), 
        .s(n10906), .op(n10830) );
  mux2_1 U12651 ( .ip1(n10831), .ip2(n10830), .s(n11188), .op(n10832) );
  and2_1 U12652 ( .ip1(n12137), .ip2(n10832), .op(n10874) );
  mux2_1 U12653 ( .ip1(\ANSWER/mem[0][5][3] ), .ip2(\ANSWER/mem[1][5][3] ), 
        .s(n10906), .op(n10834) );
  mux2_1 U12654 ( .ip1(\ANSWER/mem[2][5][3] ), .ip2(\ANSWER/mem[3][5][3] ), 
        .s(n10899), .op(n10833) );
  mux2_1 U12655 ( .ip1(n10834), .ip2(n10833), .s(n11008), .op(n10838) );
  mux2_1 U12656 ( .ip1(\ANSWER/mem[4][5][3] ), .ip2(\ANSWER/mem[5][5][3] ), 
        .s(n10899), .op(n10836) );
  mux2_1 U12657 ( .ip1(\ANSWER/mem[6][5][3] ), .ip2(\ANSWER/mem[7][5][3] ), 
        .s(n10899), .op(n10835) );
  mux2_1 U12658 ( .ip1(n10836), .ip2(n10835), .s(n11950), .op(n10837) );
  mux2_1 U12659 ( .ip1(n10838), .ip2(n10837), .s(n8821), .op(n10840) );
  mux2_1 U12660 ( .ip1(\ANSWER/mem[8][5][3] ), .ip2(\ANSWER/mem[9][5][3] ), 
        .s(n10899), .op(n10839) );
  mux2_1 U12661 ( .ip1(n10840), .ip2(n10839), .s(n11188), .op(n10841) );
  nand2_1 U12662 ( .ip1(n12127), .ip2(n10841), .op(n10872) );
  mux2_1 U12663 ( .ip1(\ANSWER/mem[0][7][3] ), .ip2(\ANSWER/mem[1][7][3] ), 
        .s(n10899), .op(n10843) );
  mux2_1 U12664 ( .ip1(\ANSWER/mem[2][7][3] ), .ip2(\ANSWER/mem[3][7][3] ), 
        .s(n10899), .op(n10842) );
  mux2_1 U12665 ( .ip1(n10843), .ip2(n10842), .s(n10968), .op(n10847) );
  mux2_1 U12666 ( .ip1(\ANSWER/mem[4][7][3] ), .ip2(\ANSWER/mem[5][7][3] ), 
        .s(n10899), .op(n10845) );
  mux2_1 U12667 ( .ip1(\ANSWER/mem[6][7][3] ), .ip2(\ANSWER/mem[7][7][3] ), 
        .s(n10899), .op(n10844) );
  mux2_1 U12668 ( .ip1(n10845), .ip2(n10844), .s(n12062), .op(n10846) );
  mux2_1 U12669 ( .ip1(n10847), .ip2(n10846), .s(n8821), .op(n10849) );
  mux2_1 U12670 ( .ip1(\ANSWER/mem[8][7][3] ), .ip2(\ANSWER/mem[9][7][3] ), 
        .s(n10906), .op(n10848) );
  mux2_1 U12671 ( .ip1(n10849), .ip2(n10848), .s(n11188), .op(n10850) );
  nand2_1 U12672 ( .ip1(n12186), .ip2(n10850), .op(n10871) );
  mux2_1 U12673 ( .ip1(\ANSWER/mem[0][4][3] ), .ip2(\ANSWER/mem[1][4][3] ), 
        .s(n10906), .op(n10852) );
  mux2_1 U12674 ( .ip1(\ANSWER/mem[2][4][3] ), .ip2(\ANSWER/mem[3][4][3] ), 
        .s(n10906), .op(n10851) );
  mux2_1 U12675 ( .ip1(n10852), .ip2(n10851), .s(n12062), .op(n10856) );
  mux2_1 U12676 ( .ip1(\ANSWER/mem[4][4][3] ), .ip2(\ANSWER/mem[5][4][3] ), 
        .s(n10906), .op(n10854) );
  mux2_1 U12677 ( .ip1(\ANSWER/mem[6][4][3] ), .ip2(\ANSWER/mem[7][4][3] ), 
        .s(n10906), .op(n10853) );
  mux2_1 U12678 ( .ip1(n10854), .ip2(n10853), .s(n11224), .op(n10855) );
  mux2_1 U12679 ( .ip1(n10856), .ip2(n10855), .s(n8821), .op(n10858) );
  mux2_1 U12680 ( .ip1(\ANSWER/mem[8][4][3] ), .ip2(\ANSWER/mem[9][4][3] ), 
        .s(n10906), .op(n10857) );
  mux2_1 U12681 ( .ip1(n10858), .ip2(n10857), .s(n11188), .op(n10859) );
  nand2_1 U12682 ( .ip1(n12176), .ip2(n10859), .op(n10870) );
  mux2_1 U12683 ( .ip1(\ANSWER/mem[0][6][3] ), .ip2(\ANSWER/mem[1][6][3] ), 
        .s(n10899), .op(n10861) );
  mux2_1 U12684 ( .ip1(\ANSWER/mem[2][6][3] ), .ip2(\ANSWER/mem[3][6][3] ), 
        .s(n10899), .op(n10860) );
  mux2_1 U12685 ( .ip1(n10861), .ip2(n10860), .s(n11842), .op(n10865) );
  mux2_1 U12686 ( .ip1(\ANSWER/mem[4][6][3] ), .ip2(\ANSWER/mem[5][6][3] ), 
        .s(n10899), .op(n10863) );
  mux2_1 U12687 ( .ip1(\ANSWER/mem[6][6][3] ), .ip2(\ANSWER/mem[7][6][3] ), 
        .s(n10899), .op(n10862) );
  mux2_1 U12688 ( .ip1(n10863), .ip2(n10862), .s(n11090), .op(n10864) );
  mux2_1 U12689 ( .ip1(n10865), .ip2(n10864), .s(n11979), .op(n10867) );
  mux2_1 U12690 ( .ip1(\ANSWER/mem[8][6][3] ), .ip2(\ANSWER/mem[9][6][3] ), 
        .s(n10899), .op(n10866) );
  mux2_1 U12691 ( .ip1(n10867), .ip2(n10866), .s(n11188), .op(n10868) );
  nand2_1 U12692 ( .ip1(n12168), .ip2(n10868), .op(n10869) );
  nand4_1 U12693 ( .ip1(n10872), .ip2(n10871), .ip3(n10870), .ip4(n10869), 
        .op(n10873) );
  not_ab_or_c_or_d U12694 ( .ip1(n12157), .ip2(n10875), .ip3(n10874), .ip4(
        n10873), .op(n10887) );
  mux2_1 U12695 ( .ip1(\ANSWER/mem[0][2][3] ), .ip2(\ANSWER/mem[1][2][3] ), 
        .s(n10878), .op(n10877) );
  mux2_1 U12696 ( .ip1(\ANSWER/mem[2][2][3] ), .ip2(\ANSWER/mem[3][2][3] ), 
        .s(n10878), .op(n10876) );
  mux2_1 U12697 ( .ip1(n10877), .ip2(n10876), .s(n11090), .op(n10882) );
  mux2_1 U12698 ( .ip1(\ANSWER/mem[4][2][3] ), .ip2(\ANSWER/mem[5][2][3] ), 
        .s(n10878), .op(n10880) );
  mux2_1 U12699 ( .ip1(\ANSWER/mem[6][2][3] ), .ip2(\ANSWER/mem[7][2][3] ), 
        .s(n10906), .op(n10879) );
  mux2_1 U12700 ( .ip1(n10880), .ip2(n10879), .s(n11183), .op(n10881) );
  mux2_1 U12701 ( .ip1(n10882), .ip2(n10881), .s(n8821), .op(n10884) );
  mux2_1 U12702 ( .ip1(\ANSWER/mem[8][2][3] ), .ip2(\ANSWER/mem[9][2][3] ), 
        .s(n10906), .op(n10883) );
  mux2_1 U12703 ( .ip1(n10884), .ip2(n10883), .s(n11188), .op(n10885) );
  nand2_1 U12704 ( .ip1(n12147), .ip2(n10885), .op(n10886) );
  nand3_1 U12705 ( .ip1(n10888), .ip2(n10887), .ip3(n10886), .op(n10889) );
  nand2_1 U12706 ( .ip1(n10889), .ip2(n12190), .op(n10912) );
  mux2_1 U12707 ( .ip1(\ANSWER/mem[0][8][3] ), .ip2(\ANSWER/mem[1][8][3] ), 
        .s(n10906), .op(n10891) );
  mux2_1 U12708 ( .ip1(\ANSWER/mem[2][8][3] ), .ip2(\ANSWER/mem[3][8][3] ), 
        .s(n10899), .op(n10890) );
  mux2_1 U12709 ( .ip1(n10891), .ip2(n10890), .s(n11735), .op(n10895) );
  mux2_1 U12710 ( .ip1(\ANSWER/mem[4][8][3] ), .ip2(\ANSWER/mem[5][8][3] ), 
        .s(n10906), .op(n10893) );
  mux2_1 U12711 ( .ip1(\ANSWER/mem[6][8][3] ), .ip2(\ANSWER/mem[7][8][3] ), 
        .s(n10906), .op(n10892) );
  mux2_1 U12712 ( .ip1(n10893), .ip2(n10892), .s(n11414), .op(n10894) );
  mux2_1 U12713 ( .ip1(n10895), .ip2(n10894), .s(n8821), .op(n10897) );
  mux2_1 U12714 ( .ip1(\ANSWER/mem[8][8][3] ), .ip2(\ANSWER/mem[9][8][3] ), 
        .s(n10906), .op(n10896) );
  mux2_1 U12715 ( .ip1(n10897), .ip2(n10896), .s(n11188), .op(n10898) );
  nand2_1 U12716 ( .ip1(n12201), .ip2(n10898), .op(n10911) );
  mux2_1 U12717 ( .ip1(\ANSWER/mem[0][9][3] ), .ip2(\ANSWER/mem[1][9][3] ), 
        .s(n10899), .op(n10901) );
  mux2_1 U12718 ( .ip1(\ANSWER/mem[2][9][3] ), .ip2(\ANSWER/mem[3][9][3] ), 
        .s(n10899), .op(n10900) );
  mux2_1 U12719 ( .ip1(n10901), .ip2(n10900), .s(n12158), .op(n10905) );
  mux2_1 U12720 ( .ip1(\ANSWER/mem[4][9][3] ), .ip2(\ANSWER/mem[5][9][3] ), 
        .s(n10906), .op(n10903) );
  mux2_1 U12721 ( .ip1(\ANSWER/mem[6][9][3] ), .ip2(\ANSWER/mem[7][9][3] ), 
        .s(n10906), .op(n10902) );
  mux2_1 U12722 ( .ip1(n10903), .ip2(n10902), .s(n11976), .op(n10904) );
  mux2_1 U12723 ( .ip1(n10905), .ip2(n10904), .s(n8821), .op(n10908) );
  mux2_1 U12724 ( .ip1(\ANSWER/mem[8][9][3] ), .ip2(\ANSWER/mem[9][9][3] ), 
        .s(n10906), .op(n10907) );
  mux2_1 U12725 ( .ip1(n10908), .ip2(n10907), .s(n11188), .op(n10909) );
  nand2_1 U12726 ( .ip1(n12215), .ip2(n10909), .op(n10910) );
  nand3_1 U12727 ( .ip1(n10912), .ip2(n10911), .ip3(n10910), .op(\ANSWER/N484 ) );
  mux2_1 U12728 ( .ip1(\ANSWER/mem[0][0][4] ), .ip2(\ANSWER/mem[1][0][4] ), 
        .s(n12204), .op(n10914) );
  mux2_1 U12729 ( .ip1(\ANSWER/mem[2][0][4] ), .ip2(\ANSWER/mem[3][0][4] ), 
        .s(n11007), .op(n10913) );
  inv_1 U12730 ( .ip(n12098), .op(n10968) );
  mux2_1 U12731 ( .ip1(n10914), .ip2(n10913), .s(n10968), .op(n10918) );
  mux2_1 U12732 ( .ip1(\ANSWER/mem[4][0][4] ), .ip2(\ANSWER/mem[5][0][4] ), 
        .s(n11223), .op(n10916) );
  mux2_1 U12733 ( .ip1(\ANSWER/mem[6][0][4] ), .ip2(\ANSWER/mem[7][0][4] ), 
        .s(n11651), .op(n10915) );
  mux2_1 U12734 ( .ip1(n10916), .ip2(n10915), .s(n10968), .op(n10917) );
  buf_1 U12735 ( .ip(n11454), .op(n12088) );
  mux2_1 U12736 ( .ip1(n10918), .ip2(n10917), .s(n12088), .op(n10920) );
  mux2_1 U12737 ( .ip1(\ANSWER/mem[8][0][4] ), .ip2(\ANSWER/mem[9][0][4] ), 
        .s(n11975), .op(n10919) );
  mux2_1 U12738 ( .ip1(n10920), .ip2(n10919), .s(n11188), .op(n10921) );
  nand2_1 U12739 ( .ip1(n10921), .ip2(n12108), .op(n10994) );
  inv_1 U12740 ( .ip(n12109), .op(n11013) );
  buf_1 U12741 ( .ip(n11013), .op(n11007) );
  mux2_1 U12742 ( .ip1(\ANSWER/mem[0][4][4] ), .ip2(\ANSWER/mem[1][4][4] ), 
        .s(n11007), .op(n10923) );
  mux2_1 U12743 ( .ip1(\ANSWER/mem[2][4][4] ), .ip2(\ANSWER/mem[3][4][4] ), 
        .s(n11007), .op(n10922) );
  mux2_1 U12744 ( .ip1(n10923), .ip2(n10922), .s(n10968), .op(n10927) );
  mux2_1 U12745 ( .ip1(\ANSWER/mem[4][4][4] ), .ip2(\ANSWER/mem[5][4][4] ), 
        .s(n11007), .op(n10925) );
  mux2_1 U12746 ( .ip1(\ANSWER/mem[6][4][4] ), .ip2(\ANSWER/mem[7][4][4] ), 
        .s(n11007), .op(n10924) );
  mux2_1 U12747 ( .ip1(n10925), .ip2(n10924), .s(n10968), .op(n10926) );
  mux2_1 U12748 ( .ip1(n10927), .ip2(n10926), .s(n12088), .op(n10929) );
  mux2_1 U12749 ( .ip1(\ANSWER/mem[8][4][4] ), .ip2(\ANSWER/mem[9][4][4] ), 
        .s(n11007), .op(n10928) );
  mux2_1 U12750 ( .ip1(n10929), .ip2(n10928), .s(n11188), .op(n10982) );
  mux2_1 U12751 ( .ip1(\ANSWER/mem[0][6][4] ), .ip2(\ANSWER/mem[1][6][4] ), 
        .s(n11013), .op(n10931) );
  mux2_1 U12752 ( .ip1(\ANSWER/mem[2][6][4] ), .ip2(\ANSWER/mem[3][6][4] ), 
        .s(n11013), .op(n10930) );
  mux2_1 U12753 ( .ip1(n10931), .ip2(n10930), .s(n10968), .op(n10935) );
  mux2_1 U12754 ( .ip1(\ANSWER/mem[4][6][4] ), .ip2(\ANSWER/mem[5][6][4] ), 
        .s(n11013), .op(n10933) );
  mux2_1 U12755 ( .ip1(\ANSWER/mem[6][6][4] ), .ip2(\ANSWER/mem[7][6][4] ), 
        .s(n11013), .op(n10932) );
  mux2_1 U12756 ( .ip1(n10933), .ip2(n10932), .s(n11008), .op(n10934) );
  mux2_1 U12757 ( .ip1(n10935), .ip2(n10934), .s(n12088), .op(n10937) );
  mux2_1 U12758 ( .ip1(\ANSWER/mem[8][6][4] ), .ip2(\ANSWER/mem[9][6][4] ), 
        .s(n11013), .op(n10936) );
  mux2_1 U12759 ( .ip1(n10937), .ip2(n10936), .s(n11188), .op(n10938) );
  and2_1 U12760 ( .ip1(n12168), .ip2(n10938), .op(n10981) );
  mux2_1 U12761 ( .ip1(\ANSWER/mem[0][2][4] ), .ip2(\ANSWER/mem[1][2][4] ), 
        .s(n11223), .op(n10940) );
  mux2_1 U12762 ( .ip1(\ANSWER/mem[2][2][4] ), .ip2(\ANSWER/mem[3][2][4] ), 
        .s(n10816), .op(n10939) );
  mux2_1 U12763 ( .ip1(n10940), .ip2(n10939), .s(n10968), .op(n10944) );
  mux2_1 U12764 ( .ip1(\ANSWER/mem[4][2][4] ), .ip2(\ANSWER/mem[5][2][4] ), 
        .s(n11651), .op(n10942) );
  mux2_1 U12765 ( .ip1(\ANSWER/mem[6][2][4] ), .ip2(\ANSWER/mem[7][2][4] ), 
        .s(n11007), .op(n10941) );
  mux2_1 U12766 ( .ip1(n10942), .ip2(n10941), .s(n10968), .op(n10943) );
  mux2_1 U12767 ( .ip1(n10944), .ip2(n10943), .s(n12088), .op(n10946) );
  mux2_1 U12768 ( .ip1(\ANSWER/mem[8][2][4] ), .ip2(\ANSWER/mem[9][2][4] ), 
        .s(n11007), .op(n10945) );
  mux2_1 U12769 ( .ip1(n10946), .ip2(n10945), .s(n11188), .op(n10947) );
  nand2_1 U12770 ( .ip1(n12147), .ip2(n10947), .op(n10979) );
  mux2_1 U12771 ( .ip1(\ANSWER/mem[0][5][4] ), .ip2(\ANSWER/mem[1][5][4] ), 
        .s(n11007), .op(n10949) );
  mux2_1 U12772 ( .ip1(\ANSWER/mem[2][5][4] ), .ip2(\ANSWER/mem[3][5][4] ), 
        .s(n11007), .op(n10948) );
  mux2_1 U12773 ( .ip1(n10949), .ip2(n10948), .s(n10968), .op(n10953) );
  mux2_1 U12774 ( .ip1(\ANSWER/mem[4][5][4] ), .ip2(\ANSWER/mem[5][5][4] ), 
        .s(n11013), .op(n10951) );
  mux2_1 U12775 ( .ip1(\ANSWER/mem[6][5][4] ), .ip2(\ANSWER/mem[7][5][4] ), 
        .s(n11013), .op(n10950) );
  mux2_1 U12776 ( .ip1(n10951), .ip2(n10950), .s(n10968), .op(n10952) );
  mux2_1 U12777 ( .ip1(n10953), .ip2(n10952), .s(n12088), .op(n10955) );
  mux2_1 U12778 ( .ip1(\ANSWER/mem[8][5][4] ), .ip2(\ANSWER/mem[9][5][4] ), 
        .s(n11013), .op(n10954) );
  mux2_1 U12779 ( .ip1(n10955), .ip2(n10954), .s(n11188), .op(n10956) );
  nand2_1 U12780 ( .ip1(n12127), .ip2(n10956), .op(n10978) );
  mux2_1 U12781 ( .ip1(\ANSWER/mem[0][1][4] ), .ip2(\ANSWER/mem[1][1][4] ), 
        .s(n11113), .op(n10958) );
  mux2_1 U12782 ( .ip1(\ANSWER/mem[2][1][4] ), .ip2(\ANSWER/mem[3][1][4] ), 
        .s(n10583), .op(n10957) );
  mux2_1 U12783 ( .ip1(n10958), .ip2(n10957), .s(n10968), .op(n10962) );
  mux2_1 U12784 ( .ip1(\ANSWER/mem[4][1][4] ), .ip2(\ANSWER/mem[5][1][4] ), 
        .s(n11007), .op(n10960) );
  mux2_1 U12785 ( .ip1(\ANSWER/mem[6][1][4] ), .ip2(\ANSWER/mem[7][1][4] ), 
        .s(n11873), .op(n10959) );
  mux2_1 U12786 ( .ip1(n10960), .ip2(n10959), .s(n10968), .op(n10961) );
  mux2_1 U12787 ( .ip1(n10962), .ip2(n10961), .s(n12088), .op(n10964) );
  mux2_1 U12788 ( .ip1(\ANSWER/mem[8][1][4] ), .ip2(\ANSWER/mem[9][1][4] ), 
        .s(n11328), .op(n10963) );
  mux2_1 U12789 ( .ip1(n10964), .ip2(n10963), .s(n11188), .op(n10965) );
  nand2_1 U12790 ( .ip1(n12157), .ip2(n10965), .op(n10977) );
  mux2_1 U12791 ( .ip1(\ANSWER/mem[0][3][4] ), .ip2(\ANSWER/mem[1][3][4] ), 
        .s(n11007), .op(n10967) );
  mux2_1 U12792 ( .ip1(\ANSWER/mem[2][3][4] ), .ip2(\ANSWER/mem[3][3][4] ), 
        .s(n11007), .op(n10966) );
  mux2_1 U12793 ( .ip1(n10967), .ip2(n10966), .s(n10968), .op(n10972) );
  mux2_1 U12794 ( .ip1(\ANSWER/mem[4][3][4] ), .ip2(\ANSWER/mem[5][3][4] ), 
        .s(n11007), .op(n10970) );
  mux2_1 U12795 ( .ip1(\ANSWER/mem[6][3][4] ), .ip2(\ANSWER/mem[7][3][4] ), 
        .s(n11007), .op(n10969) );
  mux2_1 U12796 ( .ip1(n10970), .ip2(n10969), .s(n10968), .op(n10971) );
  mux2_1 U12797 ( .ip1(n10972), .ip2(n10971), .s(n12088), .op(n10974) );
  mux2_1 U12798 ( .ip1(\ANSWER/mem[8][3][4] ), .ip2(\ANSWER/mem[9][3][4] ), 
        .s(n11007), .op(n10973) );
  mux2_1 U12799 ( .ip1(n10974), .ip2(n10973), .s(n11188), .op(n10975) );
  nand2_1 U12800 ( .ip1(n12137), .ip2(n10975), .op(n10976) );
  nand4_1 U12801 ( .ip1(n10979), .ip2(n10978), .ip3(n10977), .ip4(n10976), 
        .op(n10980) );
  not_ab_or_c_or_d U12802 ( .ip1(n12176), .ip2(n10982), .ip3(n10981), .ip4(
        n10980), .op(n10993) );
  mux2_1 U12803 ( .ip1(\ANSWER/mem[0][7][4] ), .ip2(\ANSWER/mem[1][7][4] ), 
        .s(n11013), .op(n10984) );
  mux2_1 U12804 ( .ip1(\ANSWER/mem[2][7][4] ), .ip2(\ANSWER/mem[3][7][4] ), 
        .s(n11013), .op(n10983) );
  mux2_1 U12805 ( .ip1(n10984), .ip2(n10983), .s(n11008), .op(n10988) );
  mux2_1 U12806 ( .ip1(\ANSWER/mem[4][7][4] ), .ip2(\ANSWER/mem[5][7][4] ), 
        .s(n11013), .op(n10986) );
  mux2_1 U12807 ( .ip1(\ANSWER/mem[6][7][4] ), .ip2(\ANSWER/mem[7][7][4] ), 
        .s(n11013), .op(n10985) );
  mux2_1 U12808 ( .ip1(n10986), .ip2(n10985), .s(n11008), .op(n10987) );
  mux2_1 U12809 ( .ip1(n10988), .ip2(n10987), .s(n12088), .op(n10990) );
  mux2_1 U12810 ( .ip1(\ANSWER/mem[8][7][4] ), .ip2(\ANSWER/mem[9][7][4] ), 
        .s(n11013), .op(n10989) );
  mux2_1 U12811 ( .ip1(n10990), .ip2(n10989), .s(n11188), .op(n10991) );
  nand2_1 U12812 ( .ip1(n12186), .ip2(n10991), .op(n10992) );
  nand3_1 U12813 ( .ip1(n10994), .ip2(n10993), .ip3(n10992), .op(n10995) );
  nand2_1 U12814 ( .ip1(n10995), .ip2(n12190), .op(n11019) );
  mux2_1 U12815 ( .ip1(\ANSWER/mem[0][8][4] ), .ip2(\ANSWER/mem[1][8][4] ), 
        .s(n11013), .op(n10997) );
  mux2_1 U12816 ( .ip1(\ANSWER/mem[2][8][4] ), .ip2(\ANSWER/mem[3][8][4] ), 
        .s(n11007), .op(n10996) );
  mux2_1 U12817 ( .ip1(n10997), .ip2(n10996), .s(n11008), .op(n11001) );
  mux2_1 U12818 ( .ip1(\ANSWER/mem[4][8][4] ), .ip2(\ANSWER/mem[5][8][4] ), 
        .s(n11013), .op(n10999) );
  mux2_1 U12819 ( .ip1(\ANSWER/mem[6][8][4] ), .ip2(\ANSWER/mem[7][8][4] ), 
        .s(n11013), .op(n10998) );
  mux2_1 U12820 ( .ip1(n10999), .ip2(n10998), .s(n11008), .op(n11000) );
  mux2_1 U12821 ( .ip1(n11001), .ip2(n11000), .s(n12088), .op(n11003) );
  mux2_1 U12822 ( .ip1(\ANSWER/mem[8][8][4] ), .ip2(\ANSWER/mem[9][8][4] ), 
        .s(n11013), .op(n11002) );
  mux2_1 U12823 ( .ip1(n11003), .ip2(n11002), .s(n11188), .op(n11004) );
  nand2_1 U12824 ( .ip1(n12201), .ip2(n11004), .op(n11018) );
  mux2_1 U12825 ( .ip1(\ANSWER/mem[0][9][4] ), .ip2(\ANSWER/mem[1][9][4] ), 
        .s(n11013), .op(n11006) );
  mux2_1 U12826 ( .ip1(\ANSWER/mem[2][9][4] ), .ip2(\ANSWER/mem[3][9][4] ), 
        .s(n11007), .op(n11005) );
  mux2_1 U12827 ( .ip1(n11006), .ip2(n11005), .s(n11008), .op(n11012) );
  mux2_1 U12828 ( .ip1(\ANSWER/mem[4][9][4] ), .ip2(\ANSWER/mem[5][9][4] ), 
        .s(n11013), .op(n11010) );
  mux2_1 U12829 ( .ip1(\ANSWER/mem[6][9][4] ), .ip2(\ANSWER/mem[7][9][4] ), 
        .s(n11007), .op(n11009) );
  mux2_1 U12830 ( .ip1(n11010), .ip2(n11009), .s(n11008), .op(n11011) );
  mux2_1 U12831 ( .ip1(n11012), .ip2(n11011), .s(n12088), .op(n11015) );
  mux2_1 U12832 ( .ip1(\ANSWER/mem[8][9][4] ), .ip2(\ANSWER/mem[9][9][4] ), 
        .s(n11013), .op(n11014) );
  mux2_1 U12833 ( .ip1(n11015), .ip2(n11014), .s(n11188), .op(n11016) );
  nand2_1 U12834 ( .ip1(n12215), .ip2(n11016), .op(n11017) );
  nand3_1 U12835 ( .ip1(n11019), .ip2(n11018), .ip3(n11017), .op(\ANSWER/N483 ) );
  inv_1 U12836 ( .ip(n12109), .op(n11070) );
  mux2_1 U12837 ( .ip1(\ANSWER/mem[0][0][5] ), .ip2(\ANSWER/mem[1][0][5] ), 
        .s(n11070), .op(n11021) );
  mux2_1 U12838 ( .ip1(\ANSWER/mem[2][0][5] ), .ip2(\ANSWER/mem[3][0][5] ), 
        .s(n11070), .op(n11020) );
  inv_1 U12839 ( .ip(n12098), .op(n11090) );
  mux2_1 U12840 ( .ip1(n11021), .ip2(n11020), .s(n11090), .op(n11025) );
  mux2_1 U12841 ( .ip1(\ANSWER/mem[4][0][5] ), .ip2(\ANSWER/mem[5][0][5] ), 
        .s(n11070), .op(n11023) );
  mux2_1 U12842 ( .ip1(\ANSWER/mem[6][0][5] ), .ip2(\ANSWER/mem[7][0][5] ), 
        .s(n11070), .op(n11022) );
  mux2_1 U12843 ( .ip1(n11023), .ip2(n11022), .s(n11090), .op(n11024) );
  buf_1 U12844 ( .ip(n11656), .op(n12207) );
  mux2_1 U12845 ( .ip1(n11025), .ip2(n11024), .s(n12207), .op(n11027) );
  mux2_1 U12846 ( .ip1(\ANSWER/mem[8][0][5] ), .ip2(\ANSWER/mem[9][0][5] ), 
        .s(n11070), .op(n11026) );
  mux2_1 U12847 ( .ip1(n11027), .ip2(n11026), .s(n11565), .op(n11028) );
  nand2_1 U12848 ( .ip1(n11028), .ip2(n12108), .op(n11102) );
  mux2_1 U12849 ( .ip1(\ANSWER/mem[0][2][5] ), .ip2(\ANSWER/mem[1][2][5] ), 
        .s(n11070), .op(n11030) );
  mux2_1 U12850 ( .ip1(\ANSWER/mem[2][2][5] ), .ip2(\ANSWER/mem[3][2][5] ), 
        .s(n11070), .op(n11029) );
  mux2_1 U12851 ( .ip1(n11030), .ip2(n11029), .s(n11090), .op(n11034) );
  mux2_1 U12852 ( .ip1(\ANSWER/mem[4][2][5] ), .ip2(\ANSWER/mem[5][2][5] ), 
        .s(n11070), .op(n11032) );
  inv_1 U12853 ( .ip(n12109), .op(n11120) );
  buf_1 U12854 ( .ip(n11120), .op(n11113) );
  mux2_1 U12855 ( .ip1(\ANSWER/mem[6][2][5] ), .ip2(\ANSWER/mem[7][2][5] ), 
        .s(n11113), .op(n11031) );
  mux2_1 U12856 ( .ip1(n11032), .ip2(n11031), .s(n11090), .op(n11033) );
  mux2_1 U12857 ( .ip1(n11034), .ip2(n11033), .s(n12207), .op(n11036) );
  mux2_1 U12858 ( .ip1(\ANSWER/mem[8][2][5] ), .ip2(\ANSWER/mem[9][2][5] ), 
        .s(n11113), .op(n11035) );
  mux2_1 U12859 ( .ip1(n11036), .ip2(n11035), .s(n11565), .op(n11089) );
  mux2_1 U12860 ( .ip1(\ANSWER/mem[0][4][5] ), .ip2(\ANSWER/mem[1][4][5] ), 
        .s(n11113), .op(n11038) );
  mux2_1 U12861 ( .ip1(\ANSWER/mem[2][4][5] ), .ip2(\ANSWER/mem[3][4][5] ), 
        .s(n11113), .op(n11037) );
  mux2_1 U12862 ( .ip1(n11038), .ip2(n11037), .s(n11090), .op(n11042) );
  mux2_1 U12863 ( .ip1(\ANSWER/mem[4][4][5] ), .ip2(\ANSWER/mem[5][4][5] ), 
        .s(n11113), .op(n11040) );
  mux2_1 U12864 ( .ip1(\ANSWER/mem[6][4][5] ), .ip2(\ANSWER/mem[7][4][5] ), 
        .s(n11113), .op(n11039) );
  mux2_1 U12865 ( .ip1(n11040), .ip2(n11039), .s(n11090), .op(n11041) );
  mux2_1 U12866 ( .ip1(n11042), .ip2(n11041), .s(n12207), .op(n11044) );
  mux2_1 U12867 ( .ip1(\ANSWER/mem[8][4][5] ), .ip2(\ANSWER/mem[9][4][5] ), 
        .s(n11113), .op(n11043) );
  mux2_1 U12868 ( .ip1(n11044), .ip2(n11043), .s(n11565), .op(n11045) );
  and2_1 U12869 ( .ip1(n12176), .ip2(n11045), .op(n11088) );
  mux2_1 U12870 ( .ip1(\ANSWER/mem[0][7][5] ), .ip2(\ANSWER/mem[1][7][5] ), 
        .s(n11120), .op(n11047) );
  mux2_1 U12871 ( .ip1(\ANSWER/mem[2][7][5] ), .ip2(\ANSWER/mem[3][7][5] ), 
        .s(n11120), .op(n11046) );
  mux2_1 U12872 ( .ip1(n11047), .ip2(n11046), .s(n11950), .op(n11051) );
  mux2_1 U12873 ( .ip1(\ANSWER/mem[4][7][5] ), .ip2(\ANSWER/mem[5][7][5] ), 
        .s(n11120), .op(n11049) );
  mux2_1 U12874 ( .ip1(\ANSWER/mem[6][7][5] ), .ip2(\ANSWER/mem[7][7][5] ), 
        .s(n11120), .op(n11048) );
  mux2_1 U12875 ( .ip1(n11049), .ip2(n11048), .s(n11976), .op(n11050) );
  mux2_1 U12876 ( .ip1(n11051), .ip2(n11050), .s(n12207), .op(n11053) );
  mux2_1 U12877 ( .ip1(\ANSWER/mem[8][7][5] ), .ip2(\ANSWER/mem[9][7][5] ), 
        .s(n11120), .op(n11052) );
  mux2_1 U12878 ( .ip1(n11053), .ip2(n11052), .s(n11565), .op(n11054) );
  nand2_1 U12879 ( .ip1(n12186), .ip2(n11054), .op(n11086) );
  mux2_1 U12880 ( .ip1(\ANSWER/mem[0][5][5] ), .ip2(\ANSWER/mem[1][5][5] ), 
        .s(n11113), .op(n11056) );
  mux2_1 U12881 ( .ip1(\ANSWER/mem[2][5][5] ), .ip2(\ANSWER/mem[3][5][5] ), 
        .s(n11120), .op(n11055) );
  mux2_1 U12882 ( .ip1(n11056), .ip2(n11055), .s(n11090), .op(n11060) );
  mux2_1 U12883 ( .ip1(\ANSWER/mem[4][5][5] ), .ip2(\ANSWER/mem[5][5][5] ), 
        .s(n11120), .op(n11058) );
  mux2_1 U12884 ( .ip1(\ANSWER/mem[6][5][5] ), .ip2(\ANSWER/mem[7][5][5] ), 
        .s(n11120), .op(n11057) );
  mux2_1 U12885 ( .ip1(n11058), .ip2(n11057), .s(n11090), .op(n11059) );
  mux2_1 U12886 ( .ip1(n11060), .ip2(n11059), .s(n12207), .op(n11062) );
  mux2_1 U12887 ( .ip1(\ANSWER/mem[8][5][5] ), .ip2(\ANSWER/mem[9][5][5] ), 
        .s(n11120), .op(n11061) );
  mux2_1 U12888 ( .ip1(n11062), .ip2(n11061), .s(n11565), .op(n11063) );
  nand2_1 U12889 ( .ip1(n12127), .ip2(n11063), .op(n11085) );
  mux2_1 U12890 ( .ip1(\ANSWER/mem[0][1][5] ), .ip2(\ANSWER/mem[1][1][5] ), 
        .s(n11070), .op(n11065) );
  mux2_1 U12891 ( .ip1(\ANSWER/mem[2][1][5] ), .ip2(\ANSWER/mem[3][1][5] ), 
        .s(n11070), .op(n11064) );
  mux2_1 U12892 ( .ip1(n11065), .ip2(n11064), .s(n11090), .op(n11069) );
  mux2_1 U12893 ( .ip1(\ANSWER/mem[4][1][5] ), .ip2(\ANSWER/mem[5][1][5] ), 
        .s(n11070), .op(n11067) );
  mux2_1 U12894 ( .ip1(\ANSWER/mem[6][1][5] ), .ip2(\ANSWER/mem[7][1][5] ), 
        .s(n11070), .op(n11066) );
  mux2_1 U12895 ( .ip1(n11067), .ip2(n11066), .s(n11090), .op(n11068) );
  mux2_1 U12896 ( .ip1(n11069), .ip2(n11068), .s(n12207), .op(n11072) );
  mux2_1 U12897 ( .ip1(\ANSWER/mem[8][1][5] ), .ip2(\ANSWER/mem[9][1][5] ), 
        .s(n11070), .op(n11071) );
  mux2_1 U12898 ( .ip1(n11072), .ip2(n11071), .s(n11565), .op(n11073) );
  nand2_1 U12899 ( .ip1(n12157), .ip2(n11073), .op(n11084) );
  mux2_1 U12900 ( .ip1(\ANSWER/mem[0][3][5] ), .ip2(\ANSWER/mem[1][3][5] ), 
        .s(n11113), .op(n11075) );
  mux2_1 U12901 ( .ip1(\ANSWER/mem[2][3][5] ), .ip2(\ANSWER/mem[3][3][5] ), 
        .s(n11113), .op(n11074) );
  mux2_1 U12902 ( .ip1(n11075), .ip2(n11074), .s(n11090), .op(n11079) );
  mux2_1 U12903 ( .ip1(\ANSWER/mem[4][3][5] ), .ip2(\ANSWER/mem[5][3][5] ), 
        .s(n11113), .op(n11077) );
  mux2_1 U12904 ( .ip1(\ANSWER/mem[6][3][5] ), .ip2(\ANSWER/mem[7][3][5] ), 
        .s(n11113), .op(n11076) );
  mux2_1 U12905 ( .ip1(n11077), .ip2(n11076), .s(n11090), .op(n11078) );
  mux2_1 U12906 ( .ip1(n11079), .ip2(n11078), .s(n12207), .op(n11081) );
  mux2_1 U12907 ( .ip1(\ANSWER/mem[8][3][5] ), .ip2(\ANSWER/mem[9][3][5] ), 
        .s(n11113), .op(n11080) );
  mux2_1 U12908 ( .ip1(n11081), .ip2(n11080), .s(n11188), .op(n11082) );
  nand2_1 U12909 ( .ip1(n12137), .ip2(n11082), .op(n11083) );
  nand4_1 U12910 ( .ip1(n11086), .ip2(n11085), .ip3(n11084), .ip4(n11083), 
        .op(n11087) );
  not_ab_or_c_or_d U12911 ( .ip1(n11089), .ip2(n12147), .ip3(n11088), .ip4(
        n11087), .op(n11101) );
  mux2_1 U12912 ( .ip1(\ANSWER/mem[0][6][5] ), .ip2(\ANSWER/mem[1][6][5] ), 
        .s(n11120), .op(n11092) );
  mux2_1 U12913 ( .ip1(\ANSWER/mem[2][6][5] ), .ip2(\ANSWER/mem[3][6][5] ), 
        .s(n11120), .op(n11091) );
  mux2_1 U12914 ( .ip1(n11092), .ip2(n11091), .s(n11090), .op(n11096) );
  mux2_1 U12915 ( .ip1(\ANSWER/mem[4][6][5] ), .ip2(\ANSWER/mem[5][6][5] ), 
        .s(n11120), .op(n11094) );
  mux2_1 U12916 ( .ip1(\ANSWER/mem[6][6][5] ), .ip2(\ANSWER/mem[7][6][5] ), 
        .s(n11120), .op(n11093) );
  mux2_1 U12917 ( .ip1(n11094), .ip2(n11093), .s(n11090), .op(n11095) );
  mux2_1 U12918 ( .ip1(n11096), .ip2(n11095), .s(n12207), .op(n11098) );
  mux2_1 U12919 ( .ip1(\ANSWER/mem[8][6][5] ), .ip2(\ANSWER/mem[9][6][5] ), 
        .s(n11120), .op(n11097) );
  mux2_1 U12920 ( .ip1(n11098), .ip2(n11097), .s(n11565), .op(n11099) );
  nand2_1 U12921 ( .ip1(n12168), .ip2(n11099), .op(n11100) );
  nand3_1 U12922 ( .ip1(n11102), .ip2(n11101), .ip3(n11100), .op(n11103) );
  nand2_1 U12923 ( .ip1(n11103), .ip2(n12190), .op(n11126) );
  mux2_1 U12924 ( .ip1(\ANSWER/mem[0][9][5] ), .ip2(\ANSWER/mem[1][9][5] ), 
        .s(n11120), .op(n11105) );
  mux2_1 U12925 ( .ip1(\ANSWER/mem[2][9][5] ), .ip2(\ANSWER/mem[3][9][5] ), 
        .s(n11113), .op(n11104) );
  mux2_1 U12926 ( .ip1(n11105), .ip2(n11104), .s(n12158), .op(n11109) );
  mux2_1 U12927 ( .ip1(\ANSWER/mem[4][9][5] ), .ip2(\ANSWER/mem[5][9][5] ), 
        .s(n11120), .op(n11107) );
  mux2_1 U12928 ( .ip1(\ANSWER/mem[6][9][5] ), .ip2(\ANSWER/mem[7][9][5] ), 
        .s(n11120), .op(n11106) );
  mux2_1 U12929 ( .ip1(n11107), .ip2(n11106), .s(n11090), .op(n11108) );
  mux2_1 U12930 ( .ip1(n11109), .ip2(n11108), .s(n12207), .op(n11111) );
  mux2_1 U12931 ( .ip1(\ANSWER/mem[8][9][5] ), .ip2(\ANSWER/mem[9][9][5] ), 
        .s(n11120), .op(n11110) );
  mux2_1 U12932 ( .ip1(n11111), .ip2(n11110), .s(n11565), .op(n11112) );
  nand2_1 U12933 ( .ip1(n12215), .ip2(n11112), .op(n11125) );
  mux2_1 U12934 ( .ip1(\ANSWER/mem[0][8][5] ), .ip2(\ANSWER/mem[1][8][5] ), 
        .s(n11113), .op(n11115) );
  mux2_1 U12935 ( .ip1(\ANSWER/mem[2][8][5] ), .ip2(\ANSWER/mem[3][8][5] ), 
        .s(n11113), .op(n11114) );
  mux2_1 U12936 ( .ip1(n11115), .ip2(n11114), .s(n10968), .op(n11119) );
  mux2_1 U12937 ( .ip1(\ANSWER/mem[4][8][5] ), .ip2(\ANSWER/mem[5][8][5] ), 
        .s(n11120), .op(n11117) );
  mux2_1 U12938 ( .ip1(\ANSWER/mem[6][8][5] ), .ip2(\ANSWER/mem[7][8][5] ), 
        .s(n11120), .op(n11116) );
  mux2_1 U12939 ( .ip1(n11117), .ip2(n11116), .s(n11224), .op(n11118) );
  mux2_1 U12940 ( .ip1(n11119), .ip2(n11118), .s(n12207), .op(n11122) );
  mux2_1 U12941 ( .ip1(\ANSWER/mem[8][8][5] ), .ip2(\ANSWER/mem[9][8][5] ), 
        .s(n11120), .op(n11121) );
  mux2_1 U12942 ( .ip1(n11122), .ip2(n11121), .s(n11565), .op(n11123) );
  nand2_1 U12943 ( .ip1(n12201), .ip2(n11123), .op(n11124) );
  nand3_1 U12944 ( .ip1(n11126), .ip2(n11125), .ip3(n11124), .op(\ANSWER/N482 ) );
  inv_1 U12945 ( .ip(n12109), .op(n11164) );
  mux2_1 U12946 ( .ip1(\ANSWER/mem[0][0][6] ), .ip2(\ANSWER/mem[1][0][6] ), 
        .s(n11164), .op(n11128) );
  mux2_1 U12947 ( .ip1(\ANSWER/mem[2][0][6] ), .ip2(\ANSWER/mem[3][0][6] ), 
        .s(n11164), .op(n11127) );
  inv_1 U12948 ( .ip(n12098), .op(n11183) );
  mux2_1 U12949 ( .ip1(n11128), .ip2(n11127), .s(n11183), .op(n11132) );
  mux2_1 U12950 ( .ip1(\ANSWER/mem[4][0][6] ), .ip2(\ANSWER/mem[5][0][6] ), 
        .s(n11164), .op(n11130) );
  mux2_1 U12951 ( .ip1(\ANSWER/mem[6][0][6] ), .ip2(\ANSWER/mem[7][0][6] ), 
        .s(n11164), .op(n11129) );
  mux2_1 U12952 ( .ip1(n11130), .ip2(n11129), .s(n11183), .op(n11131) );
  mux2_1 U12953 ( .ip1(n11132), .ip2(n11131), .s(n8821), .op(n11134) );
  mux2_1 U12954 ( .ip1(\ANSWER/mem[8][0][6] ), .ip2(\ANSWER/mem[9][0][6] ), 
        .s(n11164), .op(n11133) );
  mux2_1 U12955 ( .ip1(n11134), .ip2(n11133), .s(n11565), .op(n11135) );
  nand2_1 U12956 ( .ip1(n11135), .ip2(n12108), .op(n11210) );
  mux2_1 U12957 ( .ip1(\ANSWER/mem[0][1][6] ), .ip2(\ANSWER/mem[1][1][6] ), 
        .s(n11164), .op(n11137) );
  mux2_1 U12958 ( .ip1(\ANSWER/mem[2][1][6] ), .ip2(\ANSWER/mem[3][1][6] ), 
        .s(n11164), .op(n11136) );
  mux2_1 U12959 ( .ip1(n11137), .ip2(n11136), .s(n11183), .op(n11141) );
  mux2_1 U12960 ( .ip1(\ANSWER/mem[4][1][6] ), .ip2(\ANSWER/mem[5][1][6] ), 
        .s(n11164), .op(n11139) );
  mux2_1 U12961 ( .ip1(\ANSWER/mem[6][1][6] ), .ip2(\ANSWER/mem[7][1][6] ), 
        .s(n11164), .op(n11138) );
  mux2_1 U12962 ( .ip1(n11139), .ip2(n11138), .s(n11183), .op(n11140) );
  mux2_1 U12963 ( .ip1(n11141), .ip2(n11140), .s(n8821), .op(n11143) );
  mux2_1 U12964 ( .ip1(\ANSWER/mem[8][1][6] ), .ip2(\ANSWER/mem[9][1][6] ), 
        .s(n11164), .op(n11142) );
  mux2_1 U12965 ( .ip1(n11143), .ip2(n11142), .s(n11565), .op(n11198) );
  inv_1 U12966 ( .ip(n12109), .op(n11229) );
  mux2_1 U12967 ( .ip1(\ANSWER/mem[0][6][6] ), .ip2(\ANSWER/mem[1][6][6] ), 
        .s(n11229), .op(n11145) );
  mux2_1 U12968 ( .ip1(\ANSWER/mem[2][6][6] ), .ip2(\ANSWER/mem[3][6][6] ), 
        .s(n11229), .op(n11144) );
  mux2_1 U12969 ( .ip1(n11145), .ip2(n11144), .s(n11183), .op(n11149) );
  mux2_1 U12970 ( .ip1(\ANSWER/mem[4][6][6] ), .ip2(\ANSWER/mem[5][6][6] ), 
        .s(n11229), .op(n11147) );
  mux2_1 U12971 ( .ip1(\ANSWER/mem[6][6][6] ), .ip2(\ANSWER/mem[7][6][6] ), 
        .s(n11229), .op(n11146) );
  mux2_1 U12972 ( .ip1(n11147), .ip2(n11146), .s(n11224), .op(n11148) );
  mux2_1 U12973 ( .ip1(n11149), .ip2(n11148), .s(n8821), .op(n11151) );
  mux2_1 U12974 ( .ip1(\ANSWER/mem[8][6][6] ), .ip2(\ANSWER/mem[9][6][6] ), 
        .s(n11229), .op(n11150) );
  mux2_1 U12975 ( .ip1(n11151), .ip2(n11150), .s(n11565), .op(n11152) );
  and2_1 U12976 ( .ip1(n12168), .ip2(n11152), .op(n11197) );
  buf_1 U12977 ( .ip(n11229), .op(n11223) );
  mux2_1 U12978 ( .ip1(\ANSWER/mem[0][5][6] ), .ip2(\ANSWER/mem[1][5][6] ), 
        .s(n11223), .op(n11154) );
  mux2_1 U12979 ( .ip1(\ANSWER/mem[2][5][6] ), .ip2(\ANSWER/mem[3][5][6] ), 
        .s(n11229), .op(n11153) );
  mux2_1 U12980 ( .ip1(n11154), .ip2(n11153), .s(n11183), .op(n11158) );
  mux2_1 U12981 ( .ip1(\ANSWER/mem[4][5][6] ), .ip2(\ANSWER/mem[5][5][6] ), 
        .s(n11229), .op(n11156) );
  mux2_1 U12982 ( .ip1(\ANSWER/mem[6][5][6] ), .ip2(\ANSWER/mem[7][5][6] ), 
        .s(n11229), .op(n11155) );
  mux2_1 U12983 ( .ip1(n11156), .ip2(n11155), .s(n11183), .op(n11157) );
  mux2_1 U12984 ( .ip1(n11158), .ip2(n11157), .s(n8821), .op(n11160) );
  mux2_1 U12985 ( .ip1(\ANSWER/mem[8][5][6] ), .ip2(\ANSWER/mem[9][5][6] ), 
        .s(n11229), .op(n11159) );
  mux2_1 U12986 ( .ip1(n11160), .ip2(n11159), .s(n11565), .op(n11161) );
  nand2_1 U12987 ( .ip1(n12127), .ip2(n11161), .op(n11195) );
  mux2_1 U12988 ( .ip1(\ANSWER/mem[0][2][6] ), .ip2(\ANSWER/mem[1][2][6] ), 
        .s(n11164), .op(n11163) );
  mux2_1 U12989 ( .ip1(\ANSWER/mem[2][2][6] ), .ip2(\ANSWER/mem[3][2][6] ), 
        .s(n11164), .op(n11162) );
  mux2_1 U12990 ( .ip1(n11163), .ip2(n11162), .s(n11183), .op(n11168) );
  mux2_1 U12991 ( .ip1(\ANSWER/mem[4][2][6] ), .ip2(\ANSWER/mem[5][2][6] ), 
        .s(n11164), .op(n11166) );
  mux2_1 U12992 ( .ip1(\ANSWER/mem[6][2][6] ), .ip2(\ANSWER/mem[7][2][6] ), 
        .s(n11223), .op(n11165) );
  mux2_1 U12993 ( .ip1(n11166), .ip2(n11165), .s(n11183), .op(n11167) );
  mux2_1 U12994 ( .ip1(n11168), .ip2(n11167), .s(n8821), .op(n11170) );
  mux2_1 U12995 ( .ip1(\ANSWER/mem[8][2][6] ), .ip2(\ANSWER/mem[9][2][6] ), 
        .s(n11223), .op(n11169) );
  mux2_1 U12996 ( .ip1(n11170), .ip2(n11169), .s(n11565), .op(n11171) );
  nand2_1 U12997 ( .ip1(n12147), .ip2(n11171), .op(n11194) );
  mux2_1 U12998 ( .ip1(\ANSWER/mem[0][4][6] ), .ip2(\ANSWER/mem[1][4][6] ), 
        .s(n11223), .op(n11173) );
  mux2_1 U12999 ( .ip1(\ANSWER/mem[2][4][6] ), .ip2(\ANSWER/mem[3][4][6] ), 
        .s(n11223), .op(n11172) );
  mux2_1 U13000 ( .ip1(n11173), .ip2(n11172), .s(n11183), .op(n11177) );
  mux2_1 U13001 ( .ip1(\ANSWER/mem[4][4][6] ), .ip2(\ANSWER/mem[5][4][6] ), 
        .s(n11223), .op(n11175) );
  mux2_1 U13002 ( .ip1(\ANSWER/mem[6][4][6] ), .ip2(\ANSWER/mem[7][4][6] ), 
        .s(n11223), .op(n11174) );
  mux2_1 U13003 ( .ip1(n11175), .ip2(n11174), .s(n11183), .op(n11176) );
  mux2_1 U13004 ( .ip1(n11177), .ip2(n11176), .s(n11454), .op(n11179) );
  mux2_1 U13005 ( .ip1(\ANSWER/mem[8][4][6] ), .ip2(\ANSWER/mem[9][4][6] ), 
        .s(n11223), .op(n11178) );
  mux2_1 U13006 ( .ip1(n11179), .ip2(n11178), .s(n11565), .op(n11180) );
  nand2_1 U13007 ( .ip1(n12176), .ip2(n11180), .op(n11193) );
  mux2_1 U13008 ( .ip1(\ANSWER/mem[0][3][6] ), .ip2(\ANSWER/mem[1][3][6] ), 
        .s(n11223), .op(n11182) );
  mux2_1 U13009 ( .ip1(\ANSWER/mem[2][3][6] ), .ip2(\ANSWER/mem[3][3][6] ), 
        .s(n11223), .op(n11181) );
  mux2_1 U13010 ( .ip1(n11182), .ip2(n11181), .s(n11183), .op(n11187) );
  mux2_1 U13011 ( .ip1(\ANSWER/mem[4][3][6] ), .ip2(\ANSWER/mem[5][3][6] ), 
        .s(n11223), .op(n11185) );
  mux2_1 U13012 ( .ip1(\ANSWER/mem[6][3][6] ), .ip2(\ANSWER/mem[7][3][6] ), 
        .s(n11223), .op(n11184) );
  mux2_1 U13013 ( .ip1(n11185), .ip2(n11184), .s(n11183), .op(n11186) );
  mux2_1 U13014 ( .ip1(n11187), .ip2(n11186), .s(n8821), .op(n11190) );
  mux2_1 U13015 ( .ip1(\ANSWER/mem[8][3][6] ), .ip2(\ANSWER/mem[9][3][6] ), 
        .s(n11223), .op(n11189) );
  mux2_1 U13016 ( .ip1(n11190), .ip2(n11189), .s(n11188), .op(n11191) );
  nand2_1 U13017 ( .ip1(n12137), .ip2(n11191), .op(n11192) );
  nand4_1 U13018 ( .ip1(n11195), .ip2(n11194), .ip3(n11193), .ip4(n11192), 
        .op(n11196) );
  not_ab_or_c_or_d U13019 ( .ip1(n11198), .ip2(n12157), .ip3(n11197), .ip4(
        n11196), .op(n11209) );
  mux2_1 U13020 ( .ip1(\ANSWER/mem[0][7][6] ), .ip2(\ANSWER/mem[1][7][6] ), 
        .s(n11229), .op(n11200) );
  mux2_1 U13021 ( .ip1(\ANSWER/mem[2][7][6] ), .ip2(\ANSWER/mem[3][7][6] ), 
        .s(n11229), .op(n11199) );
  mux2_1 U13022 ( .ip1(n11200), .ip2(n11199), .s(n11224), .op(n11204) );
  mux2_1 U13023 ( .ip1(\ANSWER/mem[4][7][6] ), .ip2(\ANSWER/mem[5][7][6] ), 
        .s(n11229), .op(n11202) );
  mux2_1 U13024 ( .ip1(\ANSWER/mem[6][7][6] ), .ip2(\ANSWER/mem[7][7][6] ), 
        .s(n11229), .op(n11201) );
  mux2_1 U13025 ( .ip1(n11202), .ip2(n11201), .s(n11224), .op(n11203) );
  mux2_1 U13026 ( .ip1(n11204), .ip2(n11203), .s(n8821), .op(n11206) );
  mux2_1 U13027 ( .ip1(\ANSWER/mem[8][7][6] ), .ip2(\ANSWER/mem[9][7][6] ), 
        .s(n11229), .op(n11205) );
  mux2_1 U13028 ( .ip1(n11206), .ip2(n11205), .s(n11565), .op(n11207) );
  nand2_1 U13029 ( .ip1(n12186), .ip2(n11207), .op(n11208) );
  nand3_1 U13030 ( .ip1(n11210), .ip2(n11209), .ip3(n11208), .op(n11211) );
  nand2_1 U13031 ( .ip1(n11211), .ip2(n12190), .op(n11235) );
  mux2_1 U13032 ( .ip1(\ANSWER/mem[0][8][6] ), .ip2(\ANSWER/mem[1][8][6] ), 
        .s(n11229), .op(n11213) );
  mux2_1 U13033 ( .ip1(\ANSWER/mem[2][8][6] ), .ip2(\ANSWER/mem[3][8][6] ), 
        .s(n11223), .op(n11212) );
  mux2_1 U13034 ( .ip1(n11213), .ip2(n11212), .s(n11224), .op(n11217) );
  mux2_1 U13035 ( .ip1(\ANSWER/mem[4][8][6] ), .ip2(\ANSWER/mem[5][8][6] ), 
        .s(n11229), .op(n11215) );
  mux2_1 U13036 ( .ip1(\ANSWER/mem[6][8][6] ), .ip2(\ANSWER/mem[7][8][6] ), 
        .s(n11229), .op(n11214) );
  mux2_1 U13037 ( .ip1(n11215), .ip2(n11214), .s(n11224), .op(n11216) );
  mux2_1 U13038 ( .ip1(n11217), .ip2(n11216), .s(n8821), .op(n11219) );
  mux2_1 U13039 ( .ip1(\ANSWER/mem[8][8][6] ), .ip2(\ANSWER/mem[9][8][6] ), 
        .s(n11229), .op(n11218) );
  mux2_1 U13040 ( .ip1(n11219), .ip2(n11218), .s(n11565), .op(n11220) );
  nand2_1 U13041 ( .ip1(n12201), .ip2(n11220), .op(n11234) );
  mux2_1 U13042 ( .ip1(\ANSWER/mem[0][9][6] ), .ip2(\ANSWER/mem[1][9][6] ), 
        .s(n11229), .op(n11222) );
  mux2_1 U13043 ( .ip1(\ANSWER/mem[2][9][6] ), .ip2(\ANSWER/mem[3][9][6] ), 
        .s(n11223), .op(n11221) );
  mux2_1 U13044 ( .ip1(n11222), .ip2(n11221), .s(n11224), .op(n11228) );
  mux2_1 U13045 ( .ip1(\ANSWER/mem[4][9][6] ), .ip2(\ANSWER/mem[5][9][6] ), 
        .s(n11229), .op(n11226) );
  mux2_1 U13046 ( .ip1(\ANSWER/mem[6][9][6] ), .ip2(\ANSWER/mem[7][9][6] ), 
        .s(n11223), .op(n11225) );
  mux2_1 U13047 ( .ip1(n11226), .ip2(n11225), .s(n11224), .op(n11227) );
  mux2_1 U13048 ( .ip1(n11228), .ip2(n11227), .s(n8821), .op(n11231) );
  mux2_1 U13049 ( .ip1(\ANSWER/mem[8][9][6] ), .ip2(\ANSWER/mem[9][9][6] ), 
        .s(n11229), .op(n11230) );
  mux2_1 U13050 ( .ip1(n11231), .ip2(n11230), .s(n11565), .op(n11232) );
  nand2_1 U13051 ( .ip1(n12215), .ip2(n11232), .op(n11233) );
  nand3_1 U13052 ( .ip1(n11235), .ip2(n11234), .ip3(n11233), .op(\ANSWER/N481 ) );
  mux2_1 U13053 ( .ip1(\ANSWER/mem[0][0][7] ), .ip2(\ANSWER/mem[1][0][7] ), 
        .s(n8833), .op(n11237) );
  mux2_1 U13054 ( .ip1(\ANSWER/mem[2][0][7] ), .ip2(\ANSWER/mem[3][0][7] ), 
        .s(n8833), .op(n11236) );
  inv_1 U13055 ( .ip(n12098), .op(n11307) );
  mux2_1 U13056 ( .ip1(n11237), .ip2(n11236), .s(n11307), .op(n11241) );
  mux2_1 U13057 ( .ip1(\ANSWER/mem[4][0][7] ), .ip2(\ANSWER/mem[5][0][7] ), 
        .s(n8833), .op(n11239) );
  mux2_1 U13058 ( .ip1(\ANSWER/mem[6][0][7] ), .ip2(\ANSWER/mem[7][0][7] ), 
        .s(n8833), .op(n11238) );
  mux2_1 U13059 ( .ip1(n11239), .ip2(n11238), .s(n11307), .op(n11240) );
  mux2_1 U13060 ( .ip1(n11241), .ip2(n11240), .s(n11979), .op(n11243) );
  mux2_1 U13061 ( .ip1(\ANSWER/mem[8][0][7] ), .ip2(\ANSWER/mem[9][0][7] ), 
        .s(n8833), .op(n11242) );
  mux2_1 U13062 ( .ip1(n11243), .ip2(n11242), .s(n11336), .op(n11244) );
  nand2_1 U13063 ( .ip1(n12108), .ip2(n11244), .op(n11317) );
  inv_1 U13064 ( .ip(n12109), .op(n11335) );
  buf_1 U13065 ( .ip(n11335), .op(n11328) );
  mux2_1 U13066 ( .ip1(\ANSWER/mem[0][3][7] ), .ip2(\ANSWER/mem[1][3][7] ), 
        .s(n11328), .op(n11246) );
  mux2_1 U13067 ( .ip1(\ANSWER/mem[2][3][7] ), .ip2(\ANSWER/mem[3][3][7] ), 
        .s(n11328), .op(n11245) );
  mux2_1 U13068 ( .ip1(n11246), .ip2(n11245), .s(n11307), .op(n11250) );
  mux2_1 U13069 ( .ip1(\ANSWER/mem[4][3][7] ), .ip2(\ANSWER/mem[5][3][7] ), 
        .s(n11328), .op(n11248) );
  mux2_1 U13070 ( .ip1(\ANSWER/mem[6][3][7] ), .ip2(\ANSWER/mem[7][3][7] ), 
        .s(n11328), .op(n11247) );
  mux2_1 U13071 ( .ip1(n11248), .ip2(n11247), .s(n11307), .op(n11249) );
  mux2_1 U13072 ( .ip1(n11250), .ip2(n11249), .s(n11979), .op(n11252) );
  mux2_1 U13073 ( .ip1(\ANSWER/mem[8][3][7] ), .ip2(\ANSWER/mem[9][3][7] ), 
        .s(n11328), .op(n11251) );
  mux2_1 U13074 ( .ip1(n11252), .ip2(n11251), .s(n11336), .op(n11304) );
  mux2_1 U13075 ( .ip1(\ANSWER/mem[0][6][7] ), .ip2(\ANSWER/mem[1][6][7] ), 
        .s(n11335), .op(n11254) );
  mux2_1 U13076 ( .ip1(\ANSWER/mem[2][6][7] ), .ip2(\ANSWER/mem[3][6][7] ), 
        .s(n11335), .op(n11253) );
  mux2_1 U13077 ( .ip1(n11254), .ip2(n11253), .s(n11307), .op(n11258) );
  mux2_1 U13078 ( .ip1(\ANSWER/mem[4][6][7] ), .ip2(\ANSWER/mem[5][6][7] ), 
        .s(n11335), .op(n11256) );
  mux2_1 U13079 ( .ip1(\ANSWER/mem[6][6][7] ), .ip2(\ANSWER/mem[7][6][7] ), 
        .s(n11335), .op(n11255) );
  mux2_1 U13080 ( .ip1(n11256), .ip2(n11255), .s(n11507), .op(n11257) );
  mux2_1 U13081 ( .ip1(n11258), .ip2(n11257), .s(n11937), .op(n11260) );
  mux2_1 U13082 ( .ip1(\ANSWER/mem[8][6][7] ), .ip2(\ANSWER/mem[9][6][7] ), 
        .s(n11335), .op(n11259) );
  mux2_1 U13083 ( .ip1(n11260), .ip2(n11259), .s(n11336), .op(n11261) );
  and2_1 U13084 ( .ip1(n12168), .ip2(n11261), .op(n11303) );
  mux2_1 U13085 ( .ip1(\ANSWER/mem[0][5][7] ), .ip2(\ANSWER/mem[1][5][7] ), 
        .s(n11328), .op(n11263) );
  mux2_1 U13086 ( .ip1(\ANSWER/mem[2][5][7] ), .ip2(\ANSWER/mem[3][5][7] ), 
        .s(n11335), .op(n11262) );
  mux2_1 U13087 ( .ip1(n11263), .ip2(n11262), .s(n11307), .op(n11267) );
  mux2_1 U13088 ( .ip1(\ANSWER/mem[4][5][7] ), .ip2(\ANSWER/mem[5][5][7] ), 
        .s(n11335), .op(n11265) );
  mux2_1 U13089 ( .ip1(\ANSWER/mem[6][5][7] ), .ip2(\ANSWER/mem[7][5][7] ), 
        .s(n11335), .op(n11264) );
  mux2_1 U13090 ( .ip1(n11265), .ip2(n11264), .s(n11307), .op(n11266) );
  mux2_1 U13091 ( .ip1(n11267), .ip2(n11266), .s(n11937), .op(n11269) );
  mux2_1 U13092 ( .ip1(\ANSWER/mem[8][5][7] ), .ip2(\ANSWER/mem[9][5][7] ), 
        .s(n11335), .op(n11268) );
  mux2_1 U13093 ( .ip1(n11269), .ip2(n11268), .s(n11565), .op(n11270) );
  nand2_1 U13094 ( .ip1(n12127), .ip2(n11270), .op(n11301) );
  mux2_1 U13095 ( .ip1(\ANSWER/mem[0][4][7] ), .ip2(\ANSWER/mem[1][4][7] ), 
        .s(n11328), .op(n11272) );
  mux2_1 U13096 ( .ip1(\ANSWER/mem[2][4][7] ), .ip2(\ANSWER/mem[3][4][7] ), 
        .s(n11328), .op(n11271) );
  mux2_1 U13097 ( .ip1(n11272), .ip2(n11271), .s(n11307), .op(n11276) );
  mux2_1 U13098 ( .ip1(\ANSWER/mem[4][4][7] ), .ip2(\ANSWER/mem[5][4][7] ), 
        .s(n11328), .op(n11274) );
  mux2_1 U13099 ( .ip1(\ANSWER/mem[6][4][7] ), .ip2(\ANSWER/mem[7][4][7] ), 
        .s(n11328), .op(n11273) );
  mux2_1 U13100 ( .ip1(n11274), .ip2(n11273), .s(n11307), .op(n11275) );
  mux2_1 U13101 ( .ip1(n11276), .ip2(n11275), .s(n11937), .op(n11278) );
  mux2_1 U13102 ( .ip1(\ANSWER/mem[8][4][7] ), .ip2(\ANSWER/mem[9][4][7] ), 
        .s(n11328), .op(n11277) );
  mux2_1 U13103 ( .ip1(n11278), .ip2(n11277), .s(n11552), .op(n11279) );
  nand2_1 U13104 ( .ip1(n12176), .ip2(n11279), .op(n11300) );
  mux2_1 U13105 ( .ip1(\ANSWER/mem[0][7][7] ), .ip2(\ANSWER/mem[1][7][7] ), 
        .s(n11335), .op(n11281) );
  mux2_1 U13106 ( .ip1(\ANSWER/mem[2][7][7] ), .ip2(\ANSWER/mem[3][7][7] ), 
        .s(n11335), .op(n11280) );
  mux2_1 U13107 ( .ip1(n11281), .ip2(n11280), .s(n11842), .op(n11285) );
  mux2_1 U13108 ( .ip1(\ANSWER/mem[4][7][7] ), .ip2(\ANSWER/mem[5][7][7] ), 
        .s(n11335), .op(n11283) );
  mux2_1 U13109 ( .ip1(\ANSWER/mem[6][7][7] ), .ip2(\ANSWER/mem[7][7][7] ), 
        .s(n11335), .op(n11282) );
  mux2_1 U13110 ( .ip1(n11283), .ip2(n11282), .s(n12062), .op(n11284) );
  mux2_1 U13111 ( .ip1(n11285), .ip2(n11284), .s(n11937), .op(n11287) );
  mux2_1 U13112 ( .ip1(\ANSWER/mem[8][7][7] ), .ip2(\ANSWER/mem[9][7][7] ), 
        .s(n11335), .op(n11286) );
  mux2_1 U13113 ( .ip1(n11287), .ip2(n11286), .s(n11565), .op(n11288) );
  nand2_1 U13114 ( .ip1(n12186), .ip2(n11288), .op(n11299) );
  mux2_1 U13115 ( .ip1(\ANSWER/mem[0][1][7] ), .ip2(\ANSWER/mem[1][1][7] ), 
        .s(n11506), .op(n11290) );
  mux2_1 U13116 ( .ip1(\ANSWER/mem[2][1][7] ), .ip2(\ANSWER/mem[3][1][7] ), 
        .s(n8833), .op(n11289) );
  mux2_1 U13117 ( .ip1(n11290), .ip2(n11289), .s(n11307), .op(n11294) );
  mux2_1 U13118 ( .ip1(\ANSWER/mem[4][1][7] ), .ip2(\ANSWER/mem[5][1][7] ), 
        .s(n11546), .op(n11292) );
  mux2_1 U13119 ( .ip1(\ANSWER/mem[6][1][7] ), .ip2(\ANSWER/mem[7][1][7] ), 
        .s(n11506), .op(n11291) );
  mux2_1 U13120 ( .ip1(n11292), .ip2(n11291), .s(n11307), .op(n11293) );
  mux2_1 U13121 ( .ip1(n11294), .ip2(n11293), .s(n11937), .op(n11296) );
  mux2_1 U13122 ( .ip1(\ANSWER/mem[8][1][7] ), .ip2(\ANSWER/mem[9][1][7] ), 
        .s(n8833), .op(n11295) );
  mux2_1 U13123 ( .ip1(n11296), .ip2(n11295), .s(n11336), .op(n11297) );
  nand2_1 U13124 ( .ip1(n12157), .ip2(n11297), .op(n11298) );
  nand4_1 U13125 ( .ip1(n11301), .ip2(n11300), .ip3(n11299), .ip4(n11298), 
        .op(n11302) );
  not_ab_or_c_or_d U13126 ( .ip1(n11304), .ip2(n12137), .ip3(n11303), .ip4(
        n11302), .op(n11316) );
  mux2_1 U13127 ( .ip1(\ANSWER/mem[0][2][7] ), .ip2(\ANSWER/mem[1][2][7] ), 
        .s(n8833), .op(n11306) );
  mux2_1 U13128 ( .ip1(\ANSWER/mem[2][2][7] ), .ip2(\ANSWER/mem[3][2][7] ), 
        .s(n8833), .op(n11305) );
  mux2_1 U13129 ( .ip1(n11306), .ip2(n11305), .s(n11307), .op(n11311) );
  mux2_1 U13130 ( .ip1(\ANSWER/mem[4][2][7] ), .ip2(\ANSWER/mem[5][2][7] ), 
        .s(n8833), .op(n11309) );
  mux2_1 U13131 ( .ip1(\ANSWER/mem[6][2][7] ), .ip2(\ANSWER/mem[7][2][7] ), 
        .s(n11328), .op(n11308) );
  mux2_1 U13132 ( .ip1(n11309), .ip2(n11308), .s(n11307), .op(n11310) );
  mux2_1 U13133 ( .ip1(n11311), .ip2(n11310), .s(n11979), .op(n11313) );
  mux2_1 U13134 ( .ip1(\ANSWER/mem[8][2][7] ), .ip2(\ANSWER/mem[9][2][7] ), 
        .s(n11328), .op(n11312) );
  mux2_1 U13135 ( .ip1(n11313), .ip2(n11312), .s(n11336), .op(n11314) );
  nand2_1 U13136 ( .ip1(n12147), .ip2(n11314), .op(n11315) );
  nand3_1 U13137 ( .ip1(n11317), .ip2(n11316), .ip3(n11315), .op(n11318) );
  nand2_1 U13138 ( .ip1(n11318), .ip2(n12190), .op(n11342) );
  mux2_1 U13139 ( .ip1(\ANSWER/mem[0][8][7] ), .ip2(\ANSWER/mem[1][8][7] ), 
        .s(n11335), .op(n11320) );
  mux2_1 U13140 ( .ip1(\ANSWER/mem[2][8][7] ), .ip2(\ANSWER/mem[3][8][7] ), 
        .s(n11328), .op(n11319) );
  mux2_1 U13141 ( .ip1(n11320), .ip2(n11319), .s(n11307), .op(n11324) );
  mux2_1 U13142 ( .ip1(\ANSWER/mem[4][8][7] ), .ip2(\ANSWER/mem[5][8][7] ), 
        .s(n11335), .op(n11322) );
  mux2_1 U13143 ( .ip1(\ANSWER/mem[6][8][7] ), .ip2(\ANSWER/mem[7][8][7] ), 
        .s(n11335), .op(n11321) );
  mux2_1 U13144 ( .ip1(n11322), .ip2(n11321), .s(n11008), .op(n11323) );
  mux2_1 U13145 ( .ip1(n11324), .ip2(n11323), .s(n11979), .op(n11326) );
  mux2_1 U13146 ( .ip1(\ANSWER/mem[8][8][7] ), .ip2(\ANSWER/mem[9][8][7] ), 
        .s(n11335), .op(n11325) );
  mux2_1 U13147 ( .ip1(n11326), .ip2(n11325), .s(n11336), .op(n11327) );
  nand2_1 U13148 ( .ip1(n12201), .ip2(n11327), .op(n11341) );
  mux2_1 U13149 ( .ip1(\ANSWER/mem[0][9][7] ), .ip2(\ANSWER/mem[1][9][7] ), 
        .s(n11328), .op(n11330) );
  mux2_1 U13150 ( .ip1(\ANSWER/mem[2][9][7] ), .ip2(\ANSWER/mem[3][9][7] ), 
        .s(n11328), .op(n11329) );
  mux2_1 U13151 ( .ip1(n11330), .ip2(n11329), .s(n11224), .op(n11334) );
  mux2_1 U13152 ( .ip1(\ANSWER/mem[4][9][7] ), .ip2(\ANSWER/mem[5][9][7] ), 
        .s(n11335), .op(n11332) );
  mux2_1 U13153 ( .ip1(\ANSWER/mem[6][9][7] ), .ip2(\ANSWER/mem[7][9][7] ), 
        .s(n11335), .op(n11331) );
  mux2_1 U13154 ( .ip1(n11332), .ip2(n11331), .s(n11224), .op(n11333) );
  mux2_1 U13155 ( .ip1(n11334), .ip2(n11333), .s(n11979), .op(n11338) );
  mux2_1 U13156 ( .ip1(\ANSWER/mem[8][9][7] ), .ip2(\ANSWER/mem[9][9][7] ), 
        .s(n11335), .op(n11337) );
  mux2_1 U13157 ( .ip1(n11338), .ip2(n11337), .s(n11336), .op(n11339) );
  nand2_1 U13158 ( .ip1(n12215), .ip2(n11339), .op(n11340) );
  nand3_1 U13159 ( .ip1(n11342), .ip2(n11341), .ip3(n11340), .op(\ANSWER/N480 ) );
  mux2_1 U13160 ( .ip1(\ANSWER/mem[0][1][8] ), .ip2(\ANSWER/mem[1][1][8] ), 
        .s(n11758), .op(n11344) );
  mux2_1 U13161 ( .ip1(\ANSWER/mem[2][1][8] ), .ip2(\ANSWER/mem[3][1][8] ), 
        .s(n11506), .op(n11343) );
  inv_1 U13162 ( .ip(n12098), .op(n11414) );
  mux2_1 U13163 ( .ip1(n11344), .ip2(n11343), .s(n11414), .op(n11348) );
  mux2_1 U13164 ( .ip1(\ANSWER/mem[4][1][8] ), .ip2(\ANSWER/mem[5][1][8] ), 
        .s(n11070), .op(n11346) );
  mux2_1 U13165 ( .ip1(\ANSWER/mem[6][1][8] ), .ip2(\ANSWER/mem[7][1][8] ), 
        .s(n11164), .op(n11345) );
  mux2_1 U13166 ( .ip1(n11346), .ip2(n11345), .s(n11414), .op(n11347) );
  mux2_1 U13167 ( .ip1(n11348), .ip2(n11347), .s(n11440), .op(n11350) );
  mux2_1 U13168 ( .ip1(\ANSWER/mem[8][1][8] ), .ip2(\ANSWER/mem[9][1][8] ), 
        .s(n11437), .op(n11349) );
  mux2_1 U13169 ( .ip1(n11350), .ip2(n11349), .s(n11552), .op(n11351) );
  nand2_1 U13170 ( .ip1(n12157), .ip2(n11351), .op(n11424) );
  inv_1 U13171 ( .ip(n12109), .op(n11443) );
  mux2_1 U13172 ( .ip1(\ANSWER/mem[0][4][8] ), .ip2(\ANSWER/mem[1][4][8] ), 
        .s(n11443), .op(n11353) );
  mux2_1 U13173 ( .ip1(\ANSWER/mem[2][4][8] ), .ip2(\ANSWER/mem[3][4][8] ), 
        .s(n11443), .op(n11352) );
  mux2_1 U13174 ( .ip1(n11353), .ip2(n11352), .s(n11414), .op(n11357) );
  mux2_1 U13175 ( .ip1(\ANSWER/mem[4][4][8] ), .ip2(\ANSWER/mem[5][4][8] ), 
        .s(n11443), .op(n11355) );
  mux2_1 U13176 ( .ip1(\ANSWER/mem[6][4][8] ), .ip2(\ANSWER/mem[7][4][8] ), 
        .s(n11443), .op(n11354) );
  mux2_1 U13177 ( .ip1(n11355), .ip2(n11354), .s(n11414), .op(n11356) );
  mux2_1 U13178 ( .ip1(n11357), .ip2(n11356), .s(n11440), .op(n11359) );
  mux2_1 U13179 ( .ip1(\ANSWER/mem[8][4][8] ), .ip2(\ANSWER/mem[9][4][8] ), 
        .s(n11443), .op(n11358) );
  mux2_1 U13180 ( .ip1(n11359), .ip2(n11358), .s(n11552), .op(n11411) );
  mux2_1 U13181 ( .ip1(\ANSWER/mem[0][5][8] ), .ip2(\ANSWER/mem[1][5][8] ), 
        .s(n11443), .op(n11361) );
  buf_1 U13182 ( .ip(n11443), .op(n11437) );
  mux2_1 U13183 ( .ip1(\ANSWER/mem[2][5][8] ), .ip2(\ANSWER/mem[3][5][8] ), 
        .s(n11437), .op(n11360) );
  mux2_1 U13184 ( .ip1(n11361), .ip2(n11360), .s(n11414), .op(n11365) );
  mux2_1 U13185 ( .ip1(\ANSWER/mem[4][5][8] ), .ip2(\ANSWER/mem[5][5][8] ), 
        .s(n11437), .op(n11363) );
  mux2_1 U13186 ( .ip1(\ANSWER/mem[6][5][8] ), .ip2(\ANSWER/mem[7][5][8] ), 
        .s(n11437), .op(n11362) );
  mux2_1 U13187 ( .ip1(n11363), .ip2(n11362), .s(n11414), .op(n11364) );
  mux2_1 U13188 ( .ip1(n11365), .ip2(n11364), .s(n11440), .op(n11367) );
  mux2_1 U13189 ( .ip1(\ANSWER/mem[8][5][8] ), .ip2(\ANSWER/mem[9][5][8] ), 
        .s(n11437), .op(n11366) );
  mux2_1 U13190 ( .ip1(n11367), .ip2(n11366), .s(n11552), .op(n11368) );
  and2_1 U13191 ( .ip1(n12127), .ip2(n11368), .op(n11410) );
  mux2_1 U13192 ( .ip1(\ANSWER/mem[0][2][8] ), .ip2(\ANSWER/mem[1][2][8] ), 
        .s(n11164), .op(n11370) );
  mux2_1 U13193 ( .ip1(\ANSWER/mem[2][2][8] ), .ip2(\ANSWER/mem[3][2][8] ), 
        .s(n11758), .op(n11369) );
  mux2_1 U13194 ( .ip1(n11370), .ip2(n11369), .s(n11414), .op(n11374) );
  mux2_1 U13195 ( .ip1(\ANSWER/mem[4][2][8] ), .ip2(\ANSWER/mem[5][2][8] ), 
        .s(n11070), .op(n11372) );
  mux2_1 U13196 ( .ip1(\ANSWER/mem[6][2][8] ), .ip2(\ANSWER/mem[7][2][8] ), 
        .s(n11443), .op(n11371) );
  mux2_1 U13197 ( .ip1(n11372), .ip2(n11371), .s(n11414), .op(n11373) );
  mux2_1 U13198 ( .ip1(n11374), .ip2(n11373), .s(n11440), .op(n11376) );
  mux2_1 U13199 ( .ip1(\ANSWER/mem[8][2][8] ), .ip2(\ANSWER/mem[9][2][8] ), 
        .s(n11443), .op(n11375) );
  mux2_1 U13200 ( .ip1(n11376), .ip2(n11375), .s(n11552), .op(n11377) );
  nand2_1 U13201 ( .ip1(n12147), .ip2(n11377), .op(n11408) );
  mux2_1 U13202 ( .ip1(\ANSWER/mem[0][0][8] ), .ip2(\ANSWER/mem[1][0][8] ), 
        .s(n8833), .op(n11379) );
  mux2_1 U13203 ( .ip1(\ANSWER/mem[2][0][8] ), .ip2(\ANSWER/mem[3][0][8] ), 
        .s(n10816), .op(n11378) );
  mux2_1 U13204 ( .ip1(n11379), .ip2(n11378), .s(n11414), .op(n11383) );
  mux2_1 U13205 ( .ip1(\ANSWER/mem[4][0][8] ), .ip2(\ANSWER/mem[5][0][8] ), 
        .s(n11651), .op(n11381) );
  mux2_1 U13206 ( .ip1(\ANSWER/mem[6][0][8] ), .ip2(\ANSWER/mem[7][0][8] ), 
        .s(n11873), .op(n11380) );
  mux2_1 U13207 ( .ip1(n11381), .ip2(n11380), .s(n11414), .op(n11382) );
  mux2_1 U13208 ( .ip1(n11383), .ip2(n11382), .s(n11440), .op(n11385) );
  mux2_1 U13209 ( .ip1(\ANSWER/mem[8][0][8] ), .ip2(\ANSWER/mem[9][0][8] ), 
        .s(n11113), .op(n11384) );
  mux2_1 U13210 ( .ip1(n11385), .ip2(n11384), .s(n11552), .op(n11386) );
  nand2_1 U13211 ( .ip1(n12108), .ip2(n11386), .op(n11407) );
  mux2_1 U13212 ( .ip1(\ANSWER/mem[0][7][8] ), .ip2(\ANSWER/mem[1][7][8] ), 
        .s(n11437), .op(n11388) );
  mux2_1 U13213 ( .ip1(\ANSWER/mem[2][7][8] ), .ip2(\ANSWER/mem[3][7][8] ), 
        .s(n11437), .op(n11387) );
  mux2_1 U13214 ( .ip1(n11388), .ip2(n11387), .s(n11842), .op(n11392) );
  mux2_1 U13215 ( .ip1(\ANSWER/mem[4][7][8] ), .ip2(\ANSWER/mem[5][7][8] ), 
        .s(n11437), .op(n11390) );
  mux2_1 U13216 ( .ip1(\ANSWER/mem[6][7][8] ), .ip2(\ANSWER/mem[7][7][8] ), 
        .s(n11437), .op(n11389) );
  mux2_1 U13217 ( .ip1(n11390), .ip2(n11389), .s(n11507), .op(n11391) );
  mux2_1 U13218 ( .ip1(n11392), .ip2(n11391), .s(n11440), .op(n11394) );
  mux2_1 U13219 ( .ip1(\ANSWER/mem[8][7][8] ), .ip2(\ANSWER/mem[9][7][8] ), 
        .s(n11443), .op(n11393) );
  mux2_1 U13220 ( .ip1(n11394), .ip2(n11393), .s(n11552), .op(n11395) );
  nand2_1 U13221 ( .ip1(n12186), .ip2(n11395), .op(n11406) );
  mux2_1 U13222 ( .ip1(\ANSWER/mem[0][6][8] ), .ip2(\ANSWER/mem[1][6][8] ), 
        .s(n11437), .op(n11397) );
  mux2_1 U13223 ( .ip1(\ANSWER/mem[2][6][8] ), .ip2(\ANSWER/mem[3][6][8] ), 
        .s(n11437), .op(n11396) );
  mux2_1 U13224 ( .ip1(n11397), .ip2(n11396), .s(n11414), .op(n11401) );
  mux2_1 U13225 ( .ip1(\ANSWER/mem[4][6][8] ), .ip2(\ANSWER/mem[5][6][8] ), 
        .s(n11437), .op(n11399) );
  mux2_1 U13226 ( .ip1(\ANSWER/mem[6][6][8] ), .ip2(\ANSWER/mem[7][6][8] ), 
        .s(n11437), .op(n11398) );
  mux2_1 U13227 ( .ip1(n11399), .ip2(n11398), .s(n11307), .op(n11400) );
  mux2_1 U13228 ( .ip1(n11401), .ip2(n11400), .s(n11440), .op(n11403) );
  mux2_1 U13229 ( .ip1(\ANSWER/mem[8][6][8] ), .ip2(\ANSWER/mem[9][6][8] ), 
        .s(n11437), .op(n11402) );
  mux2_1 U13230 ( .ip1(n11403), .ip2(n11402), .s(n11552), .op(n11404) );
  nand2_1 U13231 ( .ip1(n12168), .ip2(n11404), .op(n11405) );
  nand4_1 U13232 ( .ip1(n11408), .ip2(n11407), .ip3(n11406), .ip4(n11405), 
        .op(n11409) );
  not_ab_or_c_or_d U13233 ( .ip1(n11411), .ip2(n12176), .ip3(n11410), .ip4(
        n11409), .op(n11423) );
  mux2_1 U13234 ( .ip1(\ANSWER/mem[0][3][8] ), .ip2(\ANSWER/mem[1][3][8] ), 
        .s(n11443), .op(n11413) );
  mux2_1 U13235 ( .ip1(\ANSWER/mem[2][3][8] ), .ip2(\ANSWER/mem[3][3][8] ), 
        .s(n11443), .op(n11412) );
  mux2_1 U13236 ( .ip1(n11413), .ip2(n11412), .s(n11414), .op(n11418) );
  mux2_1 U13237 ( .ip1(\ANSWER/mem[4][3][8] ), .ip2(\ANSWER/mem[5][3][8] ), 
        .s(n11443), .op(n11416) );
  mux2_1 U13238 ( .ip1(\ANSWER/mem[6][3][8] ), .ip2(\ANSWER/mem[7][3][8] ), 
        .s(n11443), .op(n11415) );
  mux2_1 U13239 ( .ip1(n11416), .ip2(n11415), .s(n11414), .op(n11417) );
  mux2_1 U13240 ( .ip1(n11418), .ip2(n11417), .s(n11440), .op(n11420) );
  mux2_1 U13241 ( .ip1(\ANSWER/mem[8][3][8] ), .ip2(\ANSWER/mem[9][3][8] ), 
        .s(n11443), .op(n11419) );
  mux2_1 U13242 ( .ip1(n11420), .ip2(n11419), .s(n11552), .op(n11421) );
  nand2_1 U13243 ( .ip1(n12137), .ip2(n11421), .op(n11422) );
  nand3_1 U13244 ( .ip1(n11424), .ip2(n11423), .ip3(n11422), .op(n11425) );
  nand2_1 U13245 ( .ip1(n11425), .ip2(n12190), .op(n11449) );
  mux2_1 U13246 ( .ip1(\ANSWER/mem[0][8][8] ), .ip2(\ANSWER/mem[1][8][8] ), 
        .s(n11443), .op(n11427) );
  mux2_1 U13247 ( .ip1(\ANSWER/mem[2][8][8] ), .ip2(\ANSWER/mem[3][8][8] ), 
        .s(n11437), .op(n11426) );
  mux2_1 U13248 ( .ip1(n11427), .ip2(n11426), .s(n11507), .op(n11431) );
  mux2_1 U13249 ( .ip1(\ANSWER/mem[4][8][8] ), .ip2(\ANSWER/mem[5][8][8] ), 
        .s(n11443), .op(n11429) );
  mux2_1 U13250 ( .ip1(\ANSWER/mem[6][8][8] ), .ip2(\ANSWER/mem[7][8][8] ), 
        .s(n11443), .op(n11428) );
  mux2_1 U13251 ( .ip1(n11429), .ip2(n11428), .s(n11183), .op(n11430) );
  mux2_1 U13252 ( .ip1(n11431), .ip2(n11430), .s(n11440), .op(n11433) );
  mux2_1 U13253 ( .ip1(\ANSWER/mem[8][8][8] ), .ip2(\ANSWER/mem[9][8][8] ), 
        .s(n11443), .op(n11432) );
  mux2_1 U13254 ( .ip1(n11433), .ip2(n11432), .s(n11552), .op(n11434) );
  nand2_1 U13255 ( .ip1(n12201), .ip2(n11434), .op(n11448) );
  mux2_1 U13256 ( .ip1(\ANSWER/mem[0][9][8] ), .ip2(\ANSWER/mem[1][9][8] ), 
        .s(n11443), .op(n11436) );
  mux2_1 U13257 ( .ip1(\ANSWER/mem[2][9][8] ), .ip2(\ANSWER/mem[3][9][8] ), 
        .s(n11437), .op(n11435) );
  mux2_1 U13258 ( .ip1(n11436), .ip2(n11435), .s(n11307), .op(n11442) );
  mux2_1 U13259 ( .ip1(\ANSWER/mem[4][9][8] ), .ip2(\ANSWER/mem[5][9][8] ), 
        .s(n11443), .op(n11439) );
  mux2_1 U13260 ( .ip1(\ANSWER/mem[6][9][8] ), .ip2(\ANSWER/mem[7][9][8] ), 
        .s(n11437), .op(n11438) );
  mux2_1 U13261 ( .ip1(n11439), .ip2(n11438), .s(n11090), .op(n11441) );
  mux2_1 U13262 ( .ip1(n11442), .ip2(n11441), .s(n11440), .op(n11445) );
  mux2_1 U13263 ( .ip1(\ANSWER/mem[8][9][8] ), .ip2(\ANSWER/mem[9][9][8] ), 
        .s(n11443), .op(n11444) );
  mux2_1 U13264 ( .ip1(n11445), .ip2(n11444), .s(n11552), .op(n11446) );
  nand2_1 U13265 ( .ip1(n12215), .ip2(n11446), .op(n11447) );
  nand3_1 U13266 ( .ip1(n11449), .ip2(n11448), .ip3(n11447), .op(\ANSWER/N479 ) );
  inv_1 U13267 ( .ip(n12109), .op(n11551) );
  buf_1 U13268 ( .ip(n11551), .op(n11546) );
  mux2_1 U13269 ( .ip1(\ANSWER/mem[0][5][9] ), .ip2(\ANSWER/mem[1][5][9] ), 
        .s(n11546), .op(n11451) );
  mux2_1 U13270 ( .ip1(\ANSWER/mem[2][5][9] ), .ip2(\ANSWER/mem[3][5][9] ), 
        .s(n11551), .op(n11450) );
  inv_1 U13271 ( .ip(n12098), .op(n11507) );
  mux2_1 U13272 ( .ip1(n11451), .ip2(n11450), .s(n11507), .op(n11456) );
  mux2_1 U13273 ( .ip1(\ANSWER/mem[4][5][9] ), .ip2(\ANSWER/mem[5][5][9] ), 
        .s(n11551), .op(n11453) );
  mux2_1 U13274 ( .ip1(\ANSWER/mem[6][5][9] ), .ip2(\ANSWER/mem[7][5][9] ), 
        .s(n11551), .op(n11452) );
  mux2_1 U13275 ( .ip1(n11453), .ip2(n11452), .s(n11507), .op(n11455) );
  mux2_1 U13276 ( .ip1(n11456), .ip2(n11455), .s(n11440), .op(n11458) );
  mux2_1 U13277 ( .ip1(\ANSWER/mem[8][5][9] ), .ip2(\ANSWER/mem[9][5][9] ), 
        .s(n11551), .op(n11457) );
  mux2_1 U13278 ( .ip1(n11458), .ip2(n11457), .s(n11552), .op(n11459) );
  nand2_1 U13279 ( .ip1(n11459), .ip2(n12127), .op(n11533) );
  inv_1 U13280 ( .ip(n12109), .op(n11506) );
  mux2_1 U13281 ( .ip1(\ANSWER/mem[0][0][9] ), .ip2(\ANSWER/mem[1][0][9] ), 
        .s(n11506), .op(n11461) );
  mux2_1 U13282 ( .ip1(\ANSWER/mem[2][0][9] ), .ip2(\ANSWER/mem[3][0][9] ), 
        .s(n11506), .op(n11460) );
  mux2_1 U13283 ( .ip1(n11461), .ip2(n11460), .s(n11507), .op(n11465) );
  mux2_1 U13284 ( .ip1(\ANSWER/mem[4][0][9] ), .ip2(\ANSWER/mem[5][0][9] ), 
        .s(n11506), .op(n11463) );
  mux2_1 U13285 ( .ip1(\ANSWER/mem[6][0][9] ), .ip2(\ANSWER/mem[7][0][9] ), 
        .s(n11506), .op(n11462) );
  mux2_1 U13286 ( .ip1(n11463), .ip2(n11462), .s(n11507), .op(n11464) );
  mux2_1 U13287 ( .ip1(n11465), .ip2(n11464), .s(n11454), .op(n11467) );
  mux2_1 U13288 ( .ip1(\ANSWER/mem[8][0][9] ), .ip2(\ANSWER/mem[9][0][9] ), 
        .s(n11506), .op(n11466) );
  mux2_1 U13289 ( .ip1(n11467), .ip2(n11466), .s(n11552), .op(n11521) );
  mux2_1 U13290 ( .ip1(\ANSWER/mem[0][3][9] ), .ip2(\ANSWER/mem[1][3][9] ), 
        .s(n11546), .op(n11469) );
  mux2_1 U13291 ( .ip1(\ANSWER/mem[2][3][9] ), .ip2(\ANSWER/mem[3][3][9] ), 
        .s(n11546), .op(n11468) );
  mux2_1 U13292 ( .ip1(n11469), .ip2(n11468), .s(n11507), .op(n11473) );
  mux2_1 U13293 ( .ip1(\ANSWER/mem[4][3][9] ), .ip2(\ANSWER/mem[5][3][9] ), 
        .s(n11546), .op(n11471) );
  mux2_1 U13294 ( .ip1(\ANSWER/mem[6][3][9] ), .ip2(\ANSWER/mem[7][3][9] ), 
        .s(n11546), .op(n11470) );
  mux2_1 U13295 ( .ip1(n11471), .ip2(n11470), .s(n11507), .op(n11472) );
  mux2_1 U13296 ( .ip1(n11473), .ip2(n11472), .s(n11454), .op(n11475) );
  mux2_1 U13297 ( .ip1(\ANSWER/mem[8][3][9] ), .ip2(\ANSWER/mem[9][3][9] ), 
        .s(n11546), .op(n11474) );
  mux2_1 U13298 ( .ip1(n11475), .ip2(n11474), .s(n11552), .op(n11476) );
  and2_1 U13299 ( .ip1(n12137), .ip2(n11476), .op(n11520) );
  mux2_1 U13300 ( .ip1(\ANSWER/mem[0][6][9] ), .ip2(\ANSWER/mem[1][6][9] ), 
        .s(n11551), .op(n11478) );
  mux2_1 U13301 ( .ip1(\ANSWER/mem[2][6][9] ), .ip2(\ANSWER/mem[3][6][9] ), 
        .s(n11551), .op(n11477) );
  mux2_1 U13302 ( .ip1(n11478), .ip2(n11477), .s(n11507), .op(n11482) );
  mux2_1 U13303 ( .ip1(\ANSWER/mem[4][6][9] ), .ip2(\ANSWER/mem[5][6][9] ), 
        .s(n11551), .op(n11480) );
  mux2_1 U13304 ( .ip1(\ANSWER/mem[6][6][9] ), .ip2(\ANSWER/mem[7][6][9] ), 
        .s(n11551), .op(n11479) );
  mux2_1 U13305 ( .ip1(n11480), .ip2(n11479), .s(n11842), .op(n11481) );
  mux2_1 U13306 ( .ip1(n11482), .ip2(n11481), .s(n11454), .op(n11484) );
  mux2_1 U13307 ( .ip1(\ANSWER/mem[8][6][9] ), .ip2(\ANSWER/mem[9][6][9] ), 
        .s(n11551), .op(n11483) );
  mux2_1 U13308 ( .ip1(n11484), .ip2(n11483), .s(n11552), .op(n11485) );
  nand2_1 U13309 ( .ip1(n12168), .ip2(n11485), .op(n11518) );
  mux2_1 U13310 ( .ip1(\ANSWER/mem[0][4][9] ), .ip2(\ANSWER/mem[1][4][9] ), 
        .s(n11546), .op(n11487) );
  mux2_1 U13311 ( .ip1(\ANSWER/mem[2][4][9] ), .ip2(\ANSWER/mem[3][4][9] ), 
        .s(n11546), .op(n11486) );
  mux2_1 U13312 ( .ip1(n11487), .ip2(n11486), .s(n11507), .op(n11491) );
  mux2_1 U13313 ( .ip1(\ANSWER/mem[4][4][9] ), .ip2(\ANSWER/mem[5][4][9] ), 
        .s(n11546), .op(n11489) );
  mux2_1 U13314 ( .ip1(\ANSWER/mem[6][4][9] ), .ip2(\ANSWER/mem[7][4][9] ), 
        .s(n11546), .op(n11488) );
  mux2_1 U13315 ( .ip1(n11489), .ip2(n11488), .s(n11507), .op(n11490) );
  mux2_1 U13316 ( .ip1(n11491), .ip2(n11490), .s(n11440), .op(n11493) );
  mux2_1 U13317 ( .ip1(\ANSWER/mem[8][4][9] ), .ip2(\ANSWER/mem[9][4][9] ), 
        .s(n11546), .op(n11492) );
  mux2_1 U13318 ( .ip1(n11493), .ip2(n11492), .s(n11552), .op(n11494) );
  nand2_1 U13319 ( .ip1(n12176), .ip2(n11494), .op(n11517) );
  mux2_1 U13320 ( .ip1(\ANSWER/mem[0][1][9] ), .ip2(\ANSWER/mem[1][1][9] ), 
        .s(n11506), .op(n11496) );
  mux2_1 U13321 ( .ip1(\ANSWER/mem[2][1][9] ), .ip2(\ANSWER/mem[3][1][9] ), 
        .s(n11506), .op(n11495) );
  mux2_1 U13322 ( .ip1(n11496), .ip2(n11495), .s(n11507), .op(n11500) );
  mux2_1 U13323 ( .ip1(\ANSWER/mem[4][1][9] ), .ip2(\ANSWER/mem[5][1][9] ), 
        .s(n11506), .op(n11498) );
  mux2_1 U13324 ( .ip1(\ANSWER/mem[6][1][9] ), .ip2(\ANSWER/mem[7][1][9] ), 
        .s(n11506), .op(n11497) );
  mux2_1 U13325 ( .ip1(n11498), .ip2(n11497), .s(n11507), .op(n11499) );
  mux2_1 U13326 ( .ip1(n11500), .ip2(n11499), .s(n11440), .op(n11502) );
  mux2_1 U13327 ( .ip1(\ANSWER/mem[8][1][9] ), .ip2(\ANSWER/mem[9][1][9] ), 
        .s(n11506), .op(n11501) );
  mux2_1 U13328 ( .ip1(n11502), .ip2(n11501), .s(n11552), .op(n11503) );
  nand2_1 U13329 ( .ip1(n12157), .ip2(n11503), .op(n11516) );
  mux2_1 U13330 ( .ip1(\ANSWER/mem[0][2][9] ), .ip2(\ANSWER/mem[1][2][9] ), 
        .s(n11506), .op(n11505) );
  mux2_1 U13331 ( .ip1(\ANSWER/mem[2][2][9] ), .ip2(\ANSWER/mem[3][2][9] ), 
        .s(n11506), .op(n11504) );
  mux2_1 U13332 ( .ip1(n11505), .ip2(n11504), .s(n11507), .op(n11511) );
  mux2_1 U13333 ( .ip1(\ANSWER/mem[4][2][9] ), .ip2(\ANSWER/mem[5][2][9] ), 
        .s(n11506), .op(n11509) );
  mux2_1 U13334 ( .ip1(\ANSWER/mem[6][2][9] ), .ip2(\ANSWER/mem[7][2][9] ), 
        .s(n11546), .op(n11508) );
  mux2_1 U13335 ( .ip1(n11509), .ip2(n11508), .s(n11507), .op(n11510) );
  mux2_1 U13336 ( .ip1(n11511), .ip2(n11510), .s(n11440), .op(n11513) );
  mux2_1 U13337 ( .ip1(\ANSWER/mem[8][2][9] ), .ip2(\ANSWER/mem[9][2][9] ), 
        .s(n11546), .op(n11512) );
  mux2_1 U13338 ( .ip1(n11513), .ip2(n11512), .s(n11552), .op(n11514) );
  nand2_1 U13339 ( .ip1(n12147), .ip2(n11514), .op(n11515) );
  nand4_1 U13340 ( .ip1(n11518), .ip2(n11517), .ip3(n11516), .ip4(n11515), 
        .op(n11519) );
  not_ab_or_c_or_d U13341 ( .ip1(n12108), .ip2(n11521), .ip3(n11520), .ip4(
        n11519), .op(n11532) );
  mux2_1 U13342 ( .ip1(\ANSWER/mem[0][7][9] ), .ip2(\ANSWER/mem[1][7][9] ), 
        .s(n11551), .op(n11523) );
  mux2_1 U13343 ( .ip1(\ANSWER/mem[2][7][9] ), .ip2(\ANSWER/mem[3][7][9] ), 
        .s(n11551), .op(n11522) );
  mux2_1 U13344 ( .ip1(n11523), .ip2(n11522), .s(n11183), .op(n11527) );
  mux2_1 U13345 ( .ip1(\ANSWER/mem[4][7][9] ), .ip2(\ANSWER/mem[5][7][9] ), 
        .s(n11551), .op(n11525) );
  mux2_1 U13346 ( .ip1(\ANSWER/mem[6][7][9] ), .ip2(\ANSWER/mem[7][7][9] ), 
        .s(n11551), .op(n11524) );
  mux2_1 U13347 ( .ip1(n11525), .ip2(n11524), .s(n10968), .op(n11526) );
  mux2_1 U13348 ( .ip1(n11527), .ip2(n11526), .s(n11440), .op(n11529) );
  mux2_1 U13349 ( .ip1(\ANSWER/mem[8][7][9] ), .ip2(\ANSWER/mem[9][7][9] ), 
        .s(n11551), .op(n11528) );
  mux2_1 U13350 ( .ip1(n11529), .ip2(n11528), .s(n11552), .op(n11530) );
  nand2_1 U13351 ( .ip1(n12186), .ip2(n11530), .op(n11531) );
  nand3_1 U13352 ( .ip1(n11533), .ip2(n11532), .ip3(n11531), .op(n11534) );
  nand2_1 U13353 ( .ip1(n11534), .ip2(n12190), .op(n11558) );
  mux2_1 U13354 ( .ip1(\ANSWER/mem[0][9][9] ), .ip2(\ANSWER/mem[1][9][9] ), 
        .s(n11546), .op(n11536) );
  mux2_1 U13355 ( .ip1(\ANSWER/mem[2][9][9] ), .ip2(\ANSWER/mem[3][9][9] ), 
        .s(n11551), .op(n11535) );
  mux2_1 U13356 ( .ip1(n11536), .ip2(n11535), .s(n12062), .op(n11540) );
  mux2_1 U13357 ( .ip1(\ANSWER/mem[4][9][9] ), .ip2(\ANSWER/mem[5][9][9] ), 
        .s(n11546), .op(n11538) );
  mux2_1 U13358 ( .ip1(\ANSWER/mem[6][9][9] ), .ip2(\ANSWER/mem[7][9][9] ), 
        .s(n11551), .op(n11537) );
  mux2_1 U13359 ( .ip1(n11538), .ip2(n11537), .s(n11183), .op(n11539) );
  mux2_1 U13360 ( .ip1(n11540), .ip2(n11539), .s(n11454), .op(n11542) );
  mux2_1 U13361 ( .ip1(\ANSWER/mem[8][9][9] ), .ip2(\ANSWER/mem[9][9][9] ), 
        .s(n11551), .op(n11541) );
  mux2_1 U13362 ( .ip1(n11542), .ip2(n11541), .s(n11552), .op(n11543) );
  nand2_1 U13363 ( .ip1(n12215), .ip2(n11543), .op(n11557) );
  mux2_1 U13364 ( .ip1(\ANSWER/mem[0][8][9] ), .ip2(\ANSWER/mem[1][8][9] ), 
        .s(n11551), .op(n11545) );
  mux2_1 U13365 ( .ip1(\ANSWER/mem[2][8][9] ), .ip2(\ANSWER/mem[3][8][9] ), 
        .s(n11551), .op(n11544) );
  mux2_1 U13366 ( .ip1(n11545), .ip2(n11544), .s(n11976), .op(n11550) );
  mux2_1 U13367 ( .ip1(\ANSWER/mem[4][8][9] ), .ip2(\ANSWER/mem[5][8][9] ), 
        .s(n11546), .op(n11548) );
  mux2_1 U13368 ( .ip1(\ANSWER/mem[6][8][9] ), .ip2(\ANSWER/mem[7][8][9] ), 
        .s(n11551), .op(n11547) );
  mux2_1 U13369 ( .ip1(n11548), .ip2(n11547), .s(n11507), .op(n11549) );
  mux2_1 U13370 ( .ip1(n11550), .ip2(n11549), .s(n11440), .op(n11554) );
  mux2_1 U13371 ( .ip1(\ANSWER/mem[8][8][9] ), .ip2(\ANSWER/mem[9][8][9] ), 
        .s(n11551), .op(n11553) );
  mux2_1 U13372 ( .ip1(n11554), .ip2(n11553), .s(n11552), .op(n11555) );
  nand2_1 U13373 ( .ip1(n12201), .ip2(n11555), .op(n11556) );
  nand3_1 U13374 ( .ip1(n11558), .ip2(n11557), .ip3(n11556), .op(\ANSWER/N478 ) );
  inv_1 U13375 ( .ip(n12109), .op(n11659) );
  mux2_1 U13376 ( .ip1(\ANSWER/mem[0][3][10] ), .ip2(\ANSWER/mem[1][3][10] ), 
        .s(n11659), .op(n11560) );
  mux2_1 U13377 ( .ip1(\ANSWER/mem[2][3][10] ), .ip2(\ANSWER/mem[3][3][10] ), 
        .s(n11659), .op(n11559) );
  mux2_1 U13378 ( .ip1(n11560), .ip2(n11559), .s(n10968), .op(n11564) );
  mux2_1 U13379 ( .ip1(\ANSWER/mem[4][3][10] ), .ip2(\ANSWER/mem[5][3][10] ), 
        .s(n11659), .op(n11562) );
  mux2_1 U13380 ( .ip1(\ANSWER/mem[6][3][10] ), .ip2(\ANSWER/mem[7][3][10] ), 
        .s(n11659), .op(n11561) );
  mux2_1 U13381 ( .ip1(n11562), .ip2(n11561), .s(n12158), .op(n11563) );
  mux2_1 U13382 ( .ip1(n11564), .ip2(n11563), .s(n11656), .op(n11567) );
  mux2_1 U13383 ( .ip1(\ANSWER/mem[8][3][10] ), .ip2(\ANSWER/mem[9][3][10] ), 
        .s(n11659), .op(n11566) );
  inv_1 U13384 ( .ip(n11565), .op(n11996) );
  inv_1 U13385 ( .ip(n11996), .op(n11766) );
  mux2_1 U13386 ( .ip1(n11567), .ip2(n11566), .s(n11766), .op(n11568) );
  nand2_1 U13387 ( .ip1(n12137), .ip2(n11568), .op(n11640) );
  mux2_1 U13388 ( .ip1(\ANSWER/mem[0][1][10] ), .ip2(\ANSWER/mem[1][1][10] ), 
        .s(n11506), .op(n11570) );
  mux2_1 U13389 ( .ip1(\ANSWER/mem[2][1][10] ), .ip2(\ANSWER/mem[3][1][10] ), 
        .s(n11873), .op(n11569) );
  mux2_1 U13390 ( .ip1(n11570), .ip2(n11569), .s(n11507), .op(n11574) );
  mux2_1 U13391 ( .ip1(\ANSWER/mem[4][1][10] ), .ip2(\ANSWER/mem[5][1][10] ), 
        .s(n8833), .op(n11572) );
  mux2_1 U13392 ( .ip1(\ANSWER/mem[6][1][10] ), .ip2(\ANSWER/mem[7][1][10] ), 
        .s(n11546), .op(n11571) );
  mux2_1 U13393 ( .ip1(n11572), .ip2(n11571), .s(n11090), .op(n11573) );
  mux2_1 U13394 ( .ip1(n11574), .ip2(n11573), .s(n11656), .op(n11576) );
  mux2_1 U13395 ( .ip1(\ANSWER/mem[8][1][10] ), .ip2(\ANSWER/mem[9][1][10] ), 
        .s(n11070), .op(n11575) );
  mux2_1 U13396 ( .ip1(n11576), .ip2(n11575), .s(n11766), .op(n11628) );
  mux2_1 U13397 ( .ip1(\ANSWER/mem[0][4][10] ), .ip2(\ANSWER/mem[1][4][10] ), 
        .s(n11659), .op(n11578) );
  mux2_1 U13398 ( .ip1(\ANSWER/mem[2][4][10] ), .ip2(\ANSWER/mem[3][4][10] ), 
        .s(n11659), .op(n11577) );
  mux2_1 U13399 ( .ip1(n11578), .ip2(n11577), .s(n11842), .op(n11582) );
  mux2_1 U13400 ( .ip1(\ANSWER/mem[4][4][10] ), .ip2(\ANSWER/mem[5][4][10] ), 
        .s(n11659), .op(n11580) );
  mux2_1 U13401 ( .ip1(\ANSWER/mem[6][4][10] ), .ip2(\ANSWER/mem[7][4][10] ), 
        .s(n11659), .op(n11579) );
  mux2_1 U13402 ( .ip1(n11580), .ip2(n11579), .s(n11307), .op(n11581) );
  mux2_1 U13403 ( .ip1(n11582), .ip2(n11581), .s(n11656), .op(n11584) );
  mux2_1 U13404 ( .ip1(\ANSWER/mem[8][4][10] ), .ip2(\ANSWER/mem[9][4][10] ), 
        .s(n11659), .op(n11583) );
  mux2_1 U13405 ( .ip1(n11584), .ip2(n11583), .s(n11766), .op(n11585) );
  and2_1 U13406 ( .ip1(n12176), .ip2(n11585), .op(n11627) );
  mux2_1 U13407 ( .ip1(\ANSWER/mem[0][5][10] ), .ip2(\ANSWER/mem[1][5][10] ), 
        .s(n11659), .op(n11587) );
  buf_1 U13408 ( .ip(n11659), .op(n11651) );
  mux2_1 U13409 ( .ip1(\ANSWER/mem[2][5][10] ), .ip2(\ANSWER/mem[3][5][10] ), 
        .s(n11651), .op(n11586) );
  mux2_1 U13410 ( .ip1(n11587), .ip2(n11586), .s(n11976), .op(n11591) );
  mux2_1 U13411 ( .ip1(\ANSWER/mem[4][5][10] ), .ip2(\ANSWER/mem[5][5][10] ), 
        .s(n11651), .op(n11589) );
  mux2_1 U13412 ( .ip1(\ANSWER/mem[6][5][10] ), .ip2(\ANSWER/mem[7][5][10] ), 
        .s(n11651), .op(n11588) );
  mux2_1 U13413 ( .ip1(n11589), .ip2(n11588), .s(n12062), .op(n11590) );
  mux2_1 U13414 ( .ip1(n11591), .ip2(n11590), .s(n11656), .op(n11593) );
  mux2_1 U13415 ( .ip1(\ANSWER/mem[8][5][10] ), .ip2(\ANSWER/mem[9][5][10] ), 
        .s(n11651), .op(n11592) );
  mux2_1 U13416 ( .ip1(n11593), .ip2(n11592), .s(n11766), .op(n11594) );
  nand2_1 U13417 ( .ip1(n12127), .ip2(n11594), .op(n11625) );
  mux2_1 U13418 ( .ip1(\ANSWER/mem[0][2][10] ), .ip2(\ANSWER/mem[1][2][10] ), 
        .s(n11506), .op(n11596) );
  mux2_1 U13419 ( .ip1(\ANSWER/mem[2][2][10] ), .ip2(\ANSWER/mem[3][2][10] ), 
        .s(n11437), .op(n11595) );
  mux2_1 U13420 ( .ip1(n11596), .ip2(n11595), .s(n11976), .op(n11600) );
  mux2_1 U13421 ( .ip1(\ANSWER/mem[4][2][10] ), .ip2(\ANSWER/mem[5][2][10] ), 
        .s(n11007), .op(n11598) );
  mux2_1 U13422 ( .ip1(\ANSWER/mem[6][2][10] ), .ip2(\ANSWER/mem[7][2][10] ), 
        .s(n11659), .op(n11597) );
  mux2_1 U13423 ( .ip1(n11598), .ip2(n11597), .s(n11414), .op(n11599) );
  mux2_1 U13424 ( .ip1(n11600), .ip2(n11599), .s(n11656), .op(n11602) );
  mux2_1 U13425 ( .ip1(\ANSWER/mem[8][2][10] ), .ip2(\ANSWER/mem[9][2][10] ), 
        .s(n11659), .op(n11601) );
  mux2_1 U13426 ( .ip1(n11602), .ip2(n11601), .s(n11766), .op(n11603) );
  nand2_1 U13427 ( .ip1(n12147), .ip2(n11603), .op(n11624) );
  mux2_1 U13428 ( .ip1(\ANSWER/mem[0][7][10] ), .ip2(\ANSWER/mem[1][7][10] ), 
        .s(n11651), .op(n11605) );
  mux2_1 U13429 ( .ip1(\ANSWER/mem[2][7][10] ), .ip2(\ANSWER/mem[3][7][10] ), 
        .s(n11651), .op(n11604) );
  mux2_1 U13430 ( .ip1(n11605), .ip2(n11604), .s(n11307), .op(n11609) );
  mux2_1 U13431 ( .ip1(\ANSWER/mem[4][7][10] ), .ip2(\ANSWER/mem[5][7][10] ), 
        .s(n11651), .op(n11607) );
  mux2_1 U13432 ( .ip1(\ANSWER/mem[6][7][10] ), .ip2(\ANSWER/mem[7][7][10] ), 
        .s(n11651), .op(n11606) );
  mux2_1 U13433 ( .ip1(n11607), .ip2(n11606), .s(n11183), .op(n11608) );
  mux2_1 U13434 ( .ip1(n11609), .ip2(n11608), .s(n11656), .op(n11611) );
  mux2_1 U13435 ( .ip1(\ANSWER/mem[8][7][10] ), .ip2(\ANSWER/mem[9][7][10] ), 
        .s(n11659), .op(n11610) );
  mux2_1 U13436 ( .ip1(n11611), .ip2(n11610), .s(n11766), .op(n11612) );
  nand2_1 U13437 ( .ip1(n12186), .ip2(n11612), .op(n11623) );
  mux2_1 U13438 ( .ip1(\ANSWER/mem[0][0][10] ), .ip2(\ANSWER/mem[1][0][10] ), 
        .s(n11070), .op(n11614) );
  mux2_1 U13439 ( .ip1(\ANSWER/mem[2][0][10] ), .ip2(\ANSWER/mem[3][0][10] ), 
        .s(n11975), .op(n11613) );
  mux2_1 U13440 ( .ip1(n11614), .ip2(n11613), .s(n12158), .op(n11618) );
  mux2_1 U13441 ( .ip1(\ANSWER/mem[4][0][10] ), .ip2(\ANSWER/mem[5][0][10] ), 
        .s(n11113), .op(n11616) );
  mux2_1 U13442 ( .ip1(\ANSWER/mem[6][0][10] ), .ip2(\ANSWER/mem[7][0][10] ), 
        .s(n11070), .op(n11615) );
  mux2_1 U13443 ( .ip1(n11616), .ip2(n11615), .s(n11735), .op(n11617) );
  mux2_1 U13444 ( .ip1(n11618), .ip2(n11617), .s(n11656), .op(n11620) );
  mux2_1 U13445 ( .ip1(\ANSWER/mem[8][0][10] ), .ip2(\ANSWER/mem[9][0][10] ), 
        .s(n8833), .op(n11619) );
  mux2_1 U13446 ( .ip1(n11620), .ip2(n11619), .s(n11766), .op(n11621) );
  nand2_1 U13447 ( .ip1(n12108), .ip2(n11621), .op(n11622) );
  nand4_1 U13448 ( .ip1(n11625), .ip2(n11624), .ip3(n11623), .ip4(n11622), 
        .op(n11626) );
  not_ab_or_c_or_d U13449 ( .ip1(n11628), .ip2(n12157), .ip3(n11627), .ip4(
        n11626), .op(n11639) );
  mux2_1 U13450 ( .ip1(\ANSWER/mem[0][6][10] ), .ip2(\ANSWER/mem[1][6][10] ), 
        .s(n11651), .op(n11630) );
  mux2_1 U13451 ( .ip1(\ANSWER/mem[2][6][10] ), .ip2(\ANSWER/mem[3][6][10] ), 
        .s(n11651), .op(n11629) );
  mux2_1 U13452 ( .ip1(n11630), .ip2(n11629), .s(n11183), .op(n11634) );
  mux2_1 U13453 ( .ip1(\ANSWER/mem[4][6][10] ), .ip2(\ANSWER/mem[5][6][10] ), 
        .s(n11651), .op(n11632) );
  mux2_1 U13454 ( .ip1(\ANSWER/mem[6][6][10] ), .ip2(\ANSWER/mem[7][6][10] ), 
        .s(n11651), .op(n11631) );
  mux2_1 U13455 ( .ip1(n11632), .ip2(n11631), .s(n10968), .op(n11633) );
  mux2_1 U13456 ( .ip1(n11634), .ip2(n11633), .s(n11656), .op(n11636) );
  mux2_1 U13457 ( .ip1(\ANSWER/mem[8][6][10] ), .ip2(\ANSWER/mem[9][6][10] ), 
        .s(n11651), .op(n11635) );
  mux2_1 U13458 ( .ip1(n11636), .ip2(n11635), .s(n11766), .op(n11637) );
  nand2_1 U13459 ( .ip1(n12168), .ip2(n11637), .op(n11638) );
  nand3_1 U13460 ( .ip1(n11640), .ip2(n11639), .ip3(n11638), .op(n11641) );
  nand2_1 U13461 ( .ip1(n11641), .ip2(n12190), .op(n11665) );
  mux2_1 U13462 ( .ip1(\ANSWER/mem[0][8][10] ), .ip2(\ANSWER/mem[1][8][10] ), 
        .s(n11659), .op(n11643) );
  mux2_1 U13463 ( .ip1(\ANSWER/mem[2][8][10] ), .ip2(\ANSWER/mem[3][8][10] ), 
        .s(n11651), .op(n11642) );
  mux2_1 U13464 ( .ip1(n11643), .ip2(n11642), .s(n11008), .op(n11647) );
  mux2_1 U13465 ( .ip1(\ANSWER/mem[4][8][10] ), .ip2(\ANSWER/mem[5][8][10] ), 
        .s(n11659), .op(n11645) );
  mux2_1 U13466 ( .ip1(\ANSWER/mem[6][8][10] ), .ip2(\ANSWER/mem[7][8][10] ), 
        .s(n11659), .op(n11644) );
  mux2_1 U13467 ( .ip1(n11645), .ip2(n11644), .s(n11735), .op(n11646) );
  mux2_1 U13468 ( .ip1(n11647), .ip2(n11646), .s(n11656), .op(n11649) );
  mux2_1 U13469 ( .ip1(\ANSWER/mem[8][8][10] ), .ip2(\ANSWER/mem[9][8][10] ), 
        .s(n11659), .op(n11648) );
  mux2_1 U13470 ( .ip1(n11649), .ip2(n11648), .s(n11766), .op(n11650) );
  nand2_1 U13471 ( .ip1(n12201), .ip2(n11650), .op(n11664) );
  mux2_1 U13472 ( .ip1(\ANSWER/mem[0][9][10] ), .ip2(\ANSWER/mem[1][9][10] ), 
        .s(n11651), .op(n11653) );
  mux2_1 U13473 ( .ip1(\ANSWER/mem[2][9][10] ), .ip2(\ANSWER/mem[3][9][10] ), 
        .s(n11651), .op(n11652) );
  mux2_1 U13474 ( .ip1(n11653), .ip2(n11652), .s(n11735), .op(n11658) );
  mux2_1 U13475 ( .ip1(\ANSWER/mem[4][9][10] ), .ip2(\ANSWER/mem[5][9][10] ), 
        .s(n11659), .op(n11655) );
  mux2_1 U13476 ( .ip1(\ANSWER/mem[6][9][10] ), .ip2(\ANSWER/mem[7][9][10] ), 
        .s(n11659), .op(n11654) );
  mux2_1 U13477 ( .ip1(n11655), .ip2(n11654), .s(n11414), .op(n11657) );
  mux2_1 U13478 ( .ip1(n11658), .ip2(n11657), .s(n11656), .op(n11661) );
  mux2_1 U13479 ( .ip1(\ANSWER/mem[8][9][10] ), .ip2(\ANSWER/mem[9][9][10] ), 
        .s(n11659), .op(n11660) );
  mux2_1 U13480 ( .ip1(n11661), .ip2(n11660), .s(n11766), .op(n11662) );
  nand2_1 U13481 ( .ip1(n12215), .ip2(n11662), .op(n11663) );
  nand3_1 U13482 ( .ip1(n11665), .ip2(n11664), .ip3(n11663), .op(\ANSWER/N477 ) );
  mux2_1 U13483 ( .ip1(\ANSWER/mem[0][1][11] ), .ip2(\ANSWER/mem[1][1][11] ), 
        .s(n8833), .op(n11667) );
  mux2_1 U13484 ( .ip1(\ANSWER/mem[2][1][11] ), .ip2(\ANSWER/mem[3][1][11] ), 
        .s(n8833), .op(n11666) );
  inv_1 U13485 ( .ip(n12098), .op(n11735) );
  mux2_1 U13486 ( .ip1(n11667), .ip2(n11666), .s(n11735), .op(n11671) );
  mux2_1 U13487 ( .ip1(\ANSWER/mem[4][1][11] ), .ip2(\ANSWER/mem[5][1][11] ), 
        .s(n11328), .op(n11669) );
  mux2_1 U13488 ( .ip1(\ANSWER/mem[6][1][11] ), .ip2(\ANSWER/mem[7][1][11] ), 
        .s(n12204), .op(n11668) );
  mux2_1 U13489 ( .ip1(n11669), .ip2(n11668), .s(n11735), .op(n11670) );
  mux2_1 U13490 ( .ip1(n11671), .ip2(n11670), .s(n11979), .op(n11673) );
  mux2_1 U13491 ( .ip1(\ANSWER/mem[8][1][11] ), .ip2(\ANSWER/mem[9][1][11] ), 
        .s(n12204), .op(n11672) );
  mux2_1 U13492 ( .ip1(n11673), .ip2(n11672), .s(n11766), .op(n11674) );
  nand2_1 U13493 ( .ip1(n11674), .ip2(n12157), .op(n11747) );
  mux2_1 U13494 ( .ip1(\ANSWER/mem[0][0][11] ), .ip2(\ANSWER/mem[1][0][11] ), 
        .s(n11651), .op(n11676) );
  mux2_1 U13495 ( .ip1(\ANSWER/mem[2][0][11] ), .ip2(\ANSWER/mem[3][0][11] ), 
        .s(n11070), .op(n11675) );
  mux2_1 U13496 ( .ip1(n11676), .ip2(n11675), .s(n11735), .op(n11680) );
  mux2_1 U13497 ( .ip1(\ANSWER/mem[4][0][11] ), .ip2(\ANSWER/mem[5][0][11] ), 
        .s(n12085), .op(n11678) );
  mux2_1 U13498 ( .ip1(\ANSWER/mem[6][0][11] ), .ip2(\ANSWER/mem[7][0][11] ), 
        .s(n11506), .op(n11677) );
  mux2_1 U13499 ( .ip1(n11678), .ip2(n11677), .s(n11735), .op(n11679) );
  mux2_1 U13500 ( .ip1(n11680), .ip2(n11679), .s(n12207), .op(n11682) );
  mux2_1 U13501 ( .ip1(\ANSWER/mem[8][0][11] ), .ip2(\ANSWER/mem[9][0][11] ), 
        .s(n10583), .op(n11681) );
  mux2_1 U13502 ( .ip1(n11682), .ip2(n11681), .s(n11766), .op(n11734) );
  inv_1 U13503 ( .ip(n12109), .op(n11765) );
  buf_1 U13504 ( .ip(n11765), .op(n11758) );
  mux2_1 U13505 ( .ip1(\ANSWER/mem[0][4][11] ), .ip2(\ANSWER/mem[1][4][11] ), 
        .s(n11758), .op(n11684) );
  mux2_1 U13506 ( .ip1(\ANSWER/mem[2][4][11] ), .ip2(\ANSWER/mem[3][4][11] ), 
        .s(n11758), .op(n11683) );
  mux2_1 U13507 ( .ip1(n11684), .ip2(n11683), .s(n11735), .op(n11688) );
  mux2_1 U13508 ( .ip1(\ANSWER/mem[4][4][11] ), .ip2(\ANSWER/mem[5][4][11] ), 
        .s(n11758), .op(n11686) );
  mux2_1 U13509 ( .ip1(\ANSWER/mem[6][4][11] ), .ip2(\ANSWER/mem[7][4][11] ), 
        .s(n11758), .op(n11685) );
  mux2_1 U13510 ( .ip1(n11686), .ip2(n11685), .s(n11735), .op(n11687) );
  mux2_1 U13511 ( .ip1(n11688), .ip2(n11687), .s(n11454), .op(n11690) );
  mux2_1 U13512 ( .ip1(\ANSWER/mem[8][4][11] ), .ip2(\ANSWER/mem[9][4][11] ), 
        .s(n11758), .op(n11689) );
  mux2_1 U13513 ( .ip1(n11690), .ip2(n11689), .s(n11766), .op(n11691) );
  and2_1 U13514 ( .ip1(n12176), .ip2(n11691), .op(n11733) );
  mux2_1 U13515 ( .ip1(\ANSWER/mem[0][7][11] ), .ip2(\ANSWER/mem[1][7][11] ), 
        .s(n11765), .op(n11693) );
  mux2_1 U13516 ( .ip1(\ANSWER/mem[2][7][11] ), .ip2(\ANSWER/mem[3][7][11] ), 
        .s(n11765), .op(n11692) );
  mux2_1 U13517 ( .ip1(n11693), .ip2(n11692), .s(n12158), .op(n11697) );
  mux2_1 U13518 ( .ip1(\ANSWER/mem[4][7][11] ), .ip2(\ANSWER/mem[5][7][11] ), 
        .s(n11765), .op(n11695) );
  mux2_1 U13519 ( .ip1(\ANSWER/mem[6][7][11] ), .ip2(\ANSWER/mem[7][7][11] ), 
        .s(n11765), .op(n11694) );
  mux2_1 U13520 ( .ip1(n11695), .ip2(n11694), .s(n11950), .op(n11696) );
  mux2_1 U13521 ( .ip1(n11697), .ip2(n11696), .s(n8821), .op(n11699) );
  mux2_1 U13522 ( .ip1(\ANSWER/mem[8][7][11] ), .ip2(\ANSWER/mem[9][7][11] ), 
        .s(n11765), .op(n11698) );
  mux2_1 U13523 ( .ip1(n11699), .ip2(n11698), .s(n11766), .op(n11700) );
  nand2_1 U13524 ( .ip1(n12186), .ip2(n11700), .op(n11731) );
  mux2_1 U13525 ( .ip1(\ANSWER/mem[0][5][11] ), .ip2(\ANSWER/mem[1][5][11] ), 
        .s(n11758), .op(n11702) );
  mux2_1 U13526 ( .ip1(\ANSWER/mem[2][5][11] ), .ip2(\ANSWER/mem[3][5][11] ), 
        .s(n11765), .op(n11701) );
  mux2_1 U13527 ( .ip1(n11702), .ip2(n11701), .s(n11735), .op(n11706) );
  mux2_1 U13528 ( .ip1(\ANSWER/mem[4][5][11] ), .ip2(\ANSWER/mem[5][5][11] ), 
        .s(n11765), .op(n11704) );
  mux2_1 U13529 ( .ip1(\ANSWER/mem[6][5][11] ), .ip2(\ANSWER/mem[7][5][11] ), 
        .s(n11765), .op(n11703) );
  mux2_1 U13530 ( .ip1(n11704), .ip2(n11703), .s(n11735), .op(n11705) );
  mux2_1 U13531 ( .ip1(n11706), .ip2(n11705), .s(n12207), .op(n11708) );
  mux2_1 U13532 ( .ip1(\ANSWER/mem[8][5][11] ), .ip2(\ANSWER/mem[9][5][11] ), 
        .s(n11765), .op(n11707) );
  mux2_1 U13533 ( .ip1(n11708), .ip2(n11707), .s(n11766), .op(n11709) );
  nand2_1 U13534 ( .ip1(n12127), .ip2(n11709), .op(n11730) );
  mux2_1 U13535 ( .ip1(\ANSWER/mem[0][2][11] ), .ip2(\ANSWER/mem[1][2][11] ), 
        .s(n11164), .op(n11711) );
  mux2_1 U13536 ( .ip1(\ANSWER/mem[2][2][11] ), .ip2(\ANSWER/mem[3][2][11] ), 
        .s(n11975), .op(n11710) );
  mux2_1 U13537 ( .ip1(n11711), .ip2(n11710), .s(n11735), .op(n11715) );
  mux2_1 U13538 ( .ip1(\ANSWER/mem[4][2][11] ), .ip2(\ANSWER/mem[5][2][11] ), 
        .s(n12204), .op(n11713) );
  mux2_1 U13539 ( .ip1(\ANSWER/mem[6][2][11] ), .ip2(\ANSWER/mem[7][2][11] ), 
        .s(n11758), .op(n11712) );
  mux2_1 U13540 ( .ip1(n11713), .ip2(n11712), .s(n11735), .op(n11714) );
  mux2_1 U13541 ( .ip1(n11715), .ip2(n11714), .s(n11937), .op(n11717) );
  mux2_1 U13542 ( .ip1(\ANSWER/mem[8][2][11] ), .ip2(\ANSWER/mem[9][2][11] ), 
        .s(n11758), .op(n11716) );
  mux2_1 U13543 ( .ip1(n11717), .ip2(n11716), .s(n11766), .op(n11718) );
  nand2_1 U13544 ( .ip1(n12147), .ip2(n11718), .op(n11729) );
  mux2_1 U13545 ( .ip1(\ANSWER/mem[0][3][11] ), .ip2(\ANSWER/mem[1][3][11] ), 
        .s(n11758), .op(n11720) );
  mux2_1 U13546 ( .ip1(\ANSWER/mem[2][3][11] ), .ip2(\ANSWER/mem[3][3][11] ), 
        .s(n11758), .op(n11719) );
  mux2_1 U13547 ( .ip1(n11720), .ip2(n11719), .s(n11735), .op(n11724) );
  mux2_1 U13548 ( .ip1(\ANSWER/mem[4][3][11] ), .ip2(\ANSWER/mem[5][3][11] ), 
        .s(n11758), .op(n11722) );
  mux2_1 U13549 ( .ip1(\ANSWER/mem[6][3][11] ), .ip2(\ANSWER/mem[7][3][11] ), 
        .s(n11758), .op(n11721) );
  mux2_1 U13550 ( .ip1(n11722), .ip2(n11721), .s(n11735), .op(n11723) );
  mux2_1 U13551 ( .ip1(n11724), .ip2(n11723), .s(n11454), .op(n11726) );
  mux2_1 U13552 ( .ip1(\ANSWER/mem[8][3][11] ), .ip2(\ANSWER/mem[9][3][11] ), 
        .s(n11758), .op(n11725) );
  mux2_1 U13553 ( .ip1(n11726), .ip2(n11725), .s(n11766), .op(n11727) );
  nand2_1 U13554 ( .ip1(n12137), .ip2(n11727), .op(n11728) );
  nand4_1 U13555 ( .ip1(n11731), .ip2(n11730), .ip3(n11729), .ip4(n11728), 
        .op(n11732) );
  not_ab_or_c_or_d U13556 ( .ip1(n11734), .ip2(n12108), .ip3(n11733), .ip4(
        n11732), .op(n11746) );
  mux2_1 U13557 ( .ip1(\ANSWER/mem[0][6][11] ), .ip2(\ANSWER/mem[1][6][11] ), 
        .s(n11765), .op(n11737) );
  mux2_1 U13558 ( .ip1(\ANSWER/mem[2][6][11] ), .ip2(\ANSWER/mem[3][6][11] ), 
        .s(n11765), .op(n11736) );
  mux2_1 U13559 ( .ip1(n11737), .ip2(n11736), .s(n11735), .op(n11741) );
  mux2_1 U13560 ( .ip1(\ANSWER/mem[4][6][11] ), .ip2(\ANSWER/mem[5][6][11] ), 
        .s(n11765), .op(n11739) );
  mux2_1 U13561 ( .ip1(\ANSWER/mem[6][6][11] ), .ip2(\ANSWER/mem[7][6][11] ), 
        .s(n11765), .op(n11738) );
  mux2_1 U13562 ( .ip1(n11739), .ip2(n11738), .s(n11735), .op(n11740) );
  mux2_1 U13563 ( .ip1(n11741), .ip2(n11740), .s(n12088), .op(n11743) );
  mux2_1 U13564 ( .ip1(\ANSWER/mem[8][6][11] ), .ip2(\ANSWER/mem[9][6][11] ), 
        .s(n11765), .op(n11742) );
  mux2_1 U13565 ( .ip1(n11743), .ip2(n11742), .s(n11766), .op(n11744) );
  nand2_1 U13566 ( .ip1(n12168), .ip2(n11744), .op(n11745) );
  nand3_1 U13567 ( .ip1(n11747), .ip2(n11746), .ip3(n11745), .op(n11748) );
  nand2_1 U13568 ( .ip1(n11748), .ip2(n12190), .op(n11772) );
  mux2_1 U13569 ( .ip1(\ANSWER/mem[0][8][11] ), .ip2(\ANSWER/mem[1][8][11] ), 
        .s(n11765), .op(n11750) );
  mux2_1 U13570 ( .ip1(\ANSWER/mem[2][8][11] ), .ip2(\ANSWER/mem[3][8][11] ), 
        .s(n11758), .op(n11749) );
  mux2_1 U13571 ( .ip1(n11750), .ip2(n11749), .s(n11008), .op(n11754) );
  mux2_1 U13572 ( .ip1(\ANSWER/mem[4][8][11] ), .ip2(\ANSWER/mem[5][8][11] ), 
        .s(n11765), .op(n11752) );
  mux2_1 U13573 ( .ip1(\ANSWER/mem[6][8][11] ), .ip2(\ANSWER/mem[7][8][11] ), 
        .s(n11765), .op(n11751) );
  mux2_1 U13574 ( .ip1(n11752), .ip2(n11751), .s(n11976), .op(n11753) );
  mux2_1 U13575 ( .ip1(n11754), .ip2(n11753), .s(n12088), .op(n11756) );
  mux2_1 U13576 ( .ip1(\ANSWER/mem[8][8][11] ), .ip2(\ANSWER/mem[9][8][11] ), 
        .s(n11765), .op(n11755) );
  mux2_1 U13577 ( .ip1(n11756), .ip2(n11755), .s(n11766), .op(n11757) );
  nand2_1 U13578 ( .ip1(n12201), .ip2(n11757), .op(n11771) );
  mux2_1 U13579 ( .ip1(\ANSWER/mem[0][9][11] ), .ip2(\ANSWER/mem[1][9][11] ), 
        .s(n11758), .op(n11760) );
  mux2_1 U13580 ( .ip1(\ANSWER/mem[2][9][11] ), .ip2(\ANSWER/mem[3][9][11] ), 
        .s(n11758), .op(n11759) );
  mux2_1 U13581 ( .ip1(n11760), .ip2(n11759), .s(n12062), .op(n11764) );
  mux2_1 U13582 ( .ip1(\ANSWER/mem[4][9][11] ), .ip2(\ANSWER/mem[5][9][11] ), 
        .s(n11765), .op(n11762) );
  mux2_1 U13583 ( .ip1(\ANSWER/mem[6][9][11] ), .ip2(\ANSWER/mem[7][9][11] ), 
        .s(n11765), .op(n11761) );
  mux2_1 U13584 ( .ip1(n11762), .ip2(n11761), .s(n11842), .op(n11763) );
  mux2_1 U13585 ( .ip1(n11764), .ip2(n11763), .s(n8821), .op(n11768) );
  mux2_1 U13586 ( .ip1(\ANSWER/mem[8][9][11] ), .ip2(\ANSWER/mem[9][9][11] ), 
        .s(n11765), .op(n11767) );
  mux2_1 U13587 ( .ip1(n11768), .ip2(n11767), .s(n11766), .op(n11769) );
  nand2_1 U13588 ( .ip1(n12215), .ip2(n11769), .op(n11770) );
  nand3_1 U13589 ( .ip1(n11772), .ip2(n11771), .ip3(n11770), .op(\ANSWER/N476 ) );
  inv_1 U13590 ( .ip(n12109), .op(n11867) );
  buf_1 U13591 ( .ip(n11867), .op(n11873) );
  mux2_1 U13592 ( .ip1(\ANSWER/mem[0][4][12] ), .ip2(\ANSWER/mem[1][4][12] ), 
        .s(n11873), .op(n11774) );
  mux2_1 U13593 ( .ip1(\ANSWER/mem[2][4][12] ), .ip2(\ANSWER/mem[3][4][12] ), 
        .s(n11873), .op(n11773) );
  inv_1 U13594 ( .ip(n12098), .op(n11842) );
  mux2_1 U13595 ( .ip1(n11774), .ip2(n11773), .s(n11842), .op(n11778) );
  mux2_1 U13596 ( .ip1(\ANSWER/mem[4][4][12] ), .ip2(\ANSWER/mem[5][4][12] ), 
        .s(n11873), .op(n11776) );
  mux2_1 U13597 ( .ip1(\ANSWER/mem[6][4][12] ), .ip2(\ANSWER/mem[7][4][12] ), 
        .s(n11873), .op(n11775) );
  mux2_1 U13598 ( .ip1(n11776), .ip2(n11775), .s(n11842), .op(n11777) );
  mux2_1 U13599 ( .ip1(n11778), .ip2(n11777), .s(n11454), .op(n11780) );
  mux2_1 U13600 ( .ip1(\ANSWER/mem[8][4][12] ), .ip2(\ANSWER/mem[9][4][12] ), 
        .s(n11873), .op(n11779) );
  inv_1 U13601 ( .ip(n11996), .op(n11983) );
  mux2_1 U13602 ( .ip1(n11780), .ip2(n11779), .s(n11983), .op(n11781) );
  nand2_1 U13603 ( .ip1(n12176), .ip2(n11781), .op(n11854) );
  mux2_1 U13604 ( .ip1(\ANSWER/mem[0][5][12] ), .ip2(\ANSWER/mem[1][5][12] ), 
        .s(n11873), .op(n11783) );
  mux2_1 U13605 ( .ip1(\ANSWER/mem[2][5][12] ), .ip2(\ANSWER/mem[3][5][12] ), 
        .s(n11867), .op(n11782) );
  mux2_1 U13606 ( .ip1(n11783), .ip2(n11782), .s(n11842), .op(n11787) );
  mux2_1 U13607 ( .ip1(\ANSWER/mem[4][5][12] ), .ip2(\ANSWER/mem[5][5][12] ), 
        .s(n11867), .op(n11785) );
  mux2_1 U13608 ( .ip1(\ANSWER/mem[6][5][12] ), .ip2(\ANSWER/mem[7][5][12] ), 
        .s(n11867), .op(n11784) );
  mux2_1 U13609 ( .ip1(n11785), .ip2(n11784), .s(n11842), .op(n11786) );
  mux2_1 U13610 ( .ip1(n11787), .ip2(n11786), .s(n11440), .op(n11789) );
  mux2_1 U13611 ( .ip1(\ANSWER/mem[8][5][12] ), .ip2(\ANSWER/mem[9][5][12] ), 
        .s(n11867), .op(n11788) );
  mux2_1 U13612 ( .ip1(n11789), .ip2(n11788), .s(n11983), .op(n11841) );
  mux2_1 U13613 ( .ip1(\ANSWER/mem[0][7][12] ), .ip2(\ANSWER/mem[1][7][12] ), 
        .s(n11873), .op(n11791) );
  mux2_1 U13614 ( .ip1(\ANSWER/mem[2][7][12] ), .ip2(\ANSWER/mem[3][7][12] ), 
        .s(n11867), .op(n11790) );
  mux2_1 U13615 ( .ip1(n11791), .ip2(n11790), .s(n11868), .op(n11795) );
  mux2_1 U13616 ( .ip1(\ANSWER/mem[4][7][12] ), .ip2(\ANSWER/mem[5][7][12] ), 
        .s(n11867), .op(n11793) );
  mux2_1 U13617 ( .ip1(\ANSWER/mem[6][7][12] ), .ip2(\ANSWER/mem[7][7][12] ), 
        .s(n11867), .op(n11792) );
  mux2_1 U13618 ( .ip1(n11793), .ip2(n11792), .s(n11868), .op(n11794) );
  mux2_1 U13619 ( .ip1(n11795), .ip2(n11794), .s(n11440), .op(n11797) );
  mux2_1 U13620 ( .ip1(\ANSWER/mem[8][7][12] ), .ip2(\ANSWER/mem[9][7][12] ), 
        .s(n11867), .op(n11796) );
  mux2_1 U13621 ( .ip1(n11797), .ip2(n11796), .s(n11983), .op(n11798) );
  and2_1 U13622 ( .ip1(n12186), .ip2(n11798), .op(n11840) );
  mux2_1 U13623 ( .ip1(\ANSWER/mem[0][0][12] ), .ip2(\ANSWER/mem[1][0][12] ), 
        .s(n10816), .op(n11800) );
  mux2_1 U13624 ( .ip1(\ANSWER/mem[2][0][12] ), .ip2(\ANSWER/mem[3][0][12] ), 
        .s(n10583), .op(n11799) );
  mux2_1 U13625 ( .ip1(n11800), .ip2(n11799), .s(n11842), .op(n11804) );
  mux2_1 U13626 ( .ip1(\ANSWER/mem[4][0][12] ), .ip2(\ANSWER/mem[5][0][12] ), 
        .s(n11223), .op(n11802) );
  mux2_1 U13627 ( .ip1(\ANSWER/mem[6][0][12] ), .ip2(\ANSWER/mem[7][0][12] ), 
        .s(n11437), .op(n11801) );
  mux2_1 U13628 ( .ip1(n11802), .ip2(n11801), .s(n11842), .op(n11803) );
  mux2_1 U13629 ( .ip1(n11804), .ip2(n11803), .s(n11440), .op(n11806) );
  mux2_1 U13630 ( .ip1(\ANSWER/mem[8][0][12] ), .ip2(\ANSWER/mem[9][0][12] ), 
        .s(n11328), .op(n11805) );
  mux2_1 U13631 ( .ip1(n11806), .ip2(n11805), .s(n11983), .op(n11807) );
  nand2_1 U13632 ( .ip1(n12108), .ip2(n11807), .op(n11838) );
  mux2_1 U13633 ( .ip1(\ANSWER/mem[0][1][12] ), .ip2(\ANSWER/mem[1][1][12] ), 
        .s(n11758), .op(n11809) );
  mux2_1 U13634 ( .ip1(\ANSWER/mem[2][1][12] ), .ip2(\ANSWER/mem[3][1][12] ), 
        .s(n12204), .op(n11808) );
  mux2_1 U13635 ( .ip1(n11809), .ip2(n11808), .s(n11842), .op(n11813) );
  mux2_1 U13636 ( .ip1(\ANSWER/mem[4][1][12] ), .ip2(\ANSWER/mem[5][1][12] ), 
        .s(n11328), .op(n11811) );
  mux2_1 U13637 ( .ip1(\ANSWER/mem[6][1][12] ), .ip2(\ANSWER/mem[7][1][12] ), 
        .s(n11975), .op(n11810) );
  mux2_1 U13638 ( .ip1(n11811), .ip2(n11810), .s(n11842), .op(n11812) );
  mux2_1 U13639 ( .ip1(n11813), .ip2(n11812), .s(n11454), .op(n11815) );
  mux2_1 U13640 ( .ip1(\ANSWER/mem[8][1][12] ), .ip2(\ANSWER/mem[9][1][12] ), 
        .s(n11546), .op(n11814) );
  mux2_1 U13641 ( .ip1(n11815), .ip2(n11814), .s(n11983), .op(n11816) );
  nand2_1 U13642 ( .ip1(n12157), .ip2(n11816), .op(n11837) );
  mux2_1 U13643 ( .ip1(\ANSWER/mem[0][2][12] ), .ip2(\ANSWER/mem[1][2][12] ), 
        .s(n11873), .op(n11818) );
  mux2_1 U13644 ( .ip1(\ANSWER/mem[2][2][12] ), .ip2(\ANSWER/mem[3][2][12] ), 
        .s(n11437), .op(n11817) );
  mux2_1 U13645 ( .ip1(n11818), .ip2(n11817), .s(n11842), .op(n11822) );
  mux2_1 U13646 ( .ip1(\ANSWER/mem[4][2][12] ), .ip2(\ANSWER/mem[5][2][12] ), 
        .s(n11975), .op(n11820) );
  mux2_1 U13647 ( .ip1(\ANSWER/mem[6][2][12] ), .ip2(\ANSWER/mem[7][2][12] ), 
        .s(n11873), .op(n11819) );
  mux2_1 U13648 ( .ip1(n11820), .ip2(n11819), .s(n11842), .op(n11821) );
  mux2_1 U13649 ( .ip1(n11822), .ip2(n11821), .s(n11440), .op(n11824) );
  mux2_1 U13650 ( .ip1(\ANSWER/mem[8][2][12] ), .ip2(\ANSWER/mem[9][2][12] ), 
        .s(n11873), .op(n11823) );
  mux2_1 U13651 ( .ip1(n11824), .ip2(n11823), .s(n11983), .op(n11825) );
  nand2_1 U13652 ( .ip1(n12147), .ip2(n11825), .op(n11836) );
  mux2_1 U13653 ( .ip1(\ANSWER/mem[0][3][12] ), .ip2(\ANSWER/mem[1][3][12] ), 
        .s(n11873), .op(n11827) );
  mux2_1 U13654 ( .ip1(\ANSWER/mem[2][3][12] ), .ip2(\ANSWER/mem[3][3][12] ), 
        .s(n11873), .op(n11826) );
  mux2_1 U13655 ( .ip1(n11827), .ip2(n11826), .s(n11842), .op(n11831) );
  mux2_1 U13656 ( .ip1(\ANSWER/mem[4][3][12] ), .ip2(\ANSWER/mem[5][3][12] ), 
        .s(n11873), .op(n11829) );
  mux2_1 U13657 ( .ip1(\ANSWER/mem[6][3][12] ), .ip2(\ANSWER/mem[7][3][12] ), 
        .s(n11873), .op(n11828) );
  mux2_1 U13658 ( .ip1(n11829), .ip2(n11828), .s(n11842), .op(n11830) );
  mux2_1 U13659 ( .ip1(n11831), .ip2(n11830), .s(n11440), .op(n11833) );
  mux2_1 U13660 ( .ip1(\ANSWER/mem[8][3][12] ), .ip2(\ANSWER/mem[9][3][12] ), 
        .s(n11873), .op(n11832) );
  mux2_1 U13661 ( .ip1(n11833), .ip2(n11832), .s(n11983), .op(n11834) );
  nand2_1 U13662 ( .ip1(n12137), .ip2(n11834), .op(n11835) );
  nand4_1 U13663 ( .ip1(n11838), .ip2(n11837), .ip3(n11836), .ip4(n11835), 
        .op(n11839) );
  not_ab_or_c_or_d U13664 ( .ip1(n11841), .ip2(n12127), .ip3(n11840), .ip4(
        n11839), .op(n11853) );
  mux2_1 U13665 ( .ip1(\ANSWER/mem[0][6][12] ), .ip2(\ANSWER/mem[1][6][12] ), 
        .s(n11867), .op(n11844) );
  mux2_1 U13666 ( .ip1(\ANSWER/mem[2][6][12] ), .ip2(\ANSWER/mem[3][6][12] ), 
        .s(n11867), .op(n11843) );
  mux2_1 U13667 ( .ip1(n11844), .ip2(n11843), .s(n11842), .op(n11848) );
  mux2_1 U13668 ( .ip1(\ANSWER/mem[4][6][12] ), .ip2(\ANSWER/mem[5][6][12] ), 
        .s(n11867), .op(n11846) );
  mux2_1 U13669 ( .ip1(\ANSWER/mem[6][6][12] ), .ip2(\ANSWER/mem[7][6][12] ), 
        .s(n11867), .op(n11845) );
  mux2_1 U13670 ( .ip1(n11846), .ip2(n11845), .s(n11868), .op(n11847) );
  mux2_1 U13671 ( .ip1(n11848), .ip2(n11847), .s(n11454), .op(n11850) );
  mux2_1 U13672 ( .ip1(\ANSWER/mem[8][6][12] ), .ip2(\ANSWER/mem[9][6][12] ), 
        .s(n11867), .op(n11849) );
  mux2_1 U13673 ( .ip1(n11850), .ip2(n11849), .s(n11983), .op(n11851) );
  nand2_1 U13674 ( .ip1(n12168), .ip2(n11851), .op(n11852) );
  nand3_1 U13675 ( .ip1(n11854), .ip2(n11853), .ip3(n11852), .op(n11855) );
  nand2_1 U13676 ( .ip1(n11855), .ip2(n12190), .op(n11879) );
  mux2_1 U13677 ( .ip1(\ANSWER/mem[0][9][12] ), .ip2(\ANSWER/mem[1][9][12] ), 
        .s(n11867), .op(n11857) );
  mux2_1 U13678 ( .ip1(\ANSWER/mem[2][9][12] ), .ip2(\ANSWER/mem[3][9][12] ), 
        .s(n11867), .op(n11856) );
  mux2_1 U13679 ( .ip1(n11857), .ip2(n11856), .s(n11868), .op(n11861) );
  mux2_1 U13680 ( .ip1(\ANSWER/mem[4][9][12] ), .ip2(\ANSWER/mem[5][9][12] ), 
        .s(n11867), .op(n11859) );
  mux2_1 U13681 ( .ip1(\ANSWER/mem[6][9][12] ), .ip2(\ANSWER/mem[7][9][12] ), 
        .s(n11867), .op(n11858) );
  mux2_1 U13682 ( .ip1(n11859), .ip2(n11858), .s(n11868), .op(n11860) );
  mux2_1 U13683 ( .ip1(n11861), .ip2(n11860), .s(n11656), .op(n11863) );
  mux2_1 U13684 ( .ip1(\ANSWER/mem[8][9][12] ), .ip2(\ANSWER/mem[9][9][12] ), 
        .s(n11873), .op(n11862) );
  mux2_1 U13685 ( .ip1(n11863), .ip2(n11862), .s(n11983), .op(n11864) );
  nand2_1 U13686 ( .ip1(n12215), .ip2(n11864), .op(n11878) );
  mux2_1 U13687 ( .ip1(\ANSWER/mem[0][8][12] ), .ip2(\ANSWER/mem[1][8][12] ), 
        .s(n11867), .op(n11866) );
  mux2_1 U13688 ( .ip1(\ANSWER/mem[2][8][12] ), .ip2(\ANSWER/mem[3][8][12] ), 
        .s(n11867), .op(n11865) );
  mux2_1 U13689 ( .ip1(n11866), .ip2(n11865), .s(n11868), .op(n11872) );
  mux2_1 U13690 ( .ip1(\ANSWER/mem[4][8][12] ), .ip2(\ANSWER/mem[5][8][12] ), 
        .s(n11867), .op(n11870) );
  mux2_1 U13691 ( .ip1(\ANSWER/mem[6][8][12] ), .ip2(\ANSWER/mem[7][8][12] ), 
        .s(n11867), .op(n11869) );
  mux2_1 U13692 ( .ip1(n11870), .ip2(n11869), .s(n11868), .op(n11871) );
  mux2_1 U13693 ( .ip1(n11872), .ip2(n11871), .s(n11454), .op(n11875) );
  mux2_1 U13694 ( .ip1(\ANSWER/mem[8][8][12] ), .ip2(\ANSWER/mem[9][8][12] ), 
        .s(n11873), .op(n11874) );
  mux2_1 U13695 ( .ip1(n11875), .ip2(n11874), .s(n11983), .op(n11876) );
  nand2_1 U13696 ( .ip1(n12201), .ip2(n11876), .op(n11877) );
  nand3_1 U13697 ( .ip1(n11879), .ip2(n11878), .ip3(n11877), .op(\ANSWER/N475 ) );
  mux2_1 U13698 ( .ip1(\ANSWER/mem[0][1][13] ), .ip2(\ANSWER/mem[1][1][13] ), 
        .s(n11328), .op(n11881) );
  mux2_1 U13699 ( .ip1(\ANSWER/mem[2][1][13] ), .ip2(\ANSWER/mem[3][1][13] ), 
        .s(n12204), .op(n11880) );
  inv_1 U13700 ( .ip(n12098), .op(n11950) );
  mux2_1 U13701 ( .ip1(n11881), .ip2(n11880), .s(n11950), .op(n11885) );
  mux2_1 U13702 ( .ip1(\ANSWER/mem[4][1][13] ), .ip2(\ANSWER/mem[5][1][13] ), 
        .s(n11007), .op(n11883) );
  mux2_1 U13703 ( .ip1(\ANSWER/mem[6][1][13] ), .ip2(\ANSWER/mem[7][1][13] ), 
        .s(n11013), .op(n11882) );
  mux2_1 U13704 ( .ip1(n11883), .ip2(n11882), .s(n11950), .op(n11884) );
  mux2_1 U13705 ( .ip1(n11885), .ip2(n11884), .s(n11979), .op(n11887) );
  mux2_1 U13706 ( .ip1(\ANSWER/mem[8][1][13] ), .ip2(\ANSWER/mem[9][1][13] ), 
        .s(n11651), .op(n11886) );
  mux2_1 U13707 ( .ip1(n11887), .ip2(n11886), .s(n11983), .op(n11888) );
  nand2_1 U13708 ( .ip1(n12157), .ip2(n11888), .op(n11962) );
  inv_1 U13709 ( .ip(n12109), .op(n11982) );
  buf_1 U13710 ( .ip(n11982), .op(n11975) );
  mux2_1 U13711 ( .ip1(\ANSWER/mem[0][3][13] ), .ip2(\ANSWER/mem[1][3][13] ), 
        .s(n11975), .op(n11890) );
  mux2_1 U13712 ( .ip1(\ANSWER/mem[2][3][13] ), .ip2(\ANSWER/mem[3][3][13] ), 
        .s(n11975), .op(n11889) );
  mux2_1 U13713 ( .ip1(n11890), .ip2(n11889), .s(n11950), .op(n11894) );
  mux2_1 U13714 ( .ip1(\ANSWER/mem[4][3][13] ), .ip2(\ANSWER/mem[5][3][13] ), 
        .s(n11975), .op(n11892) );
  mux2_1 U13715 ( .ip1(\ANSWER/mem[6][3][13] ), .ip2(\ANSWER/mem[7][3][13] ), 
        .s(n11975), .op(n11891) );
  mux2_1 U13716 ( .ip1(n11892), .ip2(n11891), .s(n11950), .op(n11893) );
  mux2_1 U13717 ( .ip1(n11894), .ip2(n11893), .s(n11979), .op(n11896) );
  mux2_1 U13718 ( .ip1(\ANSWER/mem[8][3][13] ), .ip2(\ANSWER/mem[9][3][13] ), 
        .s(n11975), .op(n11895) );
  mux2_1 U13719 ( .ip1(n11896), .ip2(n11895), .s(n11983), .op(n11949) );
  mux2_1 U13720 ( .ip1(\ANSWER/mem[0][7][13] ), .ip2(\ANSWER/mem[1][7][13] ), 
        .s(n11982), .op(n11898) );
  mux2_1 U13721 ( .ip1(\ANSWER/mem[2][7][13] ), .ip2(\ANSWER/mem[3][7][13] ), 
        .s(n11982), .op(n11897) );
  mux2_1 U13722 ( .ip1(n11898), .ip2(n11897), .s(n11976), .op(n11902) );
  mux2_1 U13723 ( .ip1(\ANSWER/mem[4][7][13] ), .ip2(\ANSWER/mem[5][7][13] ), 
        .s(n11982), .op(n11900) );
  mux2_1 U13724 ( .ip1(\ANSWER/mem[6][7][13] ), .ip2(\ANSWER/mem[7][7][13] ), 
        .s(n11982), .op(n11899) );
  mux2_1 U13725 ( .ip1(n11900), .ip2(n11899), .s(n11976), .op(n11901) );
  mux2_1 U13726 ( .ip1(n11902), .ip2(n11901), .s(n11937), .op(n11904) );
  mux2_1 U13727 ( .ip1(\ANSWER/mem[8][7][13] ), .ip2(\ANSWER/mem[9][7][13] ), 
        .s(n11982), .op(n11903) );
  mux2_1 U13728 ( .ip1(n11904), .ip2(n11903), .s(n11983), .op(n11905) );
  and2_1 U13729 ( .ip1(n12186), .ip2(n11905), .op(n11948) );
  mux2_1 U13730 ( .ip1(\ANSWER/mem[0][4][13] ), .ip2(\ANSWER/mem[1][4][13] ), 
        .s(n11975), .op(n11907) );
  mux2_1 U13731 ( .ip1(\ANSWER/mem[2][4][13] ), .ip2(\ANSWER/mem[3][4][13] ), 
        .s(n11975), .op(n11906) );
  mux2_1 U13732 ( .ip1(n11907), .ip2(n11906), .s(n11950), .op(n11911) );
  mux2_1 U13733 ( .ip1(\ANSWER/mem[4][4][13] ), .ip2(\ANSWER/mem[5][4][13] ), 
        .s(n11975), .op(n11909) );
  mux2_1 U13734 ( .ip1(\ANSWER/mem[6][4][13] ), .ip2(\ANSWER/mem[7][4][13] ), 
        .s(n11975), .op(n11908) );
  mux2_1 U13735 ( .ip1(n11909), .ip2(n11908), .s(n11950), .op(n11910) );
  mux2_1 U13736 ( .ip1(n11911), .ip2(n11910), .s(n11937), .op(n11913) );
  mux2_1 U13737 ( .ip1(\ANSWER/mem[8][4][13] ), .ip2(\ANSWER/mem[9][4][13] ), 
        .s(n11975), .op(n11912) );
  mux2_1 U13738 ( .ip1(n11913), .ip2(n11912), .s(n11983), .op(n11914) );
  nand2_1 U13739 ( .ip1(n12176), .ip2(n11914), .op(n11946) );
  mux2_1 U13740 ( .ip1(\ANSWER/mem[0][5][13] ), .ip2(\ANSWER/mem[1][5][13] ), 
        .s(n11975), .op(n11916) );
  mux2_1 U13741 ( .ip1(\ANSWER/mem[2][5][13] ), .ip2(\ANSWER/mem[3][5][13] ), 
        .s(n11982), .op(n11915) );
  mux2_1 U13742 ( .ip1(n11916), .ip2(n11915), .s(n11950), .op(n11920) );
  mux2_1 U13743 ( .ip1(\ANSWER/mem[4][5][13] ), .ip2(\ANSWER/mem[5][5][13] ), 
        .s(n11982), .op(n11918) );
  mux2_1 U13744 ( .ip1(\ANSWER/mem[6][5][13] ), .ip2(\ANSWER/mem[7][5][13] ), 
        .s(n11982), .op(n11917) );
  mux2_1 U13745 ( .ip1(n11918), .ip2(n11917), .s(n11950), .op(n11919) );
  mux2_1 U13746 ( .ip1(n11920), .ip2(n11919), .s(n11937), .op(n11922) );
  mux2_1 U13747 ( .ip1(\ANSWER/mem[8][5][13] ), .ip2(\ANSWER/mem[9][5][13] ), 
        .s(n11982), .op(n11921) );
  mux2_1 U13748 ( .ip1(n11922), .ip2(n11921), .s(n11983), .op(n11923) );
  nand2_1 U13749 ( .ip1(n12127), .ip2(n11923), .op(n11945) );
  mux2_1 U13750 ( .ip1(\ANSWER/mem[0][0][13] ), .ip2(\ANSWER/mem[1][0][13] ), 
        .s(n8833), .op(n11925) );
  mux2_1 U13751 ( .ip1(\ANSWER/mem[2][0][13] ), .ip2(\ANSWER/mem[3][0][13] ), 
        .s(n11651), .op(n11924) );
  mux2_1 U13752 ( .ip1(n11925), .ip2(n11924), .s(n11950), .op(n11929) );
  mux2_1 U13753 ( .ip1(\ANSWER/mem[4][0][13] ), .ip2(\ANSWER/mem[5][0][13] ), 
        .s(n10583), .op(n11927) );
  mux2_1 U13754 ( .ip1(\ANSWER/mem[6][0][13] ), .ip2(\ANSWER/mem[7][0][13] ), 
        .s(n11758), .op(n11926) );
  mux2_1 U13755 ( .ip1(n11927), .ip2(n11926), .s(n11950), .op(n11928) );
  mux2_1 U13756 ( .ip1(n11929), .ip2(n11928), .s(n11937), .op(n11931) );
  mux2_1 U13757 ( .ip1(\ANSWER/mem[8][0][13] ), .ip2(\ANSWER/mem[9][0][13] ), 
        .s(n11113), .op(n11930) );
  mux2_1 U13758 ( .ip1(n11931), .ip2(n11930), .s(n11983), .op(n11932) );
  nand2_1 U13759 ( .ip1(n12108), .ip2(n11932), .op(n11944) );
  mux2_1 U13760 ( .ip1(\ANSWER/mem[0][2][13] ), .ip2(\ANSWER/mem[1][2][13] ), 
        .s(n8833), .op(n11934) );
  mux2_1 U13761 ( .ip1(\ANSWER/mem[2][2][13] ), .ip2(\ANSWER/mem[3][2][13] ), 
        .s(n8833), .op(n11933) );
  mux2_1 U13762 ( .ip1(n11934), .ip2(n11933), .s(n11950), .op(n11939) );
  mux2_1 U13763 ( .ip1(\ANSWER/mem[4][2][13] ), .ip2(\ANSWER/mem[5][2][13] ), 
        .s(n8833), .op(n11936) );
  mux2_1 U13764 ( .ip1(\ANSWER/mem[6][2][13] ), .ip2(\ANSWER/mem[7][2][13] ), 
        .s(n11975), .op(n11935) );
  mux2_1 U13765 ( .ip1(n11936), .ip2(n11935), .s(n11950), .op(n11938) );
  mux2_1 U13766 ( .ip1(n11939), .ip2(n11938), .s(n11937), .op(n11941) );
  mux2_1 U13767 ( .ip1(\ANSWER/mem[8][2][13] ), .ip2(\ANSWER/mem[9][2][13] ), 
        .s(n11975), .op(n11940) );
  mux2_1 U13768 ( .ip1(n11941), .ip2(n11940), .s(n11983), .op(n11942) );
  nand2_1 U13769 ( .ip1(n12147), .ip2(n11942), .op(n11943) );
  nand4_1 U13770 ( .ip1(n11946), .ip2(n11945), .ip3(n11944), .ip4(n11943), 
        .op(n11947) );
  not_ab_or_c_or_d U13771 ( .ip1(n11949), .ip2(n12137), .ip3(n11948), .ip4(
        n11947), .op(n11961) );
  mux2_1 U13772 ( .ip1(\ANSWER/mem[0][6][13] ), .ip2(\ANSWER/mem[1][6][13] ), 
        .s(n11982), .op(n11952) );
  mux2_1 U13773 ( .ip1(\ANSWER/mem[2][6][13] ), .ip2(\ANSWER/mem[3][6][13] ), 
        .s(n11982), .op(n11951) );
  mux2_1 U13774 ( .ip1(n11952), .ip2(n11951), .s(n11950), .op(n11956) );
  mux2_1 U13775 ( .ip1(\ANSWER/mem[4][6][13] ), .ip2(\ANSWER/mem[5][6][13] ), 
        .s(n11982), .op(n11954) );
  mux2_1 U13776 ( .ip1(\ANSWER/mem[6][6][13] ), .ip2(\ANSWER/mem[7][6][13] ), 
        .s(n11982), .op(n11953) );
  mux2_1 U13777 ( .ip1(n11954), .ip2(n11953), .s(n11976), .op(n11955) );
  mux2_1 U13778 ( .ip1(n11956), .ip2(n11955), .s(n11979), .op(n11958) );
  mux2_1 U13779 ( .ip1(\ANSWER/mem[8][6][13] ), .ip2(\ANSWER/mem[9][6][13] ), 
        .s(n11982), .op(n11957) );
  mux2_1 U13780 ( .ip1(n11958), .ip2(n11957), .s(n11983), .op(n11959) );
  nand2_1 U13781 ( .ip1(n12168), .ip2(n11959), .op(n11960) );
  nand3_1 U13782 ( .ip1(n11962), .ip2(n11961), .ip3(n11960), .op(n11963) );
  nand2_1 U13783 ( .ip1(n11963), .ip2(n12190), .op(n11989) );
  mux2_1 U13784 ( .ip1(\ANSWER/mem[0][9][13] ), .ip2(\ANSWER/mem[1][9][13] ), 
        .s(n11975), .op(n11965) );
  mux2_1 U13785 ( .ip1(\ANSWER/mem[2][9][13] ), .ip2(\ANSWER/mem[3][9][13] ), 
        .s(n11982), .op(n11964) );
  mux2_1 U13786 ( .ip1(n11965), .ip2(n11964), .s(n11976), .op(n11969) );
  mux2_1 U13787 ( .ip1(\ANSWER/mem[4][9][13] ), .ip2(\ANSWER/mem[5][9][13] ), 
        .s(n11975), .op(n11967) );
  mux2_1 U13788 ( .ip1(\ANSWER/mem[6][9][13] ), .ip2(\ANSWER/mem[7][9][13] ), 
        .s(n11982), .op(n11966) );
  mux2_1 U13789 ( .ip1(n11967), .ip2(n11966), .s(n11976), .op(n11968) );
  mux2_1 U13790 ( .ip1(n11969), .ip2(n11968), .s(n11979), .op(n11971) );
  mux2_1 U13791 ( .ip1(\ANSWER/mem[8][9][13] ), .ip2(\ANSWER/mem[9][9][13] ), 
        .s(n11982), .op(n11970) );
  mux2_1 U13792 ( .ip1(n11971), .ip2(n11970), .s(n11983), .op(n11972) );
  nand2_1 U13793 ( .ip1(n12215), .ip2(n11972), .op(n11988) );
  mux2_1 U13794 ( .ip1(\ANSWER/mem[0][8][13] ), .ip2(\ANSWER/mem[1][8][13] ), 
        .s(n11982), .op(n11974) );
  mux2_1 U13795 ( .ip1(\ANSWER/mem[2][8][13] ), .ip2(\ANSWER/mem[3][8][13] ), 
        .s(n11982), .op(n11973) );
  mux2_1 U13796 ( .ip1(n11974), .ip2(n11973), .s(n11976), .op(n11981) );
  mux2_1 U13797 ( .ip1(\ANSWER/mem[4][8][13] ), .ip2(\ANSWER/mem[5][8][13] ), 
        .s(n11975), .op(n11978) );
  mux2_1 U13798 ( .ip1(\ANSWER/mem[6][8][13] ), .ip2(\ANSWER/mem[7][8][13] ), 
        .s(n11982), .op(n11977) );
  mux2_1 U13799 ( .ip1(n11978), .ip2(n11977), .s(n11976), .op(n11980) );
  mux2_1 U13800 ( .ip1(n11981), .ip2(n11980), .s(n11979), .op(n11985) );
  mux2_1 U13801 ( .ip1(\ANSWER/mem[8][8][13] ), .ip2(\ANSWER/mem[9][8][13] ), 
        .s(n11982), .op(n11984) );
  mux2_1 U13802 ( .ip1(n11985), .ip2(n11984), .s(n11983), .op(n11986) );
  nand2_1 U13803 ( .ip1(n12201), .ip2(n11986), .op(n11987) );
  nand3_1 U13804 ( .ip1(n11989), .ip2(n11988), .ip3(n11987), .op(\ANSWER/N474 ) );
  mux2_1 U13805 ( .ip1(\ANSWER/mem[0][0][14] ), .ip2(\ANSWER/mem[1][0][14] ), 
        .s(n11164), .op(n11991) );
  mux2_1 U13806 ( .ip1(\ANSWER/mem[2][0][14] ), .ip2(\ANSWER/mem[3][0][14] ), 
        .s(n11546), .op(n11990) );
  inv_1 U13807 ( .ip(n12098), .op(n12062) );
  mux2_1 U13808 ( .ip1(n11991), .ip2(n11990), .s(n12062), .op(n11995) );
  mux2_1 U13809 ( .ip1(\ANSWER/mem[4][0][14] ), .ip2(\ANSWER/mem[5][0][14] ), 
        .s(n11223), .op(n11993) );
  mux2_1 U13810 ( .ip1(\ANSWER/mem[6][0][14] ), .ip2(\ANSWER/mem[7][0][14] ), 
        .s(n10816), .op(n11992) );
  mux2_1 U13811 ( .ip1(n11993), .ip2(n11992), .s(n12062), .op(n11994) );
  mux2_1 U13812 ( .ip1(n11995), .ip2(n11994), .s(n12088), .op(n11998) );
  mux2_1 U13813 ( .ip1(\ANSWER/mem[8][0][14] ), .ip2(\ANSWER/mem[9][0][14] ), 
        .s(n11506), .op(n11997) );
  inv_1 U13814 ( .ip(n11996), .op(n12211) );
  mux2_1 U13815 ( .ip1(n11998), .ip2(n11997), .s(n12211), .op(n11999) );
  nand2_1 U13816 ( .ip1(n12108), .ip2(n11999), .op(n12072) );
  mux2_1 U13817 ( .ip1(\ANSWER/mem[0][2][14] ), .ip2(\ANSWER/mem[1][2][14] ), 
        .s(n11164), .op(n12001) );
  mux2_1 U13818 ( .ip1(\ANSWER/mem[2][2][14] ), .ip2(\ANSWER/mem[3][2][14] ), 
        .s(n11164), .op(n12000) );
  mux2_1 U13819 ( .ip1(n12001), .ip2(n12000), .s(n12062), .op(n12005) );
  mux2_1 U13820 ( .ip1(\ANSWER/mem[4][2][14] ), .ip2(\ANSWER/mem[5][2][14] ), 
        .s(n11164), .op(n12003) );
  inv_1 U13821 ( .ip(n12109), .op(n12091) );
  mux2_1 U13822 ( .ip1(\ANSWER/mem[6][2][14] ), .ip2(\ANSWER/mem[7][2][14] ), 
        .s(n12091), .op(n12002) );
  mux2_1 U13823 ( .ip1(n12003), .ip2(n12002), .s(n12062), .op(n12004) );
  mux2_1 U13824 ( .ip1(n12005), .ip2(n12004), .s(n12088), .op(n12007) );
  mux2_1 U13825 ( .ip1(\ANSWER/mem[8][2][14] ), .ip2(\ANSWER/mem[9][2][14] ), 
        .s(n12091), .op(n12006) );
  mux2_1 U13826 ( .ip1(n12007), .ip2(n12006), .s(n12211), .op(n12059) );
  buf_1 U13827 ( .ip(n12091), .op(n12085) );
  mux2_1 U13828 ( .ip1(\ANSWER/mem[0][7][14] ), .ip2(\ANSWER/mem[1][7][14] ), 
        .s(n12085), .op(n12009) );
  mux2_1 U13829 ( .ip1(\ANSWER/mem[2][7][14] ), .ip2(\ANSWER/mem[3][7][14] ), 
        .s(n12085), .op(n12008) );
  mux2_1 U13830 ( .ip1(n12009), .ip2(n12008), .s(n11950), .op(n12013) );
  mux2_1 U13831 ( .ip1(\ANSWER/mem[4][7][14] ), .ip2(\ANSWER/mem[5][7][14] ), 
        .s(n12085), .op(n12011) );
  mux2_1 U13832 ( .ip1(\ANSWER/mem[6][7][14] ), .ip2(\ANSWER/mem[7][7][14] ), 
        .s(n12085), .op(n12010) );
  mux2_1 U13833 ( .ip1(n12011), .ip2(n12010), .s(n11842), .op(n12012) );
  mux2_1 U13834 ( .ip1(n12013), .ip2(n12012), .s(n12088), .op(n12015) );
  mux2_1 U13835 ( .ip1(\ANSWER/mem[8][7][14] ), .ip2(\ANSWER/mem[9][7][14] ), 
        .s(n12085), .op(n12014) );
  mux2_1 U13836 ( .ip1(n12015), .ip2(n12014), .s(n12211), .op(n12016) );
  and2_1 U13837 ( .ip1(n12186), .ip2(n12016), .op(n12058) );
  mux2_1 U13838 ( .ip1(\ANSWER/mem[0][4][14] ), .ip2(\ANSWER/mem[1][4][14] ), 
        .s(n12091), .op(n12018) );
  mux2_1 U13839 ( .ip1(\ANSWER/mem[2][4][14] ), .ip2(\ANSWER/mem[3][4][14] ), 
        .s(n12091), .op(n12017) );
  mux2_1 U13840 ( .ip1(n12018), .ip2(n12017), .s(n12062), .op(n12022) );
  mux2_1 U13841 ( .ip1(\ANSWER/mem[4][4][14] ), .ip2(\ANSWER/mem[5][4][14] ), 
        .s(n12091), .op(n12020) );
  mux2_1 U13842 ( .ip1(\ANSWER/mem[6][4][14] ), .ip2(\ANSWER/mem[7][4][14] ), 
        .s(n12091), .op(n12019) );
  mux2_1 U13843 ( .ip1(n12020), .ip2(n12019), .s(n12062), .op(n12021) );
  mux2_1 U13844 ( .ip1(n12022), .ip2(n12021), .s(n12088), .op(n12024) );
  mux2_1 U13845 ( .ip1(\ANSWER/mem[8][4][14] ), .ip2(\ANSWER/mem[9][4][14] ), 
        .s(n12091), .op(n12023) );
  mux2_1 U13846 ( .ip1(n12024), .ip2(n12023), .s(n12211), .op(n12025) );
  nand2_1 U13847 ( .ip1(n12176), .ip2(n12025), .op(n12056) );
  mux2_1 U13848 ( .ip1(\ANSWER/mem[0][5][14] ), .ip2(\ANSWER/mem[1][5][14] ), 
        .s(n12091), .op(n12027) );
  mux2_1 U13849 ( .ip1(\ANSWER/mem[2][5][14] ), .ip2(\ANSWER/mem[3][5][14] ), 
        .s(n12085), .op(n12026) );
  mux2_1 U13850 ( .ip1(n12027), .ip2(n12026), .s(n12062), .op(n12031) );
  mux2_1 U13851 ( .ip1(\ANSWER/mem[4][5][14] ), .ip2(\ANSWER/mem[5][5][14] ), 
        .s(n12085), .op(n12029) );
  mux2_1 U13852 ( .ip1(\ANSWER/mem[6][5][14] ), .ip2(\ANSWER/mem[7][5][14] ), 
        .s(n12085), .op(n12028) );
  mux2_1 U13853 ( .ip1(n12029), .ip2(n12028), .s(n12062), .op(n12030) );
  mux2_1 U13854 ( .ip1(n12031), .ip2(n12030), .s(n12088), .op(n12033) );
  mux2_1 U13855 ( .ip1(\ANSWER/mem[8][5][14] ), .ip2(\ANSWER/mem[9][5][14] ), 
        .s(n12085), .op(n12032) );
  mux2_1 U13856 ( .ip1(n12033), .ip2(n12032), .s(n12211), .op(n12034) );
  nand2_1 U13857 ( .ip1(n12127), .ip2(n12034), .op(n12055) );
  mux2_1 U13858 ( .ip1(\ANSWER/mem[0][1][14] ), .ip2(\ANSWER/mem[1][1][14] ), 
        .s(n12085), .op(n12036) );
  mux2_1 U13859 ( .ip1(\ANSWER/mem[2][1][14] ), .ip2(\ANSWER/mem[3][1][14] ), 
        .s(n11328), .op(n12035) );
  mux2_1 U13860 ( .ip1(n12036), .ip2(n12035), .s(n12062), .op(n12040) );
  mux2_1 U13861 ( .ip1(\ANSWER/mem[4][1][14] ), .ip2(\ANSWER/mem[5][1][14] ), 
        .s(n8833), .op(n12038) );
  mux2_1 U13862 ( .ip1(\ANSWER/mem[6][1][14] ), .ip2(\ANSWER/mem[7][1][14] ), 
        .s(n11506), .op(n12037) );
  mux2_1 U13863 ( .ip1(n12038), .ip2(n12037), .s(n12062), .op(n12039) );
  mux2_1 U13864 ( .ip1(n12040), .ip2(n12039), .s(n12088), .op(n12042) );
  mux2_1 U13865 ( .ip1(\ANSWER/mem[8][1][14] ), .ip2(\ANSWER/mem[9][1][14] ), 
        .s(n12085), .op(n12041) );
  mux2_1 U13866 ( .ip1(n12042), .ip2(n12041), .s(n12211), .op(n12043) );
  nand2_1 U13867 ( .ip1(n12157), .ip2(n12043), .op(n12054) );
  mux2_1 U13868 ( .ip1(\ANSWER/mem[0][6][14] ), .ip2(\ANSWER/mem[1][6][14] ), 
        .s(n12085), .op(n12045) );
  mux2_1 U13869 ( .ip1(\ANSWER/mem[2][6][14] ), .ip2(\ANSWER/mem[3][6][14] ), 
        .s(n12085), .op(n12044) );
  mux2_1 U13870 ( .ip1(n12045), .ip2(n12044), .s(n12062), .op(n12049) );
  mux2_1 U13871 ( .ip1(\ANSWER/mem[4][6][14] ), .ip2(\ANSWER/mem[5][6][14] ), 
        .s(n12085), .op(n12047) );
  mux2_1 U13872 ( .ip1(\ANSWER/mem[6][6][14] ), .ip2(\ANSWER/mem[7][6][14] ), 
        .s(n12085), .op(n12046) );
  mux2_1 U13873 ( .ip1(n12047), .ip2(n12046), .s(n11008), .op(n12048) );
  mux2_1 U13874 ( .ip1(n12049), .ip2(n12048), .s(n12088), .op(n12051) );
  mux2_1 U13875 ( .ip1(\ANSWER/mem[8][6][14] ), .ip2(\ANSWER/mem[9][6][14] ), 
        .s(n12085), .op(n12050) );
  mux2_1 U13876 ( .ip1(n12051), .ip2(n12050), .s(n12211), .op(n12052) );
  nand2_1 U13877 ( .ip1(n12168), .ip2(n12052), .op(n12053) );
  nand4_1 U13878 ( .ip1(n12056), .ip2(n12055), .ip3(n12054), .ip4(n12053), 
        .op(n12057) );
  not_ab_or_c_or_d U13879 ( .ip1(n12059), .ip2(n12147), .ip3(n12058), .ip4(
        n12057), .op(n12071) );
  mux2_1 U13880 ( .ip1(\ANSWER/mem[0][3][14] ), .ip2(\ANSWER/mem[1][3][14] ), 
        .s(n12091), .op(n12061) );
  mux2_1 U13881 ( .ip1(\ANSWER/mem[2][3][14] ), .ip2(\ANSWER/mem[3][3][14] ), 
        .s(n12091), .op(n12060) );
  mux2_1 U13882 ( .ip1(n12061), .ip2(n12060), .s(n12062), .op(n12066) );
  mux2_1 U13883 ( .ip1(\ANSWER/mem[4][3][14] ), .ip2(\ANSWER/mem[5][3][14] ), 
        .s(n12091), .op(n12064) );
  mux2_1 U13884 ( .ip1(\ANSWER/mem[6][3][14] ), .ip2(\ANSWER/mem[7][3][14] ), 
        .s(n12091), .op(n12063) );
  mux2_1 U13885 ( .ip1(n12064), .ip2(n12063), .s(n12062), .op(n12065) );
  mux2_1 U13886 ( .ip1(n12066), .ip2(n12065), .s(n12088), .op(n12068) );
  mux2_1 U13887 ( .ip1(\ANSWER/mem[8][3][14] ), .ip2(\ANSWER/mem[9][3][14] ), 
        .s(n12091), .op(n12067) );
  mux2_1 U13888 ( .ip1(n12068), .ip2(n12067), .s(n12211), .op(n12069) );
  nand2_1 U13889 ( .ip1(n12137), .ip2(n12069), .op(n12070) );
  nand3_1 U13890 ( .ip1(n12072), .ip2(n12071), .ip3(n12070), .op(n12073) );
  nand2_1 U13891 ( .ip1(n12073), .ip2(n12190), .op(n12097) );
  mux2_1 U13892 ( .ip1(\ANSWER/mem[0][8][14] ), .ip2(\ANSWER/mem[1][8][14] ), 
        .s(n12085), .op(n12075) );
  mux2_1 U13893 ( .ip1(\ANSWER/mem[2][8][14] ), .ip2(\ANSWER/mem[3][8][14] ), 
        .s(n12091), .op(n12074) );
  mux2_1 U13894 ( .ip1(n12075), .ip2(n12074), .s(n11868), .op(n12079) );
  mux2_1 U13895 ( .ip1(\ANSWER/mem[4][8][14] ), .ip2(\ANSWER/mem[5][8][14] ), 
        .s(n12091), .op(n12077) );
  mux2_1 U13896 ( .ip1(\ANSWER/mem[6][8][14] ), .ip2(\ANSWER/mem[7][8][14] ), 
        .s(n12091), .op(n12076) );
  mux2_1 U13897 ( .ip1(n12077), .ip2(n12076), .s(n12062), .op(n12078) );
  mux2_1 U13898 ( .ip1(n12079), .ip2(n12078), .s(n12088), .op(n12081) );
  mux2_1 U13899 ( .ip1(\ANSWER/mem[8][8][14] ), .ip2(\ANSWER/mem[9][8][14] ), 
        .s(n12091), .op(n12080) );
  mux2_1 U13900 ( .ip1(n12081), .ip2(n12080), .s(n12211), .op(n12082) );
  nand2_1 U13901 ( .ip1(n12201), .ip2(n12082), .op(n12096) );
  mux2_1 U13902 ( .ip1(\ANSWER/mem[0][9][14] ), .ip2(\ANSWER/mem[1][9][14] ), 
        .s(n12091), .op(n12084) );
  mux2_1 U13903 ( .ip1(\ANSWER/mem[2][9][14] ), .ip2(\ANSWER/mem[3][9][14] ), 
        .s(n12091), .op(n12083) );
  mux2_1 U13904 ( .ip1(n12084), .ip2(n12083), .s(n12158), .op(n12090) );
  mux2_1 U13905 ( .ip1(\ANSWER/mem[4][9][14] ), .ip2(\ANSWER/mem[5][9][14] ), 
        .s(n12085), .op(n12087) );
  mux2_1 U13906 ( .ip1(\ANSWER/mem[6][9][14] ), .ip2(\ANSWER/mem[7][9][14] ), 
        .s(n12091), .op(n12086) );
  mux2_1 U13907 ( .ip1(n12087), .ip2(n12086), .s(n11414), .op(n12089) );
  mux2_1 U13908 ( .ip1(n12090), .ip2(n12089), .s(n12088), .op(n12093) );
  mux2_1 U13909 ( .ip1(\ANSWER/mem[8][9][14] ), .ip2(\ANSWER/mem[9][9][14] ), 
        .s(n12091), .op(n12092) );
  mux2_1 U13910 ( .ip1(n12093), .ip2(n12092), .s(n12211), .op(n12094) );
  nand2_1 U13911 ( .ip1(n12215), .ip2(n12094), .op(n12095) );
  nand3_1 U13912 ( .ip1(n12097), .ip2(n12096), .ip3(n12095), .op(\ANSWER/N473 ) );
  mux2_1 U13913 ( .ip1(\ANSWER/mem[0][0][15] ), .ip2(\ANSWER/mem[1][0][15] ), 
        .s(n11437), .op(n12100) );
  mux2_1 U13914 ( .ip1(\ANSWER/mem[2][0][15] ), .ip2(\ANSWER/mem[3][0][15] ), 
        .s(n12085), .op(n12099) );
  inv_1 U13915 ( .ip(n12098), .op(n12158) );
  mux2_1 U13916 ( .ip1(n12100), .ip2(n12099), .s(n12158), .op(n12104) );
  mux2_1 U13917 ( .ip1(\ANSWER/mem[4][0][15] ), .ip2(\ANSWER/mem[5][0][15] ), 
        .s(n11873), .op(n12102) );
  mux2_1 U13918 ( .ip1(\ANSWER/mem[6][0][15] ), .ip2(\ANSWER/mem[7][0][15] ), 
        .s(n11113), .op(n12101) );
  mux2_1 U13919 ( .ip1(n12102), .ip2(n12101), .s(n12158), .op(n12103) );
  mux2_1 U13920 ( .ip1(n12104), .ip2(n12103), .s(n12207), .op(n12106) );
  mux2_1 U13921 ( .ip1(\ANSWER/mem[8][0][15] ), .ip2(\ANSWER/mem[9][0][15] ), 
        .s(n11223), .op(n12105) );
  mux2_1 U13922 ( .ip1(n12106), .ip2(n12105), .s(n12211), .op(n12107) );
  nand2_1 U13923 ( .ip1(n12108), .ip2(n12107), .op(n12189) );
  inv_1 U13924 ( .ip(n12109), .op(n12210) );
  mux2_1 U13925 ( .ip1(\ANSWER/mem[0][4][15] ), .ip2(\ANSWER/mem[1][4][15] ), 
        .s(n12210), .op(n12111) );
  mux2_1 U13926 ( .ip1(\ANSWER/mem[2][4][15] ), .ip2(\ANSWER/mem[3][4][15] ), 
        .s(n12210), .op(n12110) );
  mux2_1 U13927 ( .ip1(n12111), .ip2(n12110), .s(n12158), .op(n12115) );
  mux2_1 U13928 ( .ip1(\ANSWER/mem[4][4][15] ), .ip2(\ANSWER/mem[5][4][15] ), 
        .s(n12210), .op(n12113) );
  mux2_1 U13929 ( .ip1(\ANSWER/mem[6][4][15] ), .ip2(\ANSWER/mem[7][4][15] ), 
        .s(n12210), .op(n12112) );
  mux2_1 U13930 ( .ip1(n12113), .ip2(n12112), .s(n12158), .op(n12114) );
  mux2_1 U13931 ( .ip1(n12115), .ip2(n12114), .s(n12207), .op(n12117) );
  mux2_1 U13932 ( .ip1(\ANSWER/mem[8][4][15] ), .ip2(\ANSWER/mem[9][4][15] ), 
        .s(n12210), .op(n12116) );
  mux2_1 U13933 ( .ip1(n12117), .ip2(n12116), .s(n12211), .op(n12175) );
  mux2_1 U13934 ( .ip1(\ANSWER/mem[0][5][15] ), .ip2(\ANSWER/mem[1][5][15] ), 
        .s(n12210), .op(n12119) );
  buf_1 U13935 ( .ip(n12210), .op(n12204) );
  mux2_1 U13936 ( .ip1(\ANSWER/mem[2][5][15] ), .ip2(\ANSWER/mem[3][5][15] ), 
        .s(n12204), .op(n12118) );
  mux2_1 U13937 ( .ip1(n12119), .ip2(n12118), .s(n12158), .op(n12123) );
  mux2_1 U13938 ( .ip1(\ANSWER/mem[4][5][15] ), .ip2(\ANSWER/mem[5][5][15] ), 
        .s(n12204), .op(n12121) );
  mux2_1 U13939 ( .ip1(\ANSWER/mem[6][5][15] ), .ip2(\ANSWER/mem[7][5][15] ), 
        .s(n12204), .op(n12120) );
  mux2_1 U13940 ( .ip1(n12121), .ip2(n12120), .s(n12158), .op(n12122) );
  mux2_1 U13941 ( .ip1(n12123), .ip2(n12122), .s(n12207), .op(n12125) );
  mux2_1 U13942 ( .ip1(\ANSWER/mem[8][5][15] ), .ip2(\ANSWER/mem[9][5][15] ), 
        .s(n12204), .op(n12124) );
  mux2_1 U13943 ( .ip1(n12125), .ip2(n12124), .s(n12211), .op(n12126) );
  and2_1 U13944 ( .ip1(n12127), .ip2(n12126), .op(n12174) );
  mux2_1 U13945 ( .ip1(\ANSWER/mem[0][3][15] ), .ip2(\ANSWER/mem[1][3][15] ), 
        .s(n12210), .op(n12129) );
  mux2_1 U13946 ( .ip1(\ANSWER/mem[2][3][15] ), .ip2(\ANSWER/mem[3][3][15] ), 
        .s(n12210), .op(n12128) );
  mux2_1 U13947 ( .ip1(n12129), .ip2(n12128), .s(n12158), .op(n12133) );
  mux2_1 U13948 ( .ip1(\ANSWER/mem[4][3][15] ), .ip2(\ANSWER/mem[5][3][15] ), 
        .s(n12210), .op(n12131) );
  mux2_1 U13949 ( .ip1(\ANSWER/mem[6][3][15] ), .ip2(\ANSWER/mem[7][3][15] ), 
        .s(n12210), .op(n12130) );
  mux2_1 U13950 ( .ip1(n12131), .ip2(n12130), .s(n12158), .op(n12132) );
  mux2_1 U13951 ( .ip1(n12133), .ip2(n12132), .s(n12207), .op(n12135) );
  mux2_1 U13952 ( .ip1(\ANSWER/mem[8][3][15] ), .ip2(\ANSWER/mem[9][3][15] ), 
        .s(n12210), .op(n12134) );
  mux2_1 U13953 ( .ip1(n12135), .ip2(n12134), .s(n12211), .op(n12136) );
  nand2_1 U13954 ( .ip1(n12137), .ip2(n12136), .op(n12172) );
  mux2_1 U13955 ( .ip1(\ANSWER/mem[0][2][15] ), .ip2(\ANSWER/mem[1][2][15] ), 
        .s(n11113), .op(n12139) );
  mux2_1 U13956 ( .ip1(\ANSWER/mem[2][2][15] ), .ip2(\ANSWER/mem[3][2][15] ), 
        .s(n11873), .op(n12138) );
  mux2_1 U13957 ( .ip1(n12139), .ip2(n12138), .s(n12158), .op(n12143) );
  mux2_1 U13958 ( .ip1(\ANSWER/mem[4][2][15] ), .ip2(\ANSWER/mem[5][2][15] ), 
        .s(n11758), .op(n12141) );
  mux2_1 U13959 ( .ip1(\ANSWER/mem[6][2][15] ), .ip2(\ANSWER/mem[7][2][15] ), 
        .s(n12210), .op(n12140) );
  mux2_1 U13960 ( .ip1(n12141), .ip2(n12140), .s(n12158), .op(n12142) );
  mux2_1 U13961 ( .ip1(n12143), .ip2(n12142), .s(n12207), .op(n12145) );
  mux2_1 U13962 ( .ip1(\ANSWER/mem[8][2][15] ), .ip2(\ANSWER/mem[9][2][15] ), 
        .s(n12210), .op(n12144) );
  mux2_1 U13963 ( .ip1(n12145), .ip2(n12144), .s(n12211), .op(n12146) );
  nand2_1 U13964 ( .ip1(n12147), .ip2(n12146), .op(n12171) );
  mux2_1 U13965 ( .ip1(\ANSWER/mem[0][1][15] ), .ip2(\ANSWER/mem[1][1][15] ), 
        .s(n11223), .op(n12149) );
  mux2_1 U13966 ( .ip1(\ANSWER/mem[2][1][15] ), .ip2(\ANSWER/mem[3][1][15] ), 
        .s(n11546), .op(n12148) );
  mux2_1 U13967 ( .ip1(n12149), .ip2(n12148), .s(n12158), .op(n12153) );
  mux2_1 U13968 ( .ip1(\ANSWER/mem[4][1][15] ), .ip2(\ANSWER/mem[5][1][15] ), 
        .s(n12085), .op(n12151) );
  mux2_1 U13969 ( .ip1(\ANSWER/mem[6][1][15] ), .ip2(\ANSWER/mem[7][1][15] ), 
        .s(n10583), .op(n12150) );
  mux2_1 U13970 ( .ip1(n12151), .ip2(n12150), .s(n12158), .op(n12152) );
  mux2_1 U13971 ( .ip1(n12153), .ip2(n12152), .s(n12207), .op(n12155) );
  mux2_1 U13972 ( .ip1(\ANSWER/mem[8][1][15] ), .ip2(\ANSWER/mem[9][1][15] ), 
        .s(n11975), .op(n12154) );
  mux2_1 U13973 ( .ip1(n12155), .ip2(n12154), .s(n12211), .op(n12156) );
  nand2_1 U13974 ( .ip1(n12157), .ip2(n12156), .op(n12170) );
  mux2_1 U13975 ( .ip1(\ANSWER/mem[0][6][15] ), .ip2(\ANSWER/mem[1][6][15] ), 
        .s(n12204), .op(n12160) );
  mux2_1 U13976 ( .ip1(\ANSWER/mem[2][6][15] ), .ip2(\ANSWER/mem[3][6][15] ), 
        .s(n12204), .op(n12159) );
  mux2_1 U13977 ( .ip1(n12160), .ip2(n12159), .s(n12158), .op(n12164) );
  mux2_1 U13978 ( .ip1(\ANSWER/mem[4][6][15] ), .ip2(\ANSWER/mem[5][6][15] ), 
        .s(n12204), .op(n12162) );
  mux2_1 U13979 ( .ip1(\ANSWER/mem[6][6][15] ), .ip2(\ANSWER/mem[7][6][15] ), 
        .s(n12204), .op(n12161) );
  mux2_1 U13980 ( .ip1(n12162), .ip2(n12161), .s(n12062), .op(n12163) );
  mux2_1 U13981 ( .ip1(n12164), .ip2(n12163), .s(n12207), .op(n12166) );
  mux2_1 U13982 ( .ip1(\ANSWER/mem[8][6][15] ), .ip2(\ANSWER/mem[9][6][15] ), 
        .s(n12204), .op(n12165) );
  mux2_1 U13983 ( .ip1(n12166), .ip2(n12165), .s(n12211), .op(n12167) );
  nand2_1 U13984 ( .ip1(n12168), .ip2(n12167), .op(n12169) );
  nand4_1 U13985 ( .ip1(n12172), .ip2(n12171), .ip3(n12170), .ip4(n12169), 
        .op(n12173) );
  not_ab_or_c_or_d U13986 ( .ip1(n12176), .ip2(n12175), .ip3(n12174), .ip4(
        n12173), .op(n12188) );
  mux2_1 U13987 ( .ip1(\ANSWER/mem[0][7][15] ), .ip2(\ANSWER/mem[1][7][15] ), 
        .s(n12204), .op(n12178) );
  mux2_1 U13988 ( .ip1(\ANSWER/mem[2][7][15] ), .ip2(\ANSWER/mem[3][7][15] ), 
        .s(n12204), .op(n12177) );
  mux2_1 U13989 ( .ip1(n12178), .ip2(n12177), .s(n11507), .op(n12182) );
  mux2_1 U13990 ( .ip1(\ANSWER/mem[4][7][15] ), .ip2(\ANSWER/mem[5][7][15] ), 
        .s(n12204), .op(n12180) );
  mux2_1 U13991 ( .ip1(\ANSWER/mem[6][7][15] ), .ip2(\ANSWER/mem[7][7][15] ), 
        .s(n12204), .op(n12179) );
  mux2_1 U13992 ( .ip1(n12180), .ip2(n12179), .s(n11183), .op(n12181) );
  mux2_1 U13993 ( .ip1(n12182), .ip2(n12181), .s(n12207), .op(n12184) );
  mux2_1 U13994 ( .ip1(\ANSWER/mem[8][7][15] ), .ip2(\ANSWER/mem[9][7][15] ), 
        .s(n12210), .op(n12183) );
  mux2_1 U13995 ( .ip1(n12184), .ip2(n12183), .s(n12211), .op(n12185) );
  nand2_1 U13996 ( .ip1(n12186), .ip2(n12185), .op(n12187) );
  nand3_1 U13997 ( .ip1(n12189), .ip2(n12188), .ip3(n12187), .op(n12191) );
  nand2_1 U13998 ( .ip1(n12191), .ip2(n12190), .op(n12218) );
  mux2_1 U13999 ( .ip1(\ANSWER/mem[0][8][15] ), .ip2(\ANSWER/mem[1][8][15] ), 
        .s(n12204), .op(n12193) );
  mux2_1 U14000 ( .ip1(\ANSWER/mem[2][8][15] ), .ip2(\ANSWER/mem[3][8][15] ), 
        .s(n12210), .op(n12192) );
  mux2_1 U14001 ( .ip1(n12193), .ip2(n12192), .s(n11950), .op(n12197) );
  mux2_1 U14002 ( .ip1(\ANSWER/mem[4][8][15] ), .ip2(\ANSWER/mem[5][8][15] ), 
        .s(n12204), .op(n12195) );
  mux2_1 U14003 ( .ip1(\ANSWER/mem[6][8][15] ), .ip2(\ANSWER/mem[7][8][15] ), 
        .s(n12210), .op(n12194) );
  mux2_1 U14004 ( .ip1(n12195), .ip2(n12194), .s(n11224), .op(n12196) );
  mux2_1 U14005 ( .ip1(n12197), .ip2(n12196), .s(n12207), .op(n12199) );
  mux2_1 U14006 ( .ip1(\ANSWER/mem[8][8][15] ), .ip2(\ANSWER/mem[9][8][15] ), 
        .s(n12210), .op(n12198) );
  mux2_1 U14007 ( .ip1(n12199), .ip2(n12198), .s(n12211), .op(n12200) );
  nand2_1 U14008 ( .ip1(n12201), .ip2(n12200), .op(n12217) );
  mux2_1 U14009 ( .ip1(\ANSWER/mem[0][9][15] ), .ip2(\ANSWER/mem[1][9][15] ), 
        .s(n12210), .op(n12203) );
  mux2_1 U14010 ( .ip1(\ANSWER/mem[2][9][15] ), .ip2(\ANSWER/mem[3][9][15] ), 
        .s(n12210), .op(n12202) );
  mux2_1 U14011 ( .ip1(n12203), .ip2(n12202), .s(n11008), .op(n12209) );
  mux2_1 U14012 ( .ip1(\ANSWER/mem[4][9][15] ), .ip2(\ANSWER/mem[5][9][15] ), 
        .s(n12204), .op(n12206) );
  mux2_1 U14013 ( .ip1(\ANSWER/mem[6][9][15] ), .ip2(\ANSWER/mem[7][9][15] ), 
        .s(n12210), .op(n12205) );
  mux2_1 U14014 ( .ip1(n12206), .ip2(n12205), .s(n11008), .op(n12208) );
  mux2_1 U14015 ( .ip1(n12209), .ip2(n12208), .s(n12207), .op(n12213) );
  mux2_1 U14016 ( .ip1(\ANSWER/mem[8][9][15] ), .ip2(\ANSWER/mem[9][9][15] ), 
        .s(n12210), .op(n12212) );
  mux2_1 U14017 ( .ip1(n12213), .ip2(n12212), .s(n12211), .op(n12214) );
  nand2_1 U14018 ( .ip1(n12215), .ip2(n12214), .op(n12216) );
  nand3_1 U14019 ( .ip1(n12218), .ip2(n12217), .ip3(n12216), .op(\ANSWER/N472 ) );
endmodule

