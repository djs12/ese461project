
module Top ( clk, reset, inputSramWe, pixels, weight1, w2SramWeOffChip, 
        weight2, weight2AddrOffChip, weight2_loadNextRow, rdata );
  input [159:0] pixels;
  input [15:0] weight1;
  input [15:0] weight2;
  input [3:0] weight2AddrOffChip;
  output [15:0] rdata;
  input clk, reset, inputSramWe, w2SramWeOffChip;
  output weight2_loadNextRow;
  wire   \INPUTSRAM/mem_i[9][15] , \INPUTSRAM/mem_i[9][14] ,
         \INPUTSRAM/mem_i[9][13] , \INPUTSRAM/mem_i[9][12] ,
         \INPUTSRAM/mem_i[9][11] , \INPUTSRAM/mem_i[9][10] ,
         \INPUTSRAM/mem_i[9][9] , \INPUTSRAM/mem_i[9][8] ,
         \INPUTSRAM/mem_i[9][7] , \INPUTSRAM/mem_i[9][6] ,
         \INPUTSRAM/mem_i[9][5] , \INPUTSRAM/mem_i[9][4] ,
         \INPUTSRAM/mem_i[9][3] , \INPUTSRAM/mem_i[9][2] ,
         \INPUTSRAM/mem_i[9][1] , \INPUTSRAM/mem_i[9][0] ,
         \INPUTSRAM/mem_i[8][15] , \INPUTSRAM/mem_i[8][14] ,
         \INPUTSRAM/mem_i[8][13] , \INPUTSRAM/mem_i[8][12] ,
         \INPUTSRAM/mem_i[8][11] , \INPUTSRAM/mem_i[8][10] ,
         \INPUTSRAM/mem_i[8][9] , \INPUTSRAM/mem_i[8][8] ,
         \INPUTSRAM/mem_i[8][7] , \INPUTSRAM/mem_i[8][6] ,
         \INPUTSRAM/mem_i[8][5] , \INPUTSRAM/mem_i[8][4] ,
         \INPUTSRAM/mem_i[8][3] , \INPUTSRAM/mem_i[8][2] ,
         \INPUTSRAM/mem_i[8][1] , \INPUTSRAM/mem_i[8][0] ,
         \INPUTSRAM/mem_i[7][15] , \INPUTSRAM/mem_i[7][14] ,
         \INPUTSRAM/mem_i[7][13] , \INPUTSRAM/mem_i[7][12] ,
         \INPUTSRAM/mem_i[7][11] , \INPUTSRAM/mem_i[7][10] ,
         \INPUTSRAM/mem_i[7][9] , \INPUTSRAM/mem_i[7][8] ,
         \INPUTSRAM/mem_i[7][7] , \INPUTSRAM/mem_i[7][6] ,
         \INPUTSRAM/mem_i[7][5] , \INPUTSRAM/mem_i[7][4] ,
         \INPUTSRAM/mem_i[7][3] , \INPUTSRAM/mem_i[7][2] ,
         \INPUTSRAM/mem_i[7][1] , \INPUTSRAM/mem_i[7][0] ,
         \INPUTSRAM/mem_i[6][15] , \INPUTSRAM/mem_i[6][14] ,
         \INPUTSRAM/mem_i[6][13] , \INPUTSRAM/mem_i[6][12] ,
         \INPUTSRAM/mem_i[6][11] , \INPUTSRAM/mem_i[6][10] ,
         \INPUTSRAM/mem_i[6][9] , \INPUTSRAM/mem_i[6][8] ,
         \INPUTSRAM/mem_i[6][7] , \INPUTSRAM/mem_i[6][6] ,
         \INPUTSRAM/mem_i[6][5] , \INPUTSRAM/mem_i[6][4] ,
         \INPUTSRAM/mem_i[6][3] , \INPUTSRAM/mem_i[6][2] ,
         \INPUTSRAM/mem_i[6][1] , \INPUTSRAM/mem_i[6][0] ,
         \INPUTSRAM/mem_i[5][15] , \INPUTSRAM/mem_i[5][14] ,
         \INPUTSRAM/mem_i[5][13] , \INPUTSRAM/mem_i[5][12] ,
         \INPUTSRAM/mem_i[5][11] , \INPUTSRAM/mem_i[5][10] ,
         \INPUTSRAM/mem_i[5][9] , \INPUTSRAM/mem_i[5][8] ,
         \INPUTSRAM/mem_i[5][7] , \INPUTSRAM/mem_i[5][6] ,
         \INPUTSRAM/mem_i[5][5] , \INPUTSRAM/mem_i[5][4] ,
         \INPUTSRAM/mem_i[5][3] , \INPUTSRAM/mem_i[5][2] ,
         \INPUTSRAM/mem_i[5][1] , \INPUTSRAM/mem_i[5][0] ,
         \INPUTSRAM/mem_i[4][15] , \INPUTSRAM/mem_i[4][14] ,
         \INPUTSRAM/mem_i[4][13] , \INPUTSRAM/mem_i[4][12] ,
         \INPUTSRAM/mem_i[4][11] , \INPUTSRAM/mem_i[4][10] ,
         \INPUTSRAM/mem_i[4][9] , \INPUTSRAM/mem_i[4][8] ,
         \INPUTSRAM/mem_i[4][7] , \INPUTSRAM/mem_i[4][6] ,
         \INPUTSRAM/mem_i[4][5] , \INPUTSRAM/mem_i[4][4] ,
         \INPUTSRAM/mem_i[4][3] , \INPUTSRAM/mem_i[4][2] ,
         \INPUTSRAM/mem_i[4][1] , \INPUTSRAM/mem_i[4][0] ,
         \INPUTSRAM/mem_i[3][15] , \INPUTSRAM/mem_i[3][14] ,
         \INPUTSRAM/mem_i[3][13] , \INPUTSRAM/mem_i[3][12] ,
         \INPUTSRAM/mem_i[3][11] , \INPUTSRAM/mem_i[3][10] ,
         \INPUTSRAM/mem_i[3][9] , \INPUTSRAM/mem_i[3][8] ,
         \INPUTSRAM/mem_i[3][7] , \INPUTSRAM/mem_i[3][6] ,
         \INPUTSRAM/mem_i[3][5] , \INPUTSRAM/mem_i[3][4] ,
         \INPUTSRAM/mem_i[3][3] , \INPUTSRAM/mem_i[3][2] ,
         \INPUTSRAM/mem_i[3][1] , \INPUTSRAM/mem_i[3][0] ,
         \INPUTSRAM/mem_i[2][14] , \INPUTSRAM/mem_i[2][13] ,
         \INPUTSRAM/mem_i[2][12] , \INPUTSRAM/mem_i[2][11] ,
         \INPUTSRAM/mem_i[2][10] , \INPUTSRAM/mem_i[2][9] ,
         \INPUTSRAM/mem_i[2][8] , \INPUTSRAM/mem_i[2][7] ,
         \INPUTSRAM/mem_i[2][6] , \INPUTSRAM/mem_i[2][5] ,
         \INPUTSRAM/mem_i[2][4] , \INPUTSRAM/mem_i[2][3] ,
         \INPUTSRAM/mem_i[2][2] , \INPUTSRAM/mem_i[2][1] ,
         \INPUTSRAM/mem_i[2][0] , \INPUTSRAM/mem_i[1][15] ,
         \INPUTSRAM/mem_i[1][14] , \INPUTSRAM/mem_i[1][13] ,
         \INPUTSRAM/mem_i[1][12] , \INPUTSRAM/mem_i[1][11] ,
         \INPUTSRAM/mem_i[1][10] , \INPUTSRAM/mem_i[1][9] ,
         \INPUTSRAM/mem_i[1][8] , \INPUTSRAM/mem_i[1][7] ,
         \INPUTSRAM/mem_i[1][6] , \INPUTSRAM/mem_i[1][5] ,
         \INPUTSRAM/mem_i[1][4] , \INPUTSRAM/mem_i[1][3] ,
         \INPUTSRAM/mem_i[1][2] , \INPUTSRAM/mem_i[1][1] ,
         \INPUTSRAM/mem_i[1][0] , \INPUTSRAM/mem_i[0][14] ,
         \INPUTSRAM/mem_i[0][13] , \INPUTSRAM/mem_i[0][12] ,
         \INPUTSRAM/mem_i[0][11] , \INPUTSRAM/mem_i[0][10] ,
         \INPUTSRAM/mem_i[0][9] , \INPUTSRAM/mem_i[0][8] ,
         \INPUTSRAM/mem_i[0][7] , \INPUTSRAM/mem_i[0][6] ,
         \INPUTSRAM/mem_i[0][5] , \INPUTSRAM/mem_i[0][4] ,
         \INPUTSRAM/mem_i[0][3] , \INPUTSRAM/mem_i[0][2] ,
         \INPUTSRAM/mem_i[0][1] , \INPUTSRAM/mem_i[0][0] , \CNTRL/N242 ,
         \CNTRL/N241 , \CNTRL/N240 , \CNTRL/N239 , \CNTRL/N238 , \CNTRL/N237 ,
         \CNTRL/N236 , \CNTRL/N235 , \CNTRL/N234 , \CNTRL/N233 ,
         \WEIGHT_2/mem_w2[9][15] , \WEIGHT_2/mem_w2[9][14] ,
         \WEIGHT_2/mem_w2[9][13] , \WEIGHT_2/mem_w2[9][12] ,
         \WEIGHT_2/mem_w2[9][11] , \WEIGHT_2/mem_w2[9][10] ,
         \WEIGHT_2/mem_w2[9][9] , \WEIGHT_2/mem_w2[9][8] ,
         \WEIGHT_2/mem_w2[9][7] , \WEIGHT_2/mem_w2[9][6] ,
         \WEIGHT_2/mem_w2[9][5] , \WEIGHT_2/mem_w2[9][4] ,
         \WEIGHT_2/mem_w2[9][3] , \WEIGHT_2/mem_w2[9][2] ,
         \WEIGHT_2/mem_w2[9][1] , \WEIGHT_2/mem_w2[9][0] ,
         \WEIGHT_2/mem_w2[8][15] , \WEIGHT_2/mem_w2[8][14] ,
         \WEIGHT_2/mem_w2[8][13] , \WEIGHT_2/mem_w2[8][12] ,
         \WEIGHT_2/mem_w2[8][11] , \WEIGHT_2/mem_w2[8][10] ,
         \WEIGHT_2/mem_w2[8][9] , \WEIGHT_2/mem_w2[8][8] ,
         \WEIGHT_2/mem_w2[8][7] , \WEIGHT_2/mem_w2[8][6] ,
         \WEIGHT_2/mem_w2[8][5] , \WEIGHT_2/mem_w2[8][4] ,
         \WEIGHT_2/mem_w2[8][3] , \WEIGHT_2/mem_w2[8][2] ,
         \WEIGHT_2/mem_w2[8][1] , \WEIGHT_2/mem_w2[8][0] ,
         \WEIGHT_2/mem_w2[7][15] , \WEIGHT_2/mem_w2[7][14] ,
         \WEIGHT_2/mem_w2[7][13] , \WEIGHT_2/mem_w2[7][12] ,
         \WEIGHT_2/mem_w2[7][11] , \WEIGHT_2/mem_w2[7][10] ,
         \WEIGHT_2/mem_w2[7][9] , \WEIGHT_2/mem_w2[7][8] ,
         \WEIGHT_2/mem_w2[7][7] , \WEIGHT_2/mem_w2[7][6] ,
         \WEIGHT_2/mem_w2[7][5] , \WEIGHT_2/mem_w2[7][4] ,
         \WEIGHT_2/mem_w2[7][3] , \WEIGHT_2/mem_w2[7][2] ,
         \WEIGHT_2/mem_w2[7][1] , \WEIGHT_2/mem_w2[7][0] ,
         \WEIGHT_2/mem_w2[6][15] , \WEIGHT_2/mem_w2[6][14] ,
         \WEIGHT_2/mem_w2[6][13] , \WEIGHT_2/mem_w2[6][12] ,
         \WEIGHT_2/mem_w2[6][11] , \WEIGHT_2/mem_w2[6][10] ,
         \WEIGHT_2/mem_w2[6][9] , \WEIGHT_2/mem_w2[6][8] ,
         \WEIGHT_2/mem_w2[6][7] , \WEIGHT_2/mem_w2[6][6] ,
         \WEIGHT_2/mem_w2[6][5] , \WEIGHT_2/mem_w2[6][4] ,
         \WEIGHT_2/mem_w2[6][3] , \WEIGHT_2/mem_w2[6][2] ,
         \WEIGHT_2/mem_w2[6][1] , \WEIGHT_2/mem_w2[6][0] ,
         \WEIGHT_2/mem_w2[5][15] , \WEIGHT_2/mem_w2[5][14] ,
         \WEIGHT_2/mem_w2[5][13] , \WEIGHT_2/mem_w2[5][12] ,
         \WEIGHT_2/mem_w2[5][11] , \WEIGHT_2/mem_w2[5][10] ,
         \WEIGHT_2/mem_w2[5][9] , \WEIGHT_2/mem_w2[5][8] ,
         \WEIGHT_2/mem_w2[5][7] , \WEIGHT_2/mem_w2[5][6] ,
         \WEIGHT_2/mem_w2[5][5] , \WEIGHT_2/mem_w2[5][4] ,
         \WEIGHT_2/mem_w2[5][3] , \WEIGHT_2/mem_w2[5][2] ,
         \WEIGHT_2/mem_w2[5][1] , \WEIGHT_2/mem_w2[5][0] ,
         \WEIGHT_2/mem_w2[4][15] , \WEIGHT_2/mem_w2[4][14] ,
         \WEIGHT_2/mem_w2[4][13] , \WEIGHT_2/mem_w2[4][12] ,
         \WEIGHT_2/mem_w2[4][11] , \WEIGHT_2/mem_w2[4][10] ,
         \WEIGHT_2/mem_w2[4][9] , \WEIGHT_2/mem_w2[4][8] ,
         \WEIGHT_2/mem_w2[4][7] , \WEIGHT_2/mem_w2[4][6] ,
         \WEIGHT_2/mem_w2[4][5] , \WEIGHT_2/mem_w2[4][4] ,
         \WEIGHT_2/mem_w2[4][3] , \WEIGHT_2/mem_w2[4][2] ,
         \WEIGHT_2/mem_w2[4][1] , \WEIGHT_2/mem_w2[4][0] ,
         \WEIGHT_2/mem_w2[3][15] , \WEIGHT_2/mem_w2[3][14] ,
         \WEIGHT_2/mem_w2[3][13] , \WEIGHT_2/mem_w2[3][12] ,
         \WEIGHT_2/mem_w2[3][11] , \WEIGHT_2/mem_w2[3][10] ,
         \WEIGHT_2/mem_w2[3][9] , \WEIGHT_2/mem_w2[3][8] ,
         \WEIGHT_2/mem_w2[3][7] , \WEIGHT_2/mem_w2[3][6] ,
         \WEIGHT_2/mem_w2[3][5] , \WEIGHT_2/mem_w2[3][4] ,
         \WEIGHT_2/mem_w2[3][3] , \WEIGHT_2/mem_w2[3][2] ,
         \WEIGHT_2/mem_w2[3][1] , \WEIGHT_2/mem_w2[3][0] ,
         \WEIGHT_2/mem_w2[2][15] , \WEIGHT_2/mem_w2[2][14] ,
         \WEIGHT_2/mem_w2[2][13] , \WEIGHT_2/mem_w2[2][12] ,
         \WEIGHT_2/mem_w2[2][11] , \WEIGHT_2/mem_w2[2][10] ,
         \WEIGHT_2/mem_w2[2][9] , \WEIGHT_2/mem_w2[2][8] ,
         \WEIGHT_2/mem_w2[2][7] , \WEIGHT_2/mem_w2[2][6] ,
         \WEIGHT_2/mem_w2[2][5] , \WEIGHT_2/mem_w2[2][4] ,
         \WEIGHT_2/mem_w2[2][3] , \WEIGHT_2/mem_w2[2][2] ,
         \WEIGHT_2/mem_w2[2][1] , \WEIGHT_2/mem_w2[2][0] ,
         \WEIGHT_2/mem_w2[1][15] , \WEIGHT_2/mem_w2[1][14] ,
         \WEIGHT_2/mem_w2[1][13] , \WEIGHT_2/mem_w2[1][12] ,
         \WEIGHT_2/mem_w2[1][11] , \WEIGHT_2/mem_w2[1][10] ,
         \WEIGHT_2/mem_w2[1][9] , \WEIGHT_2/mem_w2[1][8] ,
         \WEIGHT_2/mem_w2[1][7] , \WEIGHT_2/mem_w2[1][6] ,
         \WEIGHT_2/mem_w2[1][5] , \WEIGHT_2/mem_w2[1][4] ,
         \WEIGHT_2/mem_w2[1][3] , \WEIGHT_2/mem_w2[1][2] ,
         \WEIGHT_2/mem_w2[1][1] , \WEIGHT_2/mem_w2[1][0] ,
         \WEIGHT_2/mem_w2[0][15] , \WEIGHT_2/mem_w2[0][14] ,
         \WEIGHT_2/mem_w2[0][13] , \WEIGHT_2/mem_w2[0][12] ,
         \WEIGHT_2/mem_w2[0][11] , \WEIGHT_2/mem_w2[0][10] ,
         \WEIGHT_2/mem_w2[0][9] , \WEIGHT_2/mem_w2[0][8] ,
         \WEIGHT_2/mem_w2[0][7] , \WEIGHT_2/mem_w2[0][6] ,
         \WEIGHT_2/mem_w2[0][5] , \WEIGHT_2/mem_w2[0][4] ,
         \WEIGHT_2/mem_w2[0][3] , \WEIGHT_2/mem_w2[0][2] ,
         \WEIGHT_2/mem_w2[0][1] , \WEIGHT_2/mem_w2[0][0] , \ANSWER/N487 ,
         \ANSWER/N486 , \ANSWER/N485 , \ANSWER/N484 , \ANSWER/N483 ,
         \ANSWER/N482 , \ANSWER/N481 , \ANSWER/N480 , \ANSWER/N479 ,
         \ANSWER/N478 , \ANSWER/N477 , \ANSWER/N476 , \ANSWER/N475 ,
         \ANSWER/N474 , \ANSWER/N473 , \ANSWER/N472 , \ANSWER/mem[9][9][15] ,
         \ANSWER/mem[9][9][14] , \ANSWER/mem[9][9][13] ,
         \ANSWER/mem[9][9][12] , \ANSWER/mem[9][9][11] ,
         \ANSWER/mem[9][9][10] , \ANSWER/mem[9][9][9] , \ANSWER/mem[9][9][8] ,
         \ANSWER/mem[9][9][7] , \ANSWER/mem[9][9][6] , \ANSWER/mem[9][9][5] ,
         \ANSWER/mem[9][9][4] , \ANSWER/mem[9][9][3] , \ANSWER/mem[9][9][2] ,
         \ANSWER/mem[9][9][1] , \ANSWER/mem[9][9][0] , \ANSWER/mem[9][8][15] ,
         \ANSWER/mem[9][8][14] , \ANSWER/mem[9][8][13] ,
         \ANSWER/mem[9][8][12] , \ANSWER/mem[9][8][11] ,
         \ANSWER/mem[9][8][10] , \ANSWER/mem[9][8][9] , \ANSWER/mem[9][8][8] ,
         \ANSWER/mem[9][8][7] , \ANSWER/mem[9][8][6] , \ANSWER/mem[9][8][5] ,
         \ANSWER/mem[9][8][4] , \ANSWER/mem[9][8][3] , \ANSWER/mem[9][8][2] ,
         \ANSWER/mem[9][8][1] , \ANSWER/mem[9][8][0] , \ANSWER/mem[9][7][15] ,
         \ANSWER/mem[9][7][14] , \ANSWER/mem[9][7][13] ,
         \ANSWER/mem[9][7][12] , \ANSWER/mem[9][7][11] ,
         \ANSWER/mem[9][7][10] , \ANSWER/mem[9][7][9] , \ANSWER/mem[9][7][8] ,
         \ANSWER/mem[9][7][7] , \ANSWER/mem[9][7][6] , \ANSWER/mem[9][7][5] ,
         \ANSWER/mem[9][7][4] , \ANSWER/mem[9][7][3] , \ANSWER/mem[9][7][2] ,
         \ANSWER/mem[9][7][1] , \ANSWER/mem[9][7][0] , \ANSWER/mem[9][6][15] ,
         \ANSWER/mem[9][6][14] , \ANSWER/mem[9][6][13] ,
         \ANSWER/mem[9][6][12] , \ANSWER/mem[9][6][11] ,
         \ANSWER/mem[9][6][10] , \ANSWER/mem[9][6][9] , \ANSWER/mem[9][6][8] ,
         \ANSWER/mem[9][6][7] , \ANSWER/mem[9][6][6] , \ANSWER/mem[9][6][5] ,
         \ANSWER/mem[9][6][4] , \ANSWER/mem[9][6][3] , \ANSWER/mem[9][6][2] ,
         \ANSWER/mem[9][6][1] , \ANSWER/mem[9][6][0] , \ANSWER/mem[9][5][15] ,
         \ANSWER/mem[9][5][14] , \ANSWER/mem[9][5][13] ,
         \ANSWER/mem[9][5][12] , \ANSWER/mem[9][5][11] ,
         \ANSWER/mem[9][5][10] , \ANSWER/mem[9][5][9] , \ANSWER/mem[9][5][8] ,
         \ANSWER/mem[9][5][7] , \ANSWER/mem[9][5][6] , \ANSWER/mem[9][5][5] ,
         \ANSWER/mem[9][5][4] , \ANSWER/mem[9][5][3] , \ANSWER/mem[9][5][2] ,
         \ANSWER/mem[9][5][1] , \ANSWER/mem[9][5][0] , \ANSWER/mem[9][4][15] ,
         \ANSWER/mem[9][4][14] , \ANSWER/mem[9][4][13] ,
         \ANSWER/mem[9][4][12] , \ANSWER/mem[9][4][11] ,
         \ANSWER/mem[9][4][10] , \ANSWER/mem[9][4][9] , \ANSWER/mem[9][4][8] ,
         \ANSWER/mem[9][4][7] , \ANSWER/mem[9][4][6] , \ANSWER/mem[9][4][5] ,
         \ANSWER/mem[9][4][4] , \ANSWER/mem[9][4][3] , \ANSWER/mem[9][4][2] ,
         \ANSWER/mem[9][4][1] , \ANSWER/mem[9][4][0] , \ANSWER/mem[9][3][15] ,
         \ANSWER/mem[9][3][14] , \ANSWER/mem[9][3][13] ,
         \ANSWER/mem[9][3][12] , \ANSWER/mem[9][3][11] ,
         \ANSWER/mem[9][3][10] , \ANSWER/mem[9][3][9] , \ANSWER/mem[9][3][8] ,
         \ANSWER/mem[9][3][7] , \ANSWER/mem[9][3][6] , \ANSWER/mem[9][3][5] ,
         \ANSWER/mem[9][3][4] , \ANSWER/mem[9][3][3] , \ANSWER/mem[9][3][2] ,
         \ANSWER/mem[9][3][1] , \ANSWER/mem[9][3][0] , \ANSWER/mem[9][2][15] ,
         \ANSWER/mem[9][2][14] , \ANSWER/mem[9][2][13] ,
         \ANSWER/mem[9][2][12] , \ANSWER/mem[9][2][11] ,
         \ANSWER/mem[9][2][10] , \ANSWER/mem[9][2][9] , \ANSWER/mem[9][2][8] ,
         \ANSWER/mem[9][2][7] , \ANSWER/mem[9][2][6] , \ANSWER/mem[9][2][5] ,
         \ANSWER/mem[9][2][4] , \ANSWER/mem[9][2][3] , \ANSWER/mem[9][2][2] ,
         \ANSWER/mem[9][2][1] , \ANSWER/mem[9][2][0] , \ANSWER/mem[9][1][15] ,
         \ANSWER/mem[9][1][14] , \ANSWER/mem[9][1][13] ,
         \ANSWER/mem[9][1][12] , \ANSWER/mem[9][1][11] ,
         \ANSWER/mem[9][1][10] , \ANSWER/mem[9][1][9] , \ANSWER/mem[9][1][8] ,
         \ANSWER/mem[9][1][7] , \ANSWER/mem[9][1][6] , \ANSWER/mem[9][1][5] ,
         \ANSWER/mem[9][1][4] , \ANSWER/mem[9][1][3] , \ANSWER/mem[9][1][2] ,
         \ANSWER/mem[9][1][1] , \ANSWER/mem[9][1][0] , \ANSWER/mem[9][0][15] ,
         \ANSWER/mem[9][0][14] , \ANSWER/mem[9][0][13] ,
         \ANSWER/mem[9][0][12] , \ANSWER/mem[9][0][11] ,
         \ANSWER/mem[9][0][10] , \ANSWER/mem[9][0][9] , \ANSWER/mem[9][0][8] ,
         \ANSWER/mem[9][0][7] , \ANSWER/mem[9][0][6] , \ANSWER/mem[9][0][5] ,
         \ANSWER/mem[9][0][4] , \ANSWER/mem[9][0][3] , \ANSWER/mem[9][0][2] ,
         \ANSWER/mem[9][0][1] , \ANSWER/mem[9][0][0] , \ANSWER/mem[8][9][15] ,
         \ANSWER/mem[8][9][14] , \ANSWER/mem[8][9][13] ,
         \ANSWER/mem[8][9][12] , \ANSWER/mem[8][9][11] ,
         \ANSWER/mem[8][9][10] , \ANSWER/mem[8][9][9] , \ANSWER/mem[8][9][8] ,
         \ANSWER/mem[8][9][7] , \ANSWER/mem[8][9][6] , \ANSWER/mem[8][9][5] ,
         \ANSWER/mem[8][9][4] , \ANSWER/mem[8][9][3] , \ANSWER/mem[8][9][2] ,
         \ANSWER/mem[8][9][1] , \ANSWER/mem[8][9][0] , \ANSWER/mem[8][8][15] ,
         \ANSWER/mem[8][8][14] , \ANSWER/mem[8][8][13] ,
         \ANSWER/mem[8][8][12] , \ANSWER/mem[8][8][11] ,
         \ANSWER/mem[8][8][10] , \ANSWER/mem[8][8][9] , \ANSWER/mem[8][8][8] ,
         \ANSWER/mem[8][8][7] , \ANSWER/mem[8][8][6] , \ANSWER/mem[8][8][5] ,
         \ANSWER/mem[8][8][4] , \ANSWER/mem[8][8][3] , \ANSWER/mem[8][8][2] ,
         \ANSWER/mem[8][8][1] , \ANSWER/mem[8][8][0] , \ANSWER/mem[8][7][15] ,
         \ANSWER/mem[8][7][14] , \ANSWER/mem[8][7][13] ,
         \ANSWER/mem[8][7][12] , \ANSWER/mem[8][7][11] ,
         \ANSWER/mem[8][7][10] , \ANSWER/mem[8][7][9] , \ANSWER/mem[8][7][8] ,
         \ANSWER/mem[8][7][7] , \ANSWER/mem[8][7][6] , \ANSWER/mem[8][7][5] ,
         \ANSWER/mem[8][7][4] , \ANSWER/mem[8][7][3] , \ANSWER/mem[8][7][2] ,
         \ANSWER/mem[8][7][1] , \ANSWER/mem[8][7][0] , \ANSWER/mem[8][6][15] ,
         \ANSWER/mem[8][6][14] , \ANSWER/mem[8][6][13] ,
         \ANSWER/mem[8][6][12] , \ANSWER/mem[8][6][11] ,
         \ANSWER/mem[8][6][10] , \ANSWER/mem[8][6][9] , \ANSWER/mem[8][6][8] ,
         \ANSWER/mem[8][6][7] , \ANSWER/mem[8][6][6] , \ANSWER/mem[8][6][5] ,
         \ANSWER/mem[8][6][4] , \ANSWER/mem[8][6][3] , \ANSWER/mem[8][6][2] ,
         \ANSWER/mem[8][6][1] , \ANSWER/mem[8][6][0] , \ANSWER/mem[8][5][15] ,
         \ANSWER/mem[8][5][14] , \ANSWER/mem[8][5][13] ,
         \ANSWER/mem[8][5][12] , \ANSWER/mem[8][5][11] ,
         \ANSWER/mem[8][5][10] , \ANSWER/mem[8][5][9] , \ANSWER/mem[8][5][8] ,
         \ANSWER/mem[8][5][7] , \ANSWER/mem[8][5][6] , \ANSWER/mem[8][5][5] ,
         \ANSWER/mem[8][5][4] , \ANSWER/mem[8][5][3] , \ANSWER/mem[8][5][2] ,
         \ANSWER/mem[8][5][1] , \ANSWER/mem[8][5][0] , \ANSWER/mem[8][4][15] ,
         \ANSWER/mem[8][4][14] , \ANSWER/mem[8][4][13] ,
         \ANSWER/mem[8][4][12] , \ANSWER/mem[8][4][11] ,
         \ANSWER/mem[8][4][10] , \ANSWER/mem[8][4][9] , \ANSWER/mem[8][4][8] ,
         \ANSWER/mem[8][4][7] , \ANSWER/mem[8][4][6] , \ANSWER/mem[8][4][5] ,
         \ANSWER/mem[8][4][4] , \ANSWER/mem[8][4][3] , \ANSWER/mem[8][4][2] ,
         \ANSWER/mem[8][4][1] , \ANSWER/mem[8][4][0] , \ANSWER/mem[8][3][15] ,
         \ANSWER/mem[8][3][14] , \ANSWER/mem[8][3][13] ,
         \ANSWER/mem[8][3][12] , \ANSWER/mem[8][3][11] ,
         \ANSWER/mem[8][3][10] , \ANSWER/mem[8][3][9] , \ANSWER/mem[8][3][8] ,
         \ANSWER/mem[8][3][7] , \ANSWER/mem[8][3][6] , \ANSWER/mem[8][3][5] ,
         \ANSWER/mem[8][3][4] , \ANSWER/mem[8][3][3] , \ANSWER/mem[8][3][2] ,
         \ANSWER/mem[8][3][1] , \ANSWER/mem[8][3][0] , \ANSWER/mem[8][2][15] ,
         \ANSWER/mem[8][2][14] , \ANSWER/mem[8][2][13] ,
         \ANSWER/mem[8][2][12] , \ANSWER/mem[8][2][11] ,
         \ANSWER/mem[8][2][10] , \ANSWER/mem[8][2][9] , \ANSWER/mem[8][2][8] ,
         \ANSWER/mem[8][2][7] , \ANSWER/mem[8][2][6] , \ANSWER/mem[8][2][5] ,
         \ANSWER/mem[8][2][4] , \ANSWER/mem[8][2][3] , \ANSWER/mem[8][2][2] ,
         \ANSWER/mem[8][2][1] , \ANSWER/mem[8][2][0] , \ANSWER/mem[8][1][15] ,
         \ANSWER/mem[8][1][14] , \ANSWER/mem[8][1][13] ,
         \ANSWER/mem[8][1][12] , \ANSWER/mem[8][1][11] ,
         \ANSWER/mem[8][1][10] , \ANSWER/mem[8][1][9] , \ANSWER/mem[8][1][8] ,
         \ANSWER/mem[8][1][7] , \ANSWER/mem[8][1][6] , \ANSWER/mem[8][1][5] ,
         \ANSWER/mem[8][1][4] , \ANSWER/mem[8][1][3] , \ANSWER/mem[8][1][2] ,
         \ANSWER/mem[8][1][1] , \ANSWER/mem[8][1][0] , \ANSWER/mem[8][0][15] ,
         \ANSWER/mem[8][0][14] , \ANSWER/mem[8][0][13] ,
         \ANSWER/mem[8][0][12] , \ANSWER/mem[8][0][11] ,
         \ANSWER/mem[8][0][10] , \ANSWER/mem[8][0][9] , \ANSWER/mem[8][0][8] ,
         \ANSWER/mem[8][0][7] , \ANSWER/mem[8][0][6] , \ANSWER/mem[8][0][5] ,
         \ANSWER/mem[8][0][4] , \ANSWER/mem[8][0][3] , \ANSWER/mem[8][0][2] ,
         \ANSWER/mem[8][0][1] , \ANSWER/mem[8][0][0] , \ANSWER/mem[7][9][15] ,
         \ANSWER/mem[7][9][14] , \ANSWER/mem[7][9][13] ,
         \ANSWER/mem[7][9][12] , \ANSWER/mem[7][9][11] ,
         \ANSWER/mem[7][9][10] , \ANSWER/mem[7][9][9] , \ANSWER/mem[7][9][8] ,
         \ANSWER/mem[7][9][7] , \ANSWER/mem[7][9][6] , \ANSWER/mem[7][9][5] ,
         \ANSWER/mem[7][9][4] , \ANSWER/mem[7][9][3] , \ANSWER/mem[7][9][2] ,
         \ANSWER/mem[7][9][1] , \ANSWER/mem[7][9][0] , \ANSWER/mem[7][8][15] ,
         \ANSWER/mem[7][8][14] , \ANSWER/mem[7][8][13] ,
         \ANSWER/mem[7][8][12] , \ANSWER/mem[7][8][11] ,
         \ANSWER/mem[7][8][10] , \ANSWER/mem[7][8][9] , \ANSWER/mem[7][8][8] ,
         \ANSWER/mem[7][8][7] , \ANSWER/mem[7][8][6] , \ANSWER/mem[7][8][5] ,
         \ANSWER/mem[7][8][4] , \ANSWER/mem[7][8][3] , \ANSWER/mem[7][8][2] ,
         \ANSWER/mem[7][8][1] , \ANSWER/mem[7][8][0] , \ANSWER/mem[7][7][15] ,
         \ANSWER/mem[7][7][14] , \ANSWER/mem[7][7][13] ,
         \ANSWER/mem[7][7][12] , \ANSWER/mem[7][7][11] ,
         \ANSWER/mem[7][7][10] , \ANSWER/mem[7][7][9] , \ANSWER/mem[7][7][8] ,
         \ANSWER/mem[7][7][7] , \ANSWER/mem[7][7][6] , \ANSWER/mem[7][7][5] ,
         \ANSWER/mem[7][7][4] , \ANSWER/mem[7][7][3] , \ANSWER/mem[7][7][2] ,
         \ANSWER/mem[7][7][1] , \ANSWER/mem[7][7][0] , \ANSWER/mem[7][6][15] ,
         \ANSWER/mem[7][6][14] , \ANSWER/mem[7][6][13] ,
         \ANSWER/mem[7][6][12] , \ANSWER/mem[7][6][11] ,
         \ANSWER/mem[7][6][10] , \ANSWER/mem[7][6][9] , \ANSWER/mem[7][6][8] ,
         \ANSWER/mem[7][6][7] , \ANSWER/mem[7][6][6] , \ANSWER/mem[7][6][5] ,
         \ANSWER/mem[7][6][4] , \ANSWER/mem[7][6][3] , \ANSWER/mem[7][6][2] ,
         \ANSWER/mem[7][6][1] , \ANSWER/mem[7][6][0] , \ANSWER/mem[7][5][15] ,
         \ANSWER/mem[7][5][14] , \ANSWER/mem[7][5][13] ,
         \ANSWER/mem[7][5][12] , \ANSWER/mem[7][5][11] ,
         \ANSWER/mem[7][5][10] , \ANSWER/mem[7][5][9] , \ANSWER/mem[7][5][8] ,
         \ANSWER/mem[7][5][7] , \ANSWER/mem[7][5][6] , \ANSWER/mem[7][5][5] ,
         \ANSWER/mem[7][5][4] , \ANSWER/mem[7][5][3] , \ANSWER/mem[7][5][2] ,
         \ANSWER/mem[7][5][1] , \ANSWER/mem[7][5][0] , \ANSWER/mem[7][4][15] ,
         \ANSWER/mem[7][4][14] , \ANSWER/mem[7][4][13] ,
         \ANSWER/mem[7][4][12] , \ANSWER/mem[7][4][11] ,
         \ANSWER/mem[7][4][10] , \ANSWER/mem[7][4][9] , \ANSWER/mem[7][4][8] ,
         \ANSWER/mem[7][4][7] , \ANSWER/mem[7][4][6] , \ANSWER/mem[7][4][5] ,
         \ANSWER/mem[7][4][4] , \ANSWER/mem[7][4][3] , \ANSWER/mem[7][4][2] ,
         \ANSWER/mem[7][4][1] , \ANSWER/mem[7][4][0] , \ANSWER/mem[7][3][15] ,
         \ANSWER/mem[7][3][14] , \ANSWER/mem[7][3][13] ,
         \ANSWER/mem[7][3][12] , \ANSWER/mem[7][3][11] ,
         \ANSWER/mem[7][3][10] , \ANSWER/mem[7][3][9] , \ANSWER/mem[7][3][8] ,
         \ANSWER/mem[7][3][7] , \ANSWER/mem[7][3][6] , \ANSWER/mem[7][3][5] ,
         \ANSWER/mem[7][3][4] , \ANSWER/mem[7][3][3] , \ANSWER/mem[7][3][2] ,
         \ANSWER/mem[7][3][1] , \ANSWER/mem[7][3][0] , \ANSWER/mem[7][2][15] ,
         \ANSWER/mem[7][2][14] , \ANSWER/mem[7][2][13] ,
         \ANSWER/mem[7][2][12] , \ANSWER/mem[7][2][11] ,
         \ANSWER/mem[7][2][10] , \ANSWER/mem[7][2][9] , \ANSWER/mem[7][2][8] ,
         \ANSWER/mem[7][2][7] , \ANSWER/mem[7][2][6] , \ANSWER/mem[7][2][5] ,
         \ANSWER/mem[7][2][4] , \ANSWER/mem[7][2][3] , \ANSWER/mem[7][2][2] ,
         \ANSWER/mem[7][2][1] , \ANSWER/mem[7][2][0] , \ANSWER/mem[7][1][15] ,
         \ANSWER/mem[7][1][14] , \ANSWER/mem[7][1][13] ,
         \ANSWER/mem[7][1][12] , \ANSWER/mem[7][1][11] ,
         \ANSWER/mem[7][1][10] , \ANSWER/mem[7][1][9] , \ANSWER/mem[7][1][8] ,
         \ANSWER/mem[7][1][7] , \ANSWER/mem[7][1][6] , \ANSWER/mem[7][1][5] ,
         \ANSWER/mem[7][1][4] , \ANSWER/mem[7][1][3] , \ANSWER/mem[7][1][2] ,
         \ANSWER/mem[7][1][1] , \ANSWER/mem[7][1][0] , \ANSWER/mem[7][0][15] ,
         \ANSWER/mem[7][0][14] , \ANSWER/mem[7][0][13] ,
         \ANSWER/mem[7][0][12] , \ANSWER/mem[7][0][11] ,
         \ANSWER/mem[7][0][10] , \ANSWER/mem[7][0][9] , \ANSWER/mem[7][0][8] ,
         \ANSWER/mem[7][0][7] , \ANSWER/mem[7][0][6] , \ANSWER/mem[7][0][5] ,
         \ANSWER/mem[7][0][4] , \ANSWER/mem[7][0][3] , \ANSWER/mem[7][0][2] ,
         \ANSWER/mem[7][0][1] , \ANSWER/mem[7][0][0] , \ANSWER/mem[6][9][15] ,
         \ANSWER/mem[6][9][14] , \ANSWER/mem[6][9][13] ,
         \ANSWER/mem[6][9][12] , \ANSWER/mem[6][9][11] ,
         \ANSWER/mem[6][9][10] , \ANSWER/mem[6][9][9] , \ANSWER/mem[6][9][8] ,
         \ANSWER/mem[6][9][7] , \ANSWER/mem[6][9][6] , \ANSWER/mem[6][9][5] ,
         \ANSWER/mem[6][9][4] , \ANSWER/mem[6][9][3] , \ANSWER/mem[6][9][2] ,
         \ANSWER/mem[6][9][1] , \ANSWER/mem[6][9][0] , \ANSWER/mem[6][8][15] ,
         \ANSWER/mem[6][8][14] , \ANSWER/mem[6][8][13] ,
         \ANSWER/mem[6][8][12] , \ANSWER/mem[6][8][11] ,
         \ANSWER/mem[6][8][10] , \ANSWER/mem[6][8][9] , \ANSWER/mem[6][8][8] ,
         \ANSWER/mem[6][8][7] , \ANSWER/mem[6][8][6] , \ANSWER/mem[6][8][5] ,
         \ANSWER/mem[6][8][4] , \ANSWER/mem[6][8][3] , \ANSWER/mem[6][8][2] ,
         \ANSWER/mem[6][8][1] , \ANSWER/mem[6][8][0] , \ANSWER/mem[6][7][15] ,
         \ANSWER/mem[6][7][14] , \ANSWER/mem[6][7][13] ,
         \ANSWER/mem[6][7][12] , \ANSWER/mem[6][7][11] ,
         \ANSWER/mem[6][7][10] , \ANSWER/mem[6][7][9] , \ANSWER/mem[6][7][8] ,
         \ANSWER/mem[6][7][7] , \ANSWER/mem[6][7][6] , \ANSWER/mem[6][7][5] ,
         \ANSWER/mem[6][7][4] , \ANSWER/mem[6][7][3] , \ANSWER/mem[6][7][2] ,
         \ANSWER/mem[6][7][1] , \ANSWER/mem[6][7][0] , \ANSWER/mem[6][6][15] ,
         \ANSWER/mem[6][6][14] , \ANSWER/mem[6][6][13] ,
         \ANSWER/mem[6][6][12] , \ANSWER/mem[6][6][11] ,
         \ANSWER/mem[6][6][10] , \ANSWER/mem[6][6][9] , \ANSWER/mem[6][6][8] ,
         \ANSWER/mem[6][6][7] , \ANSWER/mem[6][6][6] , \ANSWER/mem[6][6][5] ,
         \ANSWER/mem[6][6][4] , \ANSWER/mem[6][6][3] , \ANSWER/mem[6][6][2] ,
         \ANSWER/mem[6][6][1] , \ANSWER/mem[6][6][0] , \ANSWER/mem[6][5][15] ,
         \ANSWER/mem[6][5][14] , \ANSWER/mem[6][5][13] ,
         \ANSWER/mem[6][5][12] , \ANSWER/mem[6][5][11] ,
         \ANSWER/mem[6][5][10] , \ANSWER/mem[6][5][9] , \ANSWER/mem[6][5][8] ,
         \ANSWER/mem[6][5][7] , \ANSWER/mem[6][5][6] , \ANSWER/mem[6][5][5] ,
         \ANSWER/mem[6][5][4] , \ANSWER/mem[6][5][3] , \ANSWER/mem[6][5][2] ,
         \ANSWER/mem[6][5][1] , \ANSWER/mem[6][5][0] , \ANSWER/mem[6][4][15] ,
         \ANSWER/mem[6][4][14] , \ANSWER/mem[6][4][13] ,
         \ANSWER/mem[6][4][12] , \ANSWER/mem[6][4][11] ,
         \ANSWER/mem[6][4][10] , \ANSWER/mem[6][4][9] , \ANSWER/mem[6][4][8] ,
         \ANSWER/mem[6][4][7] , \ANSWER/mem[6][4][6] , \ANSWER/mem[6][4][5] ,
         \ANSWER/mem[6][4][4] , \ANSWER/mem[6][4][3] , \ANSWER/mem[6][4][2] ,
         \ANSWER/mem[6][4][1] , \ANSWER/mem[6][4][0] , \ANSWER/mem[6][3][15] ,
         \ANSWER/mem[6][3][14] , \ANSWER/mem[6][3][13] ,
         \ANSWER/mem[6][3][12] , \ANSWER/mem[6][3][11] ,
         \ANSWER/mem[6][3][10] , \ANSWER/mem[6][3][9] , \ANSWER/mem[6][3][8] ,
         \ANSWER/mem[6][3][7] , \ANSWER/mem[6][3][6] , \ANSWER/mem[6][3][5] ,
         \ANSWER/mem[6][3][4] , \ANSWER/mem[6][3][3] , \ANSWER/mem[6][3][2] ,
         \ANSWER/mem[6][3][1] , \ANSWER/mem[6][3][0] , \ANSWER/mem[6][2][15] ,
         \ANSWER/mem[6][2][14] , \ANSWER/mem[6][2][13] ,
         \ANSWER/mem[6][2][12] , \ANSWER/mem[6][2][11] ,
         \ANSWER/mem[6][2][10] , \ANSWER/mem[6][2][9] , \ANSWER/mem[6][2][8] ,
         \ANSWER/mem[6][2][7] , \ANSWER/mem[6][2][6] , \ANSWER/mem[6][2][5] ,
         \ANSWER/mem[6][2][4] , \ANSWER/mem[6][2][3] , \ANSWER/mem[6][2][2] ,
         \ANSWER/mem[6][2][1] , \ANSWER/mem[6][2][0] , \ANSWER/mem[6][1][15] ,
         \ANSWER/mem[6][1][14] , \ANSWER/mem[6][1][13] ,
         \ANSWER/mem[6][1][12] , \ANSWER/mem[6][1][11] ,
         \ANSWER/mem[6][1][10] , \ANSWER/mem[6][1][9] , \ANSWER/mem[6][1][8] ,
         \ANSWER/mem[6][1][7] , \ANSWER/mem[6][1][6] , \ANSWER/mem[6][1][5] ,
         \ANSWER/mem[6][1][4] , \ANSWER/mem[6][1][3] , \ANSWER/mem[6][1][2] ,
         \ANSWER/mem[6][1][1] , \ANSWER/mem[6][1][0] , \ANSWER/mem[6][0][15] ,
         \ANSWER/mem[6][0][14] , \ANSWER/mem[6][0][13] ,
         \ANSWER/mem[6][0][12] , \ANSWER/mem[6][0][11] ,
         \ANSWER/mem[6][0][10] , \ANSWER/mem[6][0][9] , \ANSWER/mem[6][0][8] ,
         \ANSWER/mem[6][0][7] , \ANSWER/mem[6][0][6] , \ANSWER/mem[6][0][5] ,
         \ANSWER/mem[6][0][4] , \ANSWER/mem[6][0][3] , \ANSWER/mem[6][0][2] ,
         \ANSWER/mem[6][0][1] , \ANSWER/mem[6][0][0] , \ANSWER/mem[5][9][15] ,
         \ANSWER/mem[5][9][14] , \ANSWER/mem[5][9][13] ,
         \ANSWER/mem[5][9][12] , \ANSWER/mem[5][9][11] ,
         \ANSWER/mem[5][9][10] , \ANSWER/mem[5][9][9] , \ANSWER/mem[5][9][8] ,
         \ANSWER/mem[5][9][7] , \ANSWER/mem[5][9][6] , \ANSWER/mem[5][9][5] ,
         \ANSWER/mem[5][9][4] , \ANSWER/mem[5][9][3] , \ANSWER/mem[5][9][2] ,
         \ANSWER/mem[5][9][1] , \ANSWER/mem[5][9][0] , \ANSWER/mem[5][8][15] ,
         \ANSWER/mem[5][8][14] , \ANSWER/mem[5][8][13] ,
         \ANSWER/mem[5][8][12] , \ANSWER/mem[5][8][11] ,
         \ANSWER/mem[5][8][10] , \ANSWER/mem[5][8][9] , \ANSWER/mem[5][8][8] ,
         \ANSWER/mem[5][8][7] , \ANSWER/mem[5][8][6] , \ANSWER/mem[5][8][5] ,
         \ANSWER/mem[5][8][4] , \ANSWER/mem[5][8][3] , \ANSWER/mem[5][8][2] ,
         \ANSWER/mem[5][8][1] , \ANSWER/mem[5][8][0] , \ANSWER/mem[5][7][15] ,
         \ANSWER/mem[5][7][14] , \ANSWER/mem[5][7][13] ,
         \ANSWER/mem[5][7][12] , \ANSWER/mem[5][7][11] ,
         \ANSWER/mem[5][7][10] , \ANSWER/mem[5][7][9] , \ANSWER/mem[5][7][8] ,
         \ANSWER/mem[5][7][7] , \ANSWER/mem[5][7][6] , \ANSWER/mem[5][7][5] ,
         \ANSWER/mem[5][7][4] , \ANSWER/mem[5][7][3] , \ANSWER/mem[5][7][2] ,
         \ANSWER/mem[5][7][1] , \ANSWER/mem[5][7][0] , \ANSWER/mem[5][6][15] ,
         \ANSWER/mem[5][6][14] , \ANSWER/mem[5][6][13] ,
         \ANSWER/mem[5][6][12] , \ANSWER/mem[5][6][11] ,
         \ANSWER/mem[5][6][10] , \ANSWER/mem[5][6][9] , \ANSWER/mem[5][6][8] ,
         \ANSWER/mem[5][6][7] , \ANSWER/mem[5][6][6] , \ANSWER/mem[5][6][5] ,
         \ANSWER/mem[5][6][4] , \ANSWER/mem[5][6][3] , \ANSWER/mem[5][6][2] ,
         \ANSWER/mem[5][6][1] , \ANSWER/mem[5][6][0] , \ANSWER/mem[5][5][15] ,
         \ANSWER/mem[5][5][14] , \ANSWER/mem[5][5][13] ,
         \ANSWER/mem[5][5][12] , \ANSWER/mem[5][5][11] ,
         \ANSWER/mem[5][5][10] , \ANSWER/mem[5][5][9] , \ANSWER/mem[5][5][8] ,
         \ANSWER/mem[5][5][7] , \ANSWER/mem[5][5][6] , \ANSWER/mem[5][5][5] ,
         \ANSWER/mem[5][5][4] , \ANSWER/mem[5][5][3] , \ANSWER/mem[5][5][2] ,
         \ANSWER/mem[5][5][1] , \ANSWER/mem[5][5][0] , \ANSWER/mem[5][4][15] ,
         \ANSWER/mem[5][4][14] , \ANSWER/mem[5][4][13] ,
         \ANSWER/mem[5][4][12] , \ANSWER/mem[5][4][11] ,
         \ANSWER/mem[5][4][10] , \ANSWER/mem[5][4][9] , \ANSWER/mem[5][4][8] ,
         \ANSWER/mem[5][4][7] , \ANSWER/mem[5][4][6] , \ANSWER/mem[5][4][5] ,
         \ANSWER/mem[5][4][4] , \ANSWER/mem[5][4][3] , \ANSWER/mem[5][4][2] ,
         \ANSWER/mem[5][4][1] , \ANSWER/mem[5][4][0] , \ANSWER/mem[5][3][15] ,
         \ANSWER/mem[5][3][14] , \ANSWER/mem[5][3][13] ,
         \ANSWER/mem[5][3][12] , \ANSWER/mem[5][3][11] ,
         \ANSWER/mem[5][3][10] , \ANSWER/mem[5][3][9] , \ANSWER/mem[5][3][8] ,
         \ANSWER/mem[5][3][7] , \ANSWER/mem[5][3][6] , \ANSWER/mem[5][3][5] ,
         \ANSWER/mem[5][3][4] , \ANSWER/mem[5][3][3] , \ANSWER/mem[5][3][2] ,
         \ANSWER/mem[5][3][1] , \ANSWER/mem[5][3][0] , \ANSWER/mem[5][2][15] ,
         \ANSWER/mem[5][2][14] , \ANSWER/mem[5][2][13] ,
         \ANSWER/mem[5][2][12] , \ANSWER/mem[5][2][11] ,
         \ANSWER/mem[5][2][10] , \ANSWER/mem[5][2][9] , \ANSWER/mem[5][2][8] ,
         \ANSWER/mem[5][2][7] , \ANSWER/mem[5][2][6] , \ANSWER/mem[5][2][5] ,
         \ANSWER/mem[5][2][4] , \ANSWER/mem[5][2][3] , \ANSWER/mem[5][2][2] ,
         \ANSWER/mem[5][2][1] , \ANSWER/mem[5][2][0] , \ANSWER/mem[5][1][15] ,
         \ANSWER/mem[5][1][14] , \ANSWER/mem[5][1][13] ,
         \ANSWER/mem[5][1][12] , \ANSWER/mem[5][1][11] ,
         \ANSWER/mem[5][1][10] , \ANSWER/mem[5][1][9] , \ANSWER/mem[5][1][8] ,
         \ANSWER/mem[5][1][7] , \ANSWER/mem[5][1][6] , \ANSWER/mem[5][1][5] ,
         \ANSWER/mem[5][1][4] , \ANSWER/mem[5][1][3] , \ANSWER/mem[5][1][2] ,
         \ANSWER/mem[5][1][1] , \ANSWER/mem[5][1][0] , \ANSWER/mem[5][0][15] ,
         \ANSWER/mem[5][0][14] , \ANSWER/mem[5][0][13] ,
         \ANSWER/mem[5][0][12] , \ANSWER/mem[5][0][11] ,
         \ANSWER/mem[5][0][10] , \ANSWER/mem[5][0][9] , \ANSWER/mem[5][0][8] ,
         \ANSWER/mem[5][0][7] , \ANSWER/mem[5][0][6] , \ANSWER/mem[5][0][5] ,
         \ANSWER/mem[5][0][4] , \ANSWER/mem[5][0][3] , \ANSWER/mem[5][0][2] ,
         \ANSWER/mem[5][0][1] , \ANSWER/mem[5][0][0] , \ANSWER/mem[4][9][15] ,
         \ANSWER/mem[4][9][14] , \ANSWER/mem[4][9][13] ,
         \ANSWER/mem[4][9][12] , \ANSWER/mem[4][9][11] ,
         \ANSWER/mem[4][9][10] , \ANSWER/mem[4][9][9] , \ANSWER/mem[4][9][8] ,
         \ANSWER/mem[4][9][7] , \ANSWER/mem[4][9][6] , \ANSWER/mem[4][9][5] ,
         \ANSWER/mem[4][9][4] , \ANSWER/mem[4][9][3] , \ANSWER/mem[4][9][2] ,
         \ANSWER/mem[4][9][1] , \ANSWER/mem[4][9][0] , \ANSWER/mem[4][8][15] ,
         \ANSWER/mem[4][8][14] , \ANSWER/mem[4][8][13] ,
         \ANSWER/mem[4][8][12] , \ANSWER/mem[4][8][11] ,
         \ANSWER/mem[4][8][10] , \ANSWER/mem[4][8][9] , \ANSWER/mem[4][8][8] ,
         \ANSWER/mem[4][8][7] , \ANSWER/mem[4][8][6] , \ANSWER/mem[4][8][5] ,
         \ANSWER/mem[4][8][4] , \ANSWER/mem[4][8][3] , \ANSWER/mem[4][8][2] ,
         \ANSWER/mem[4][8][1] , \ANSWER/mem[4][8][0] , \ANSWER/mem[4][7][15] ,
         \ANSWER/mem[4][7][14] , \ANSWER/mem[4][7][13] ,
         \ANSWER/mem[4][7][12] , \ANSWER/mem[4][7][11] ,
         \ANSWER/mem[4][7][10] , \ANSWER/mem[4][7][9] , \ANSWER/mem[4][7][8] ,
         \ANSWER/mem[4][7][7] , \ANSWER/mem[4][7][6] , \ANSWER/mem[4][7][5] ,
         \ANSWER/mem[4][7][4] , \ANSWER/mem[4][7][3] , \ANSWER/mem[4][7][2] ,
         \ANSWER/mem[4][7][1] , \ANSWER/mem[4][7][0] , \ANSWER/mem[4][6][15] ,
         \ANSWER/mem[4][6][14] , \ANSWER/mem[4][6][13] ,
         \ANSWER/mem[4][6][12] , \ANSWER/mem[4][6][11] ,
         \ANSWER/mem[4][6][10] , \ANSWER/mem[4][6][9] , \ANSWER/mem[4][6][8] ,
         \ANSWER/mem[4][6][7] , \ANSWER/mem[4][6][6] , \ANSWER/mem[4][6][5] ,
         \ANSWER/mem[4][6][4] , \ANSWER/mem[4][6][3] , \ANSWER/mem[4][6][2] ,
         \ANSWER/mem[4][6][1] , \ANSWER/mem[4][6][0] , \ANSWER/mem[4][5][15] ,
         \ANSWER/mem[4][5][14] , \ANSWER/mem[4][5][13] ,
         \ANSWER/mem[4][5][12] , \ANSWER/mem[4][5][11] ,
         \ANSWER/mem[4][5][10] , \ANSWER/mem[4][5][9] , \ANSWER/mem[4][5][8] ,
         \ANSWER/mem[4][5][7] , \ANSWER/mem[4][5][6] , \ANSWER/mem[4][5][5] ,
         \ANSWER/mem[4][5][4] , \ANSWER/mem[4][5][3] , \ANSWER/mem[4][5][2] ,
         \ANSWER/mem[4][5][1] , \ANSWER/mem[4][5][0] , \ANSWER/mem[4][4][15] ,
         \ANSWER/mem[4][4][14] , \ANSWER/mem[4][4][13] ,
         \ANSWER/mem[4][4][12] , \ANSWER/mem[4][4][11] ,
         \ANSWER/mem[4][4][10] , \ANSWER/mem[4][4][9] , \ANSWER/mem[4][4][8] ,
         \ANSWER/mem[4][4][7] , \ANSWER/mem[4][4][6] , \ANSWER/mem[4][4][5] ,
         \ANSWER/mem[4][4][4] , \ANSWER/mem[4][4][3] , \ANSWER/mem[4][4][2] ,
         \ANSWER/mem[4][4][1] , \ANSWER/mem[4][4][0] , \ANSWER/mem[4][3][15] ,
         \ANSWER/mem[4][3][14] , \ANSWER/mem[4][3][13] ,
         \ANSWER/mem[4][3][12] , \ANSWER/mem[4][3][11] ,
         \ANSWER/mem[4][3][10] , \ANSWER/mem[4][3][9] , \ANSWER/mem[4][3][8] ,
         \ANSWER/mem[4][3][7] , \ANSWER/mem[4][3][6] , \ANSWER/mem[4][3][5] ,
         \ANSWER/mem[4][3][4] , \ANSWER/mem[4][3][3] , \ANSWER/mem[4][3][2] ,
         \ANSWER/mem[4][3][1] , \ANSWER/mem[4][3][0] , \ANSWER/mem[4][2][15] ,
         \ANSWER/mem[4][2][14] , \ANSWER/mem[4][2][13] ,
         \ANSWER/mem[4][2][12] , \ANSWER/mem[4][2][11] ,
         \ANSWER/mem[4][2][10] , \ANSWER/mem[4][2][9] , \ANSWER/mem[4][2][8] ,
         \ANSWER/mem[4][2][7] , \ANSWER/mem[4][2][6] , \ANSWER/mem[4][2][5] ,
         \ANSWER/mem[4][2][4] , \ANSWER/mem[4][2][3] , \ANSWER/mem[4][2][2] ,
         \ANSWER/mem[4][2][1] , \ANSWER/mem[4][2][0] , \ANSWER/mem[4][1][15] ,
         \ANSWER/mem[4][1][14] , \ANSWER/mem[4][1][13] ,
         \ANSWER/mem[4][1][12] , \ANSWER/mem[4][1][11] ,
         \ANSWER/mem[4][1][10] , \ANSWER/mem[4][1][9] , \ANSWER/mem[4][1][8] ,
         \ANSWER/mem[4][1][7] , \ANSWER/mem[4][1][6] , \ANSWER/mem[4][1][5] ,
         \ANSWER/mem[4][1][4] , \ANSWER/mem[4][1][3] , \ANSWER/mem[4][1][2] ,
         \ANSWER/mem[4][1][1] , \ANSWER/mem[4][1][0] , \ANSWER/mem[4][0][15] ,
         \ANSWER/mem[4][0][14] , \ANSWER/mem[4][0][13] ,
         \ANSWER/mem[4][0][12] , \ANSWER/mem[4][0][11] ,
         \ANSWER/mem[4][0][10] , \ANSWER/mem[4][0][9] , \ANSWER/mem[4][0][8] ,
         \ANSWER/mem[4][0][7] , \ANSWER/mem[4][0][6] , \ANSWER/mem[4][0][5] ,
         \ANSWER/mem[4][0][4] , \ANSWER/mem[4][0][3] , \ANSWER/mem[4][0][2] ,
         \ANSWER/mem[4][0][1] , \ANSWER/mem[4][0][0] , \ANSWER/mem[3][9][15] ,
         \ANSWER/mem[3][9][14] , \ANSWER/mem[3][9][13] ,
         \ANSWER/mem[3][9][12] , \ANSWER/mem[3][9][11] ,
         \ANSWER/mem[3][9][10] , \ANSWER/mem[3][9][9] , \ANSWER/mem[3][9][8] ,
         \ANSWER/mem[3][9][7] , \ANSWER/mem[3][9][6] , \ANSWER/mem[3][9][5] ,
         \ANSWER/mem[3][9][4] , \ANSWER/mem[3][9][3] , \ANSWER/mem[3][9][2] ,
         \ANSWER/mem[3][9][1] , \ANSWER/mem[3][9][0] , \ANSWER/mem[3][8][15] ,
         \ANSWER/mem[3][8][14] , \ANSWER/mem[3][8][13] ,
         \ANSWER/mem[3][8][12] , \ANSWER/mem[3][8][11] ,
         \ANSWER/mem[3][8][10] , \ANSWER/mem[3][8][9] , \ANSWER/mem[3][8][8] ,
         \ANSWER/mem[3][8][7] , \ANSWER/mem[3][8][6] , \ANSWER/mem[3][8][5] ,
         \ANSWER/mem[3][8][4] , \ANSWER/mem[3][8][3] , \ANSWER/mem[3][8][2] ,
         \ANSWER/mem[3][8][1] , \ANSWER/mem[3][8][0] , \ANSWER/mem[3][7][15] ,
         \ANSWER/mem[3][7][14] , \ANSWER/mem[3][7][13] ,
         \ANSWER/mem[3][7][12] , \ANSWER/mem[3][7][11] ,
         \ANSWER/mem[3][7][10] , \ANSWER/mem[3][7][9] , \ANSWER/mem[3][7][8] ,
         \ANSWER/mem[3][7][7] , \ANSWER/mem[3][7][6] , \ANSWER/mem[3][7][5] ,
         \ANSWER/mem[3][7][4] , \ANSWER/mem[3][7][3] , \ANSWER/mem[3][7][2] ,
         \ANSWER/mem[3][7][1] , \ANSWER/mem[3][7][0] , \ANSWER/mem[3][6][15] ,
         \ANSWER/mem[3][6][14] , \ANSWER/mem[3][6][13] ,
         \ANSWER/mem[3][6][12] , \ANSWER/mem[3][6][11] ,
         \ANSWER/mem[3][6][10] , \ANSWER/mem[3][6][9] , \ANSWER/mem[3][6][8] ,
         \ANSWER/mem[3][6][7] , \ANSWER/mem[3][6][6] , \ANSWER/mem[3][6][5] ,
         \ANSWER/mem[3][6][4] , \ANSWER/mem[3][6][3] , \ANSWER/mem[3][6][2] ,
         \ANSWER/mem[3][6][1] , \ANSWER/mem[3][6][0] , \ANSWER/mem[3][5][15] ,
         \ANSWER/mem[3][5][14] , \ANSWER/mem[3][5][13] ,
         \ANSWER/mem[3][5][12] , \ANSWER/mem[3][5][11] ,
         \ANSWER/mem[3][5][10] , \ANSWER/mem[3][5][9] , \ANSWER/mem[3][5][8] ,
         \ANSWER/mem[3][5][7] , \ANSWER/mem[3][5][6] , \ANSWER/mem[3][5][5] ,
         \ANSWER/mem[3][5][4] , \ANSWER/mem[3][5][3] , \ANSWER/mem[3][5][2] ,
         \ANSWER/mem[3][5][1] , \ANSWER/mem[3][5][0] , \ANSWER/mem[3][4][15] ,
         \ANSWER/mem[3][4][14] , \ANSWER/mem[3][4][13] ,
         \ANSWER/mem[3][4][12] , \ANSWER/mem[3][4][11] ,
         \ANSWER/mem[3][4][10] , \ANSWER/mem[3][4][9] , \ANSWER/mem[3][4][8] ,
         \ANSWER/mem[3][4][7] , \ANSWER/mem[3][4][6] , \ANSWER/mem[3][4][5] ,
         \ANSWER/mem[3][4][4] , \ANSWER/mem[3][4][3] , \ANSWER/mem[3][4][2] ,
         \ANSWER/mem[3][4][1] , \ANSWER/mem[3][4][0] , \ANSWER/mem[3][3][15] ,
         \ANSWER/mem[3][3][14] , \ANSWER/mem[3][3][13] ,
         \ANSWER/mem[3][3][12] , \ANSWER/mem[3][3][11] ,
         \ANSWER/mem[3][3][10] , \ANSWER/mem[3][3][9] , \ANSWER/mem[3][3][8] ,
         \ANSWER/mem[3][3][7] , \ANSWER/mem[3][3][6] , \ANSWER/mem[3][3][5] ,
         \ANSWER/mem[3][3][4] , \ANSWER/mem[3][3][3] , \ANSWER/mem[3][3][2] ,
         \ANSWER/mem[3][3][1] , \ANSWER/mem[3][3][0] , \ANSWER/mem[3][2][15] ,
         \ANSWER/mem[3][2][14] , \ANSWER/mem[3][2][13] ,
         \ANSWER/mem[3][2][12] , \ANSWER/mem[3][2][11] ,
         \ANSWER/mem[3][2][10] , \ANSWER/mem[3][2][9] , \ANSWER/mem[3][2][8] ,
         \ANSWER/mem[3][2][7] , \ANSWER/mem[3][2][6] , \ANSWER/mem[3][2][5] ,
         \ANSWER/mem[3][2][4] , \ANSWER/mem[3][2][3] , \ANSWER/mem[3][2][2] ,
         \ANSWER/mem[3][2][1] , \ANSWER/mem[3][2][0] , \ANSWER/mem[3][1][15] ,
         \ANSWER/mem[3][1][14] , \ANSWER/mem[3][1][13] ,
         \ANSWER/mem[3][1][12] , \ANSWER/mem[3][1][11] ,
         \ANSWER/mem[3][1][10] , \ANSWER/mem[3][1][9] , \ANSWER/mem[3][1][8] ,
         \ANSWER/mem[3][1][7] , \ANSWER/mem[3][1][6] , \ANSWER/mem[3][1][5] ,
         \ANSWER/mem[3][1][4] , \ANSWER/mem[3][1][3] , \ANSWER/mem[3][1][2] ,
         \ANSWER/mem[3][1][1] , \ANSWER/mem[3][1][0] , \ANSWER/mem[3][0][15] ,
         \ANSWER/mem[3][0][14] , \ANSWER/mem[3][0][13] ,
         \ANSWER/mem[3][0][12] , \ANSWER/mem[3][0][11] ,
         \ANSWER/mem[3][0][10] , \ANSWER/mem[3][0][9] , \ANSWER/mem[3][0][8] ,
         \ANSWER/mem[3][0][7] , \ANSWER/mem[3][0][6] , \ANSWER/mem[3][0][5] ,
         \ANSWER/mem[3][0][4] , \ANSWER/mem[3][0][3] , \ANSWER/mem[3][0][2] ,
         \ANSWER/mem[3][0][1] , \ANSWER/mem[3][0][0] , \ANSWER/mem[2][9][15] ,
         \ANSWER/mem[2][9][14] , \ANSWER/mem[2][9][13] ,
         \ANSWER/mem[2][9][12] , \ANSWER/mem[2][9][11] ,
         \ANSWER/mem[2][9][10] , \ANSWER/mem[2][9][9] , \ANSWER/mem[2][9][8] ,
         \ANSWER/mem[2][9][7] , \ANSWER/mem[2][9][6] , \ANSWER/mem[2][9][5] ,
         \ANSWER/mem[2][9][4] , \ANSWER/mem[2][9][3] , \ANSWER/mem[2][9][2] ,
         \ANSWER/mem[2][9][1] , \ANSWER/mem[2][9][0] , \ANSWER/mem[2][8][15] ,
         \ANSWER/mem[2][8][14] , \ANSWER/mem[2][8][13] ,
         \ANSWER/mem[2][8][12] , \ANSWER/mem[2][8][11] ,
         \ANSWER/mem[2][8][10] , \ANSWER/mem[2][8][9] , \ANSWER/mem[2][8][8] ,
         \ANSWER/mem[2][8][7] , \ANSWER/mem[2][8][6] , \ANSWER/mem[2][8][5] ,
         \ANSWER/mem[2][8][4] , \ANSWER/mem[2][8][3] , \ANSWER/mem[2][8][2] ,
         \ANSWER/mem[2][8][1] , \ANSWER/mem[2][8][0] , \ANSWER/mem[2][7][15] ,
         \ANSWER/mem[2][7][14] , \ANSWER/mem[2][7][13] ,
         \ANSWER/mem[2][7][12] , \ANSWER/mem[2][7][11] ,
         \ANSWER/mem[2][7][10] , \ANSWER/mem[2][7][9] , \ANSWER/mem[2][7][8] ,
         \ANSWER/mem[2][7][7] , \ANSWER/mem[2][7][6] , \ANSWER/mem[2][7][5] ,
         \ANSWER/mem[2][7][4] , \ANSWER/mem[2][7][3] , \ANSWER/mem[2][7][2] ,
         \ANSWER/mem[2][7][1] , \ANSWER/mem[2][7][0] , \ANSWER/mem[2][6][15] ,
         \ANSWER/mem[2][6][14] , \ANSWER/mem[2][6][13] ,
         \ANSWER/mem[2][6][12] , \ANSWER/mem[2][6][11] ,
         \ANSWER/mem[2][6][10] , \ANSWER/mem[2][6][9] , \ANSWER/mem[2][6][8] ,
         \ANSWER/mem[2][6][7] , \ANSWER/mem[2][6][6] , \ANSWER/mem[2][6][5] ,
         \ANSWER/mem[2][6][4] , \ANSWER/mem[2][6][3] , \ANSWER/mem[2][6][2] ,
         \ANSWER/mem[2][6][1] , \ANSWER/mem[2][6][0] , \ANSWER/mem[2][5][15] ,
         \ANSWER/mem[2][5][14] , \ANSWER/mem[2][5][13] ,
         \ANSWER/mem[2][5][12] , \ANSWER/mem[2][5][11] ,
         \ANSWER/mem[2][5][10] , \ANSWER/mem[2][5][9] , \ANSWER/mem[2][5][8] ,
         \ANSWER/mem[2][5][7] , \ANSWER/mem[2][5][6] , \ANSWER/mem[2][5][5] ,
         \ANSWER/mem[2][5][4] , \ANSWER/mem[2][5][3] , \ANSWER/mem[2][5][2] ,
         \ANSWER/mem[2][5][1] , \ANSWER/mem[2][5][0] , \ANSWER/mem[2][4][15] ,
         \ANSWER/mem[2][4][14] , \ANSWER/mem[2][4][13] ,
         \ANSWER/mem[2][4][12] , \ANSWER/mem[2][4][11] ,
         \ANSWER/mem[2][4][10] , \ANSWER/mem[2][4][9] , \ANSWER/mem[2][4][8] ,
         \ANSWER/mem[2][4][7] , \ANSWER/mem[2][4][6] , \ANSWER/mem[2][4][5] ,
         \ANSWER/mem[2][4][4] , \ANSWER/mem[2][4][3] , \ANSWER/mem[2][4][2] ,
         \ANSWER/mem[2][4][1] , \ANSWER/mem[2][4][0] , \ANSWER/mem[2][3][15] ,
         \ANSWER/mem[2][3][14] , \ANSWER/mem[2][3][13] ,
         \ANSWER/mem[2][3][12] , \ANSWER/mem[2][3][11] ,
         \ANSWER/mem[2][3][10] , \ANSWER/mem[2][3][9] , \ANSWER/mem[2][3][8] ,
         \ANSWER/mem[2][3][7] , \ANSWER/mem[2][3][6] , \ANSWER/mem[2][3][5] ,
         \ANSWER/mem[2][3][4] , \ANSWER/mem[2][3][3] , \ANSWER/mem[2][3][2] ,
         \ANSWER/mem[2][3][1] , \ANSWER/mem[2][3][0] , \ANSWER/mem[2][2][15] ,
         \ANSWER/mem[2][2][14] , \ANSWER/mem[2][2][13] ,
         \ANSWER/mem[2][2][12] , \ANSWER/mem[2][2][11] ,
         \ANSWER/mem[2][2][10] , \ANSWER/mem[2][2][9] , \ANSWER/mem[2][2][8] ,
         \ANSWER/mem[2][2][7] , \ANSWER/mem[2][2][6] , \ANSWER/mem[2][2][5] ,
         \ANSWER/mem[2][2][4] , \ANSWER/mem[2][2][3] , \ANSWER/mem[2][2][2] ,
         \ANSWER/mem[2][2][1] , \ANSWER/mem[2][2][0] , \ANSWER/mem[2][1][15] ,
         \ANSWER/mem[2][1][14] , \ANSWER/mem[2][1][13] ,
         \ANSWER/mem[2][1][12] , \ANSWER/mem[2][1][11] ,
         \ANSWER/mem[2][1][10] , \ANSWER/mem[2][1][9] , \ANSWER/mem[2][1][8] ,
         \ANSWER/mem[2][1][7] , \ANSWER/mem[2][1][6] , \ANSWER/mem[2][1][5] ,
         \ANSWER/mem[2][1][4] , \ANSWER/mem[2][1][3] , \ANSWER/mem[2][1][2] ,
         \ANSWER/mem[2][1][1] , \ANSWER/mem[2][1][0] , \ANSWER/mem[2][0][15] ,
         \ANSWER/mem[2][0][14] , \ANSWER/mem[2][0][13] ,
         \ANSWER/mem[2][0][12] , \ANSWER/mem[2][0][11] ,
         \ANSWER/mem[2][0][10] , \ANSWER/mem[2][0][9] , \ANSWER/mem[2][0][8] ,
         \ANSWER/mem[2][0][7] , \ANSWER/mem[2][0][6] , \ANSWER/mem[2][0][5] ,
         \ANSWER/mem[2][0][4] , \ANSWER/mem[2][0][3] , \ANSWER/mem[2][0][2] ,
         \ANSWER/mem[2][0][1] , \ANSWER/mem[2][0][0] , \ANSWER/mem[1][9][15] ,
         \ANSWER/mem[1][9][14] , \ANSWER/mem[1][9][13] ,
         \ANSWER/mem[1][9][12] , \ANSWER/mem[1][9][11] ,
         \ANSWER/mem[1][9][10] , \ANSWER/mem[1][9][9] , \ANSWER/mem[1][9][8] ,
         \ANSWER/mem[1][9][7] , \ANSWER/mem[1][9][6] , \ANSWER/mem[1][9][5] ,
         \ANSWER/mem[1][9][4] , \ANSWER/mem[1][9][3] , \ANSWER/mem[1][9][2] ,
         \ANSWER/mem[1][9][1] , \ANSWER/mem[1][9][0] , \ANSWER/mem[1][8][15] ,
         \ANSWER/mem[1][8][14] , \ANSWER/mem[1][8][13] ,
         \ANSWER/mem[1][8][12] , \ANSWER/mem[1][8][11] ,
         \ANSWER/mem[1][8][10] , \ANSWER/mem[1][8][9] , \ANSWER/mem[1][8][8] ,
         \ANSWER/mem[1][8][7] , \ANSWER/mem[1][8][6] , \ANSWER/mem[1][8][5] ,
         \ANSWER/mem[1][8][4] , \ANSWER/mem[1][8][3] , \ANSWER/mem[1][8][2] ,
         \ANSWER/mem[1][8][1] , \ANSWER/mem[1][8][0] , \ANSWER/mem[1][7][15] ,
         \ANSWER/mem[1][7][14] , \ANSWER/mem[1][7][13] ,
         \ANSWER/mem[1][7][12] , \ANSWER/mem[1][7][11] ,
         \ANSWER/mem[1][7][10] , \ANSWER/mem[1][7][9] , \ANSWER/mem[1][7][8] ,
         \ANSWER/mem[1][7][7] , \ANSWER/mem[1][7][6] , \ANSWER/mem[1][7][5] ,
         \ANSWER/mem[1][7][4] , \ANSWER/mem[1][7][3] , \ANSWER/mem[1][7][2] ,
         \ANSWER/mem[1][7][1] , \ANSWER/mem[1][7][0] , \ANSWER/mem[1][6][15] ,
         \ANSWER/mem[1][6][14] , \ANSWER/mem[1][6][13] ,
         \ANSWER/mem[1][6][12] , \ANSWER/mem[1][6][11] ,
         \ANSWER/mem[1][6][10] , \ANSWER/mem[1][6][9] , \ANSWER/mem[1][6][8] ,
         \ANSWER/mem[1][6][7] , \ANSWER/mem[1][6][6] , \ANSWER/mem[1][6][5] ,
         \ANSWER/mem[1][6][4] , \ANSWER/mem[1][6][3] , \ANSWER/mem[1][6][2] ,
         \ANSWER/mem[1][6][1] , \ANSWER/mem[1][6][0] , \ANSWER/mem[1][5][15] ,
         \ANSWER/mem[1][5][14] , \ANSWER/mem[1][5][13] ,
         \ANSWER/mem[1][5][12] , \ANSWER/mem[1][5][11] ,
         \ANSWER/mem[1][5][10] , \ANSWER/mem[1][5][9] , \ANSWER/mem[1][5][8] ,
         \ANSWER/mem[1][5][7] , \ANSWER/mem[1][5][6] , \ANSWER/mem[1][5][5] ,
         \ANSWER/mem[1][5][4] , \ANSWER/mem[1][5][3] , \ANSWER/mem[1][5][2] ,
         \ANSWER/mem[1][5][1] , \ANSWER/mem[1][5][0] , \ANSWER/mem[1][4][15] ,
         \ANSWER/mem[1][4][14] , \ANSWER/mem[1][4][13] ,
         \ANSWER/mem[1][4][12] , \ANSWER/mem[1][4][11] ,
         \ANSWER/mem[1][4][10] , \ANSWER/mem[1][4][9] , \ANSWER/mem[1][4][8] ,
         \ANSWER/mem[1][4][7] , \ANSWER/mem[1][4][6] , \ANSWER/mem[1][4][5] ,
         \ANSWER/mem[1][4][4] , \ANSWER/mem[1][4][3] , \ANSWER/mem[1][4][2] ,
         \ANSWER/mem[1][4][1] , \ANSWER/mem[1][4][0] , \ANSWER/mem[1][3][15] ,
         \ANSWER/mem[1][3][14] , \ANSWER/mem[1][3][13] ,
         \ANSWER/mem[1][3][12] , \ANSWER/mem[1][3][11] ,
         \ANSWER/mem[1][3][10] , \ANSWER/mem[1][3][9] , \ANSWER/mem[1][3][8] ,
         \ANSWER/mem[1][3][7] , \ANSWER/mem[1][3][6] , \ANSWER/mem[1][3][5] ,
         \ANSWER/mem[1][3][4] , \ANSWER/mem[1][3][3] , \ANSWER/mem[1][3][2] ,
         \ANSWER/mem[1][3][1] , \ANSWER/mem[1][3][0] , \ANSWER/mem[1][2][15] ,
         \ANSWER/mem[1][2][14] , \ANSWER/mem[1][2][13] ,
         \ANSWER/mem[1][2][12] , \ANSWER/mem[1][2][11] ,
         \ANSWER/mem[1][2][10] , \ANSWER/mem[1][2][9] , \ANSWER/mem[1][2][8] ,
         \ANSWER/mem[1][2][7] , \ANSWER/mem[1][2][6] , \ANSWER/mem[1][2][5] ,
         \ANSWER/mem[1][2][4] , \ANSWER/mem[1][2][3] , \ANSWER/mem[1][2][2] ,
         \ANSWER/mem[1][2][1] , \ANSWER/mem[1][2][0] , \ANSWER/mem[1][1][15] ,
         \ANSWER/mem[1][1][14] , \ANSWER/mem[1][1][13] ,
         \ANSWER/mem[1][1][12] , \ANSWER/mem[1][1][11] ,
         \ANSWER/mem[1][1][10] , \ANSWER/mem[1][1][9] , \ANSWER/mem[1][1][8] ,
         \ANSWER/mem[1][1][7] , \ANSWER/mem[1][1][6] , \ANSWER/mem[1][1][5] ,
         \ANSWER/mem[1][1][4] , \ANSWER/mem[1][1][3] , \ANSWER/mem[1][1][2] ,
         \ANSWER/mem[1][1][1] , \ANSWER/mem[1][1][0] , \ANSWER/mem[1][0][15] ,
         \ANSWER/mem[1][0][14] , \ANSWER/mem[1][0][13] ,
         \ANSWER/mem[1][0][12] , \ANSWER/mem[1][0][11] ,
         \ANSWER/mem[1][0][10] , \ANSWER/mem[1][0][9] , \ANSWER/mem[1][0][8] ,
         \ANSWER/mem[1][0][7] , \ANSWER/mem[1][0][6] , \ANSWER/mem[1][0][5] ,
         \ANSWER/mem[1][0][4] , \ANSWER/mem[1][0][3] , \ANSWER/mem[1][0][2] ,
         \ANSWER/mem[1][0][1] , \ANSWER/mem[1][0][0] , \ANSWER/mem[0][9][15] ,
         \ANSWER/mem[0][9][14] , \ANSWER/mem[0][9][13] ,
         \ANSWER/mem[0][9][12] , \ANSWER/mem[0][9][11] ,
         \ANSWER/mem[0][9][10] , \ANSWER/mem[0][9][9] , \ANSWER/mem[0][9][8] ,
         \ANSWER/mem[0][9][7] , \ANSWER/mem[0][9][6] , \ANSWER/mem[0][9][5] ,
         \ANSWER/mem[0][9][4] , \ANSWER/mem[0][9][3] , \ANSWER/mem[0][9][2] ,
         \ANSWER/mem[0][9][1] , \ANSWER/mem[0][9][0] , \ANSWER/mem[0][8][15] ,
         \ANSWER/mem[0][8][14] , \ANSWER/mem[0][8][13] ,
         \ANSWER/mem[0][8][12] , \ANSWER/mem[0][8][11] ,
         \ANSWER/mem[0][8][10] , \ANSWER/mem[0][8][9] , \ANSWER/mem[0][8][8] ,
         \ANSWER/mem[0][8][7] , \ANSWER/mem[0][8][6] , \ANSWER/mem[0][8][5] ,
         \ANSWER/mem[0][8][4] , \ANSWER/mem[0][8][3] , \ANSWER/mem[0][8][2] ,
         \ANSWER/mem[0][8][1] , \ANSWER/mem[0][8][0] , \ANSWER/mem[0][7][15] ,
         \ANSWER/mem[0][7][14] , \ANSWER/mem[0][7][13] ,
         \ANSWER/mem[0][7][12] , \ANSWER/mem[0][7][11] ,
         \ANSWER/mem[0][7][10] , \ANSWER/mem[0][7][9] , \ANSWER/mem[0][7][8] ,
         \ANSWER/mem[0][7][7] , \ANSWER/mem[0][7][6] , \ANSWER/mem[0][7][5] ,
         \ANSWER/mem[0][7][4] , \ANSWER/mem[0][7][3] , \ANSWER/mem[0][7][2] ,
         \ANSWER/mem[0][7][1] , \ANSWER/mem[0][7][0] , \ANSWER/mem[0][6][15] ,
         \ANSWER/mem[0][6][14] , \ANSWER/mem[0][6][13] ,
         \ANSWER/mem[0][6][12] , \ANSWER/mem[0][6][11] ,
         \ANSWER/mem[0][6][10] , \ANSWER/mem[0][6][9] , \ANSWER/mem[0][6][8] ,
         \ANSWER/mem[0][6][7] , \ANSWER/mem[0][6][6] , \ANSWER/mem[0][6][5] ,
         \ANSWER/mem[0][6][4] , \ANSWER/mem[0][6][3] , \ANSWER/mem[0][6][2] ,
         \ANSWER/mem[0][6][1] , \ANSWER/mem[0][6][0] , \ANSWER/mem[0][5][15] ,
         \ANSWER/mem[0][5][14] , \ANSWER/mem[0][5][13] ,
         \ANSWER/mem[0][5][12] , \ANSWER/mem[0][5][11] ,
         \ANSWER/mem[0][5][10] , \ANSWER/mem[0][5][9] , \ANSWER/mem[0][5][8] ,
         \ANSWER/mem[0][5][7] , \ANSWER/mem[0][5][6] , \ANSWER/mem[0][5][5] ,
         \ANSWER/mem[0][5][4] , \ANSWER/mem[0][5][3] , \ANSWER/mem[0][5][2] ,
         \ANSWER/mem[0][5][1] , \ANSWER/mem[0][5][0] , \ANSWER/mem[0][4][15] ,
         \ANSWER/mem[0][4][14] , \ANSWER/mem[0][4][13] ,
         \ANSWER/mem[0][4][12] , \ANSWER/mem[0][4][11] ,
         \ANSWER/mem[0][4][10] , \ANSWER/mem[0][4][9] , \ANSWER/mem[0][4][8] ,
         \ANSWER/mem[0][4][7] , \ANSWER/mem[0][4][6] , \ANSWER/mem[0][4][5] ,
         \ANSWER/mem[0][4][4] , \ANSWER/mem[0][4][3] , \ANSWER/mem[0][4][2] ,
         \ANSWER/mem[0][4][1] , \ANSWER/mem[0][4][0] , \ANSWER/mem[0][3][15] ,
         \ANSWER/mem[0][3][14] , \ANSWER/mem[0][3][13] ,
         \ANSWER/mem[0][3][12] , \ANSWER/mem[0][3][11] ,
         \ANSWER/mem[0][3][10] , \ANSWER/mem[0][3][9] , \ANSWER/mem[0][3][8] ,
         \ANSWER/mem[0][3][7] , \ANSWER/mem[0][3][6] , \ANSWER/mem[0][3][5] ,
         \ANSWER/mem[0][3][4] , \ANSWER/mem[0][3][3] , \ANSWER/mem[0][3][2] ,
         \ANSWER/mem[0][3][1] , \ANSWER/mem[0][3][0] , \ANSWER/mem[0][2][15] ,
         \ANSWER/mem[0][2][14] , \ANSWER/mem[0][2][13] ,
         \ANSWER/mem[0][2][12] , \ANSWER/mem[0][2][11] ,
         \ANSWER/mem[0][2][10] , \ANSWER/mem[0][2][9] , \ANSWER/mem[0][2][8] ,
         \ANSWER/mem[0][2][7] , \ANSWER/mem[0][2][6] , \ANSWER/mem[0][2][5] ,
         \ANSWER/mem[0][2][4] , \ANSWER/mem[0][2][3] , \ANSWER/mem[0][2][2] ,
         \ANSWER/mem[0][2][1] , \ANSWER/mem[0][2][0] , \ANSWER/mem[0][1][15] ,
         \ANSWER/mem[0][1][14] , \ANSWER/mem[0][1][13] ,
         \ANSWER/mem[0][1][12] , \ANSWER/mem[0][1][11] ,
         \ANSWER/mem[0][1][10] , \ANSWER/mem[0][1][9] , \ANSWER/mem[0][1][8] ,
         \ANSWER/mem[0][1][7] , \ANSWER/mem[0][1][6] , \ANSWER/mem[0][1][5] ,
         \ANSWER/mem[0][1][4] , \ANSWER/mem[0][1][3] , \ANSWER/mem[0][1][2] ,
         \ANSWER/mem[0][1][1] , \ANSWER/mem[0][1][0] , \ANSWER/mem[0][0][15] ,
         \ANSWER/mem[0][0][14] , \ANSWER/mem[0][0][13] ,
         \ANSWER/mem[0][0][12] , \ANSWER/mem[0][0][11] ,
         \ANSWER/mem[0][0][10] , \ANSWER/mem[0][0][9] , \ANSWER/mem[0][0][8] ,
         \ANSWER/mem[0][0][7] , \ANSWER/mem[0][0][6] , \ANSWER/mem[0][0][5] ,
         \ANSWER/mem[0][0][4] , \ANSWER/mem[0][0][3] , \ANSWER/mem[0][0][2] ,
         \ANSWER/mem[0][0][1] , \ANSWER/mem[0][0][0] , \SIGMOID/N64 ,
         \SIGMOID/sign_bit , n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4111, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
         n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
         n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822,
         n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
         n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918,
         n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
         n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
         n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966,
         n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
         n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982,
         n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990,
         n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
         n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
         n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014,
         n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
         n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030,
         n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038,
         n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
         n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054,
         n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062,
         n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070,
         n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078,
         n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086,
         n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
         n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102,
         n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110,
         n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
         n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126,
         n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134,
         n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142,
         n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150,
         n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158,
         n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
         n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
         n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182,
         n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
         n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206,
         n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214,
         n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222,
         n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230,
         n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
         n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
         n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254,
         n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
         n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270,
         n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
         n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
         n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
         n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
         n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
         n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
         n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
         n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
         n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
         n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
         n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
         n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558,
         n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566,
         n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
         n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
         n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
         n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614,
         n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
         n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630,
         n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
         n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
         n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654,
         n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662,
         n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670,
         n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
         n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686,
         n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
         n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702,
         n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710,
         n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
         n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726,
         n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
         n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
         n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
         n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
         n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
         n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
         n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
         n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814,
         n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
         n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
         n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
         n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
         n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
         n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
         n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
         n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
         n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
         n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950,
         n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
         n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998,
         n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006,
         n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
         n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022,
         n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030,
         n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
         n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
         n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
         n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
         n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070,
         n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078,
         n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086,
         n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094,
         n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
         n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110,
         n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118,
         n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
         n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
         n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142,
         n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150,
         n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
         n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166,
         n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
         n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
         n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190,
         n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
         n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
         n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214,
         n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
         n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230,
         n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238,
         n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
         n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
         n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262,
         n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
         n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278,
         n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
         n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
         n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
         n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
         n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
         n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
         n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
         n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
         n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
         n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
         n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
         n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
         n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
         n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366,
         n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
         n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
         n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
         n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
         n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
         n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
         n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
         n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
         n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
         n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
         n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
         n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
         n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
         n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
         n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
         n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
         n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
         n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
         n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
         n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
         n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686,
         n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
         n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702,
         n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
         n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
         n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
         n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734,
         n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
         n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
         n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758,
         n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
         n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774,
         n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
         n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
         n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798,
         n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
         n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
         n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
         n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830,
         n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
         n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
         n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
         n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
         n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
         n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
         n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
         n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918;
  wire   [159:0] m1Inputs;
  wire   [159:0] column;
  wire   [15:0] m2DataIn;
  wire   [15:0] q_w2;
  wire   [15:0] \STAGE_1/weightReg ;
  wire   [15:0] \STAGE_1/M1/sum ;
  wire   [15:0] \STAGE_1/M2/sum ;
  wire   [15:0] \STAGE_1/M3/sum ;
  wire   [15:0] \STAGE_1/M4/sum ;
  wire   [15:0] \STAGE_1/M5/sum ;
  wire   [15:0] \STAGE_1/M6/sum ;
  wire   [15:0] \STAGE_1/M7/sum ;
  wire   [15:0] \STAGE_1/M8/sum ;
  wire   [15:0] \STAGE_1/M9/sum ;
  wire   [15:0] \STAGE_1/M10/sum ;
  wire   [4:0] \CNTRL/count_20Q ;
  wire   [3:0] \CNTRL/count_10_2Q ;
  wire   [3:0] \CNTRL/count_10Q ;
  wire   [7:0] \CNTRL/count_layer1_200Q ;
  wire   [9:0] \CNTRL/count_layer1_784Q ;
  wire   [3:0] \CNTRL/currentState ;
  wire   [159:0] \ROUTEDATA/regData ;
  wire   [15:0] \SIGMOID/lut_out ;

  dp_1 \STAGE_1/weightReg_reg[0]  ( .ip(weight1[0]), .ck(clk), .q(
        \STAGE_1/weightReg [0]) );
  dp_1 \STAGE_1/weightReg_reg[1]  ( .ip(weight1[1]), .ck(clk), .q(
        \STAGE_1/weightReg [1]) );
  dp_1 \STAGE_1/weightReg_reg[2]  ( .ip(weight1[2]), .ck(clk), .q(
        \STAGE_1/weightReg [2]) );
  dp_1 \STAGE_1/weightReg_reg[4]  ( .ip(weight1[4]), .ck(clk), .q(
        \STAGE_1/weightReg [4]) );
  dp_1 \STAGE_1/weightReg_reg[5]  ( .ip(weight1[5]), .ck(clk), .q(
        \STAGE_1/weightReg [5]) );
  dp_1 \STAGE_1/weightReg_reg[8]  ( .ip(weight1[8]), .ck(clk), .q(
        \STAGE_1/weightReg [8]) );
  dp_1 \STAGE_1/weightReg_reg[9]  ( .ip(weight1[9]), .ck(clk), .q(
        \STAGE_1/weightReg [9]) );
  dp_1 \STAGE_1/weightReg_reg[10]  ( .ip(weight1[10]), .ck(clk), .q(
        \STAGE_1/weightReg [10]) );
  dp_1 \STAGE_1/weightReg_reg[11]  ( .ip(weight1[11]), .ck(clk), .q(
        \STAGE_1/weightReg [11]) );
  dp_1 \STAGE_1/weightReg_reg[12]  ( .ip(weight1[12]), .ck(clk), .q(
        \STAGE_1/weightReg [12]) );
  dp_1 \STAGE_1/weightReg_reg[13]  ( .ip(weight1[13]), .ck(clk), .q(
        \STAGE_1/weightReg [13]) );
  dp_1 \STAGE_1/weightReg_reg[14]  ( .ip(weight1[14]), .ck(clk), .q(
        \STAGE_1/weightReg [14]) );
  dp_1 \STAGE_1/M1/result_reg[0]  ( .ip(\STAGE_1/M1/sum [0]), .ck(clk), .q(
        column[0]) );
  dp_1 \STAGE_1/M1/result_reg[1]  ( .ip(\STAGE_1/M1/sum [1]), .ck(clk), .q(
        column[1]) );
  dp_1 \STAGE_1/M1/result_reg[2]  ( .ip(\STAGE_1/M1/sum [2]), .ck(clk), .q(
        column[2]) );
  dp_1 \STAGE_1/M1/result_reg[3]  ( .ip(\STAGE_1/M1/sum [3]), .ck(clk), .q(
        column[3]) );
  dp_1 \STAGE_1/M1/result_reg[4]  ( .ip(\STAGE_1/M1/sum [4]), .ck(clk), .q(
        column[4]) );
  dp_1 \STAGE_1/M1/result_reg[5]  ( .ip(\STAGE_1/M1/sum [5]), .ck(clk), .q(
        column[5]) );
  dp_1 \STAGE_1/M1/result_reg[6]  ( .ip(\STAGE_1/M1/sum [6]), .ck(clk), .q(
        column[6]) );
  dp_1 \STAGE_1/M1/result_reg[7]  ( .ip(\STAGE_1/M1/sum [7]), .ck(clk), .q(
        column[7]) );
  dp_1 \STAGE_1/M1/result_reg[8]  ( .ip(\STAGE_1/M1/sum [8]), .ck(clk), .q(
        column[8]) );
  dp_1 \STAGE_1/M1/result_reg[9]  ( .ip(\STAGE_1/M1/sum [9]), .ck(clk), .q(
        column[9]) );
  dp_1 \STAGE_1/M1/result_reg[10]  ( .ip(\STAGE_1/M1/sum [10]), .ck(clk), .q(
        column[10]) );
  dp_1 \STAGE_1/M1/result_reg[11]  ( .ip(\STAGE_1/M1/sum [11]), .ck(clk), .q(
        column[11]) );
  dp_1 \STAGE_1/M1/result_reg[12]  ( .ip(\STAGE_1/M1/sum [12]), .ck(clk), .q(
        column[12]) );
  dp_1 \STAGE_1/M1/result_reg[13]  ( .ip(\STAGE_1/M1/sum [13]), .ck(clk), .q(
        column[13]) );
  dp_1 \STAGE_1/M1/result_reg[14]  ( .ip(\STAGE_1/M1/sum [14]), .ck(clk), .q(
        column[14]) );
  dp_1 \STAGE_1/M1/result_reg[15]  ( .ip(\STAGE_1/M1/sum [15]), .ck(clk), .q(
        column[15]) );
  dp_1 \STAGE_1/M2/result_reg[0]  ( .ip(\STAGE_1/M2/sum [0]), .ck(clk), .q(
        column[16]) );
  dp_1 \STAGE_1/M2/result_reg[1]  ( .ip(\STAGE_1/M2/sum [1]), .ck(clk), .q(
        column[17]) );
  dp_1 \STAGE_1/M2/result_reg[2]  ( .ip(\STAGE_1/M2/sum [2]), .ck(clk), .q(
        column[18]) );
  dp_1 \STAGE_1/M2/result_reg[3]  ( .ip(\STAGE_1/M2/sum [3]), .ck(clk), .q(
        column[19]) );
  dp_1 \STAGE_1/M2/result_reg[4]  ( .ip(\STAGE_1/M2/sum [4]), .ck(clk), .q(
        column[20]) );
  dp_1 \STAGE_1/M2/result_reg[5]  ( .ip(\STAGE_1/M2/sum [5]), .ck(clk), .q(
        column[21]) );
  dp_1 \STAGE_1/M2/result_reg[6]  ( .ip(\STAGE_1/M2/sum [6]), .ck(clk), .q(
        column[22]) );
  dp_1 \STAGE_1/M2/result_reg[7]  ( .ip(\STAGE_1/M2/sum [7]), .ck(clk), .q(
        column[23]) );
  dp_1 \STAGE_1/M2/result_reg[8]  ( .ip(\STAGE_1/M2/sum [8]), .ck(clk), .q(
        column[24]) );
  dp_1 \STAGE_1/M2/result_reg[9]  ( .ip(\STAGE_1/M2/sum [9]), .ck(clk), .q(
        column[25]) );
  dp_1 \STAGE_1/M2/result_reg[10]  ( .ip(\STAGE_1/M2/sum [10]), .ck(clk), .q(
        column[26]) );
  dp_1 \STAGE_1/M2/result_reg[11]  ( .ip(\STAGE_1/M2/sum [11]), .ck(clk), .q(
        column[27]) );
  dp_1 \STAGE_1/M2/result_reg[12]  ( .ip(\STAGE_1/M2/sum [12]), .ck(clk), .q(
        column[28]) );
  dp_1 \STAGE_1/M2/result_reg[13]  ( .ip(\STAGE_1/M2/sum [13]), .ck(clk), .q(
        column[29]) );
  dp_1 \STAGE_1/M2/result_reg[14]  ( .ip(\STAGE_1/M2/sum [14]), .ck(clk), .q(
        column[30]) );
  dp_1 \STAGE_1/M2/result_reg[15]  ( .ip(\STAGE_1/M2/sum [15]), .ck(clk), .q(
        column[31]) );
  dp_1 \STAGE_1/M3/result_reg[0]  ( .ip(\STAGE_1/M3/sum [0]), .ck(clk), .q(
        column[32]) );
  dp_1 \STAGE_1/M3/result_reg[1]  ( .ip(\STAGE_1/M3/sum [1]), .ck(clk), .q(
        column[33]) );
  dp_1 \STAGE_1/M3/result_reg[2]  ( .ip(\STAGE_1/M3/sum [2]), .ck(clk), .q(
        column[34]) );
  dp_1 \STAGE_1/M3/result_reg[3]  ( .ip(\STAGE_1/M3/sum [3]), .ck(clk), .q(
        column[35]) );
  dp_1 \STAGE_1/M3/result_reg[4]  ( .ip(\STAGE_1/M3/sum [4]), .ck(clk), .q(
        column[36]) );
  dp_1 \STAGE_1/M3/result_reg[5]  ( .ip(\STAGE_1/M3/sum [5]), .ck(clk), .q(
        column[37]) );
  dp_1 \STAGE_1/M3/result_reg[6]  ( .ip(\STAGE_1/M3/sum [6]), .ck(clk), .q(
        column[38]) );
  dp_1 \STAGE_1/M3/result_reg[7]  ( .ip(\STAGE_1/M3/sum [7]), .ck(clk), .q(
        column[39]) );
  dp_1 \STAGE_1/M3/result_reg[8]  ( .ip(\STAGE_1/M3/sum [8]), .ck(clk), .q(
        column[40]) );
  dp_1 \STAGE_1/M3/result_reg[9]  ( .ip(\STAGE_1/M3/sum [9]), .ck(clk), .q(
        column[41]) );
  dp_1 \STAGE_1/M3/result_reg[10]  ( .ip(\STAGE_1/M3/sum [10]), .ck(clk), .q(
        column[42]) );
  dp_1 \STAGE_1/M3/result_reg[11]  ( .ip(\STAGE_1/M3/sum [11]), .ck(clk), .q(
        column[43]) );
  dp_1 \STAGE_1/M3/result_reg[12]  ( .ip(\STAGE_1/M3/sum [12]), .ck(clk), .q(
        column[44]) );
  dp_1 \STAGE_1/M3/result_reg[13]  ( .ip(\STAGE_1/M3/sum [13]), .ck(clk), .q(
        column[45]) );
  dp_1 \STAGE_1/M3/result_reg[14]  ( .ip(\STAGE_1/M3/sum [14]), .ck(clk), .q(
        column[46]) );
  dp_1 \STAGE_1/M3/result_reg[15]  ( .ip(\STAGE_1/M3/sum [15]), .ck(clk), .q(
        column[47]) );
  dp_1 \STAGE_1/M4/result_reg[0]  ( .ip(\STAGE_1/M4/sum [0]), .ck(clk), .q(
        column[48]) );
  dp_1 \STAGE_1/M4/result_reg[1]  ( .ip(\STAGE_1/M4/sum [1]), .ck(clk), .q(
        column[49]) );
  dp_1 \STAGE_1/M4/result_reg[2]  ( .ip(\STAGE_1/M4/sum [2]), .ck(clk), .q(
        column[50]) );
  dp_1 \STAGE_1/M4/result_reg[3]  ( .ip(\STAGE_1/M4/sum [3]), .ck(clk), .q(
        column[51]) );
  dp_1 \STAGE_1/M4/result_reg[4]  ( .ip(\STAGE_1/M4/sum [4]), .ck(clk), .q(
        column[52]) );
  dp_1 \STAGE_1/M4/result_reg[5]  ( .ip(\STAGE_1/M4/sum [5]), .ck(clk), .q(
        column[53]) );
  dp_1 \STAGE_1/M4/result_reg[6]  ( .ip(\STAGE_1/M4/sum [6]), .ck(clk), .q(
        column[54]) );
  dp_1 \STAGE_1/M4/result_reg[7]  ( .ip(\STAGE_1/M4/sum [7]), .ck(clk), .q(
        column[55]) );
  dp_1 \STAGE_1/M4/result_reg[8]  ( .ip(\STAGE_1/M4/sum [8]), .ck(clk), .q(
        column[56]) );
  dp_1 \STAGE_1/M4/result_reg[9]  ( .ip(\STAGE_1/M4/sum [9]), .ck(clk), .q(
        column[57]) );
  dp_1 \STAGE_1/M4/result_reg[10]  ( .ip(\STAGE_1/M4/sum [10]), .ck(clk), .q(
        column[58]) );
  dp_1 \STAGE_1/M4/result_reg[11]  ( .ip(\STAGE_1/M4/sum [11]), .ck(clk), .q(
        column[59]) );
  dp_1 \STAGE_1/M4/result_reg[12]  ( .ip(\STAGE_1/M4/sum [12]), .ck(clk), .q(
        column[60]) );
  dp_1 \STAGE_1/M4/result_reg[13]  ( .ip(\STAGE_1/M4/sum [13]), .ck(clk), .q(
        column[61]) );
  dp_1 \STAGE_1/M4/result_reg[14]  ( .ip(\STAGE_1/M4/sum [14]), .ck(clk), .q(
        column[62]) );
  dp_1 \STAGE_1/M4/result_reg[15]  ( .ip(\STAGE_1/M4/sum [15]), .ck(clk), .q(
        column[63]) );
  dp_1 \STAGE_1/M5/result_reg[0]  ( .ip(\STAGE_1/M5/sum [0]), .ck(clk), .q(
        column[64]) );
  dp_1 \STAGE_1/M5/result_reg[1]  ( .ip(\STAGE_1/M5/sum [1]), .ck(clk), .q(
        column[65]) );
  dp_1 \STAGE_1/M5/result_reg[2]  ( .ip(\STAGE_1/M5/sum [2]), .ck(clk), .q(
        column[66]) );
  dp_1 \STAGE_1/M5/result_reg[3]  ( .ip(\STAGE_1/M5/sum [3]), .ck(clk), .q(
        column[67]) );
  dp_1 \STAGE_1/M5/result_reg[4]  ( .ip(\STAGE_1/M5/sum [4]), .ck(clk), .q(
        column[68]) );
  dp_1 \STAGE_1/M5/result_reg[5]  ( .ip(\STAGE_1/M5/sum [5]), .ck(clk), .q(
        column[69]) );
  dp_1 \STAGE_1/M5/result_reg[6]  ( .ip(\STAGE_1/M5/sum [6]), .ck(clk), .q(
        column[70]) );
  dp_1 \STAGE_1/M5/result_reg[7]  ( .ip(\STAGE_1/M5/sum [7]), .ck(clk), .q(
        column[71]) );
  dp_1 \STAGE_1/M5/result_reg[8]  ( .ip(\STAGE_1/M5/sum [8]), .ck(clk), .q(
        column[72]) );
  dp_1 \STAGE_1/M5/result_reg[9]  ( .ip(\STAGE_1/M5/sum [9]), .ck(clk), .q(
        column[73]) );
  dp_1 \STAGE_1/M5/result_reg[10]  ( .ip(\STAGE_1/M5/sum [10]), .ck(clk), .q(
        column[74]) );
  dp_1 \STAGE_1/M5/result_reg[11]  ( .ip(\STAGE_1/M5/sum [11]), .ck(clk), .q(
        column[75]) );
  dp_1 \STAGE_1/M5/result_reg[12]  ( .ip(\STAGE_1/M5/sum [12]), .ck(clk), .q(
        column[76]) );
  dp_1 \STAGE_1/M5/result_reg[13]  ( .ip(\STAGE_1/M5/sum [13]), .ck(clk), .q(
        column[77]) );
  dp_1 \STAGE_1/M5/result_reg[14]  ( .ip(\STAGE_1/M5/sum [14]), .ck(clk), .q(
        column[78]) );
  dp_1 \STAGE_1/M5/result_reg[15]  ( .ip(\STAGE_1/M5/sum [15]), .ck(clk), .q(
        column[79]) );
  dp_1 \STAGE_1/M6/result_reg[0]  ( .ip(\STAGE_1/M6/sum [0]), .ck(clk), .q(
        column[80]) );
  dp_1 \STAGE_1/M6/result_reg[1]  ( .ip(\STAGE_1/M6/sum [1]), .ck(clk), .q(
        column[81]) );
  dp_1 \STAGE_1/M6/result_reg[2]  ( .ip(\STAGE_1/M6/sum [2]), .ck(clk), .q(
        column[82]) );
  dp_1 \STAGE_1/M6/result_reg[3]  ( .ip(\STAGE_1/M6/sum [3]), .ck(clk), .q(
        column[83]) );
  dp_1 \STAGE_1/M6/result_reg[4]  ( .ip(\STAGE_1/M6/sum [4]), .ck(clk), .q(
        column[84]) );
  dp_1 \STAGE_1/M6/result_reg[5]  ( .ip(\STAGE_1/M6/sum [5]), .ck(clk), .q(
        column[85]) );
  dp_1 \STAGE_1/M6/result_reg[6]  ( .ip(\STAGE_1/M6/sum [6]), .ck(clk), .q(
        column[86]) );
  dp_1 \STAGE_1/M6/result_reg[7]  ( .ip(\STAGE_1/M6/sum [7]), .ck(clk), .q(
        column[87]) );
  dp_1 \STAGE_1/M6/result_reg[8]  ( .ip(\STAGE_1/M6/sum [8]), .ck(clk), .q(
        column[88]) );
  dp_1 \STAGE_1/M6/result_reg[9]  ( .ip(\STAGE_1/M6/sum [9]), .ck(clk), .q(
        column[89]) );
  dp_1 \STAGE_1/M6/result_reg[10]  ( .ip(\STAGE_1/M6/sum [10]), .ck(clk), .q(
        column[90]) );
  dp_1 \STAGE_1/M6/result_reg[11]  ( .ip(\STAGE_1/M6/sum [11]), .ck(clk), .q(
        column[91]) );
  dp_1 \STAGE_1/M6/result_reg[12]  ( .ip(\STAGE_1/M6/sum [12]), .ck(clk), .q(
        column[92]) );
  dp_1 \STAGE_1/M6/result_reg[13]  ( .ip(\STAGE_1/M6/sum [13]), .ck(clk), .q(
        column[93]) );
  dp_1 \STAGE_1/M6/result_reg[14]  ( .ip(\STAGE_1/M6/sum [14]), .ck(clk), .q(
        column[94]) );
  dp_1 \STAGE_1/M6/result_reg[15]  ( .ip(\STAGE_1/M6/sum [15]), .ck(clk), .q(
        column[95]) );
  dp_1 \STAGE_1/M7/result_reg[0]  ( .ip(\STAGE_1/M7/sum [0]), .ck(clk), .q(
        column[96]) );
  dp_1 \STAGE_1/M7/result_reg[1]  ( .ip(\STAGE_1/M7/sum [1]), .ck(clk), .q(
        column[97]) );
  dp_1 \STAGE_1/M7/result_reg[2]  ( .ip(\STAGE_1/M7/sum [2]), .ck(clk), .q(
        column[98]) );
  dp_1 \STAGE_1/M7/result_reg[3]  ( .ip(\STAGE_1/M7/sum [3]), .ck(clk), .q(
        column[99]) );
  dp_1 \STAGE_1/M7/result_reg[4]  ( .ip(\STAGE_1/M7/sum [4]), .ck(clk), .q(
        column[100]) );
  dp_1 \STAGE_1/M7/result_reg[5]  ( .ip(\STAGE_1/M7/sum [5]), .ck(clk), .q(
        column[101]) );
  dp_1 \STAGE_1/M7/result_reg[6]  ( .ip(\STAGE_1/M7/sum [6]), .ck(clk), .q(
        column[102]) );
  dp_1 \STAGE_1/M7/result_reg[7]  ( .ip(\STAGE_1/M7/sum [7]), .ck(clk), .q(
        column[103]) );
  dp_1 \STAGE_1/M7/result_reg[8]  ( .ip(\STAGE_1/M7/sum [8]), .ck(clk), .q(
        column[104]) );
  dp_1 \STAGE_1/M7/result_reg[9]  ( .ip(\STAGE_1/M7/sum [9]), .ck(clk), .q(
        column[105]) );
  dp_1 \STAGE_1/M7/result_reg[10]  ( .ip(\STAGE_1/M7/sum [10]), .ck(clk), .q(
        column[106]) );
  dp_1 \STAGE_1/M7/result_reg[11]  ( .ip(\STAGE_1/M7/sum [11]), .ck(clk), .q(
        column[107]) );
  dp_1 \STAGE_1/M7/result_reg[12]  ( .ip(\STAGE_1/M7/sum [12]), .ck(clk), .q(
        column[108]) );
  dp_1 \STAGE_1/M7/result_reg[13]  ( .ip(\STAGE_1/M7/sum [13]), .ck(clk), .q(
        column[109]) );
  dp_1 \STAGE_1/M7/result_reg[14]  ( .ip(\STAGE_1/M7/sum [14]), .ck(clk), .q(
        column[110]) );
  dp_1 \STAGE_1/M7/result_reg[15]  ( .ip(\STAGE_1/M7/sum [15]), .ck(clk), .q(
        column[111]) );
  dp_1 \STAGE_1/M8/result_reg[0]  ( .ip(\STAGE_1/M8/sum [0]), .ck(clk), .q(
        column[112]) );
  dp_1 \STAGE_1/M8/result_reg[1]  ( .ip(\STAGE_1/M8/sum [1]), .ck(clk), .q(
        column[113]) );
  dp_1 \STAGE_1/M8/result_reg[2]  ( .ip(\STAGE_1/M8/sum [2]), .ck(clk), .q(
        column[114]) );
  dp_1 \STAGE_1/M8/result_reg[3]  ( .ip(\STAGE_1/M8/sum [3]), .ck(clk), .q(
        column[115]) );
  dp_1 \STAGE_1/M8/result_reg[4]  ( .ip(\STAGE_1/M8/sum [4]), .ck(clk), .q(
        column[116]) );
  dp_1 \STAGE_1/M8/result_reg[5]  ( .ip(\STAGE_1/M8/sum [5]), .ck(clk), .q(
        column[117]) );
  dp_1 \STAGE_1/M8/result_reg[6]  ( .ip(\STAGE_1/M8/sum [6]), .ck(clk), .q(
        column[118]) );
  dp_1 \STAGE_1/M8/result_reg[7]  ( .ip(\STAGE_1/M8/sum [7]), .ck(clk), .q(
        column[119]) );
  dp_1 \STAGE_1/M8/result_reg[8]  ( .ip(\STAGE_1/M8/sum [8]), .ck(clk), .q(
        column[120]) );
  dp_1 \STAGE_1/M8/result_reg[9]  ( .ip(\STAGE_1/M8/sum [9]), .ck(clk), .q(
        column[121]) );
  dp_1 \STAGE_1/M8/result_reg[10]  ( .ip(\STAGE_1/M8/sum [10]), .ck(clk), .q(
        column[122]) );
  dp_1 \STAGE_1/M8/result_reg[11]  ( .ip(\STAGE_1/M8/sum [11]), .ck(clk), .q(
        column[123]) );
  dp_1 \STAGE_1/M8/result_reg[12]  ( .ip(\STAGE_1/M8/sum [12]), .ck(clk), .q(
        column[124]) );
  dp_1 \STAGE_1/M8/result_reg[13]  ( .ip(\STAGE_1/M8/sum [13]), .ck(clk), .q(
        column[125]) );
  dp_1 \STAGE_1/M8/result_reg[14]  ( .ip(\STAGE_1/M8/sum [14]), .ck(clk), .q(
        column[126]) );
  dp_1 \STAGE_1/M8/result_reg[15]  ( .ip(\STAGE_1/M8/sum [15]), .ck(clk), .q(
        column[127]) );
  dp_1 \STAGE_1/M9/result_reg[0]  ( .ip(\STAGE_1/M9/sum [0]), .ck(clk), .q(
        column[128]) );
  dp_1 \STAGE_1/M9/result_reg[1]  ( .ip(\STAGE_1/M9/sum [1]), .ck(clk), .q(
        column[129]) );
  dp_1 \STAGE_1/M9/result_reg[2]  ( .ip(\STAGE_1/M9/sum [2]), .ck(clk), .q(
        column[130]) );
  dp_1 \STAGE_1/M9/result_reg[3]  ( .ip(\STAGE_1/M9/sum [3]), .ck(clk), .q(
        column[131]) );
  dp_1 \STAGE_1/M9/result_reg[4]  ( .ip(\STAGE_1/M9/sum [4]), .ck(clk), .q(
        column[132]) );
  dp_1 \STAGE_1/M9/result_reg[5]  ( .ip(\STAGE_1/M9/sum [5]), .ck(clk), .q(
        column[133]) );
  dp_1 \STAGE_1/M9/result_reg[6]  ( .ip(\STAGE_1/M9/sum [6]), .ck(clk), .q(
        column[134]) );
  dp_1 \STAGE_1/M9/result_reg[7]  ( .ip(\STAGE_1/M9/sum [7]), .ck(clk), .q(
        column[135]) );
  dp_1 \STAGE_1/M9/result_reg[8]  ( .ip(\STAGE_1/M9/sum [8]), .ck(clk), .q(
        column[136]) );
  dp_1 \STAGE_1/M9/result_reg[9]  ( .ip(\STAGE_1/M9/sum [9]), .ck(clk), .q(
        column[137]) );
  dp_1 \STAGE_1/M9/result_reg[10]  ( .ip(\STAGE_1/M9/sum [10]), .ck(clk), .q(
        column[138]) );
  dp_1 \STAGE_1/M9/result_reg[11]  ( .ip(\STAGE_1/M9/sum [11]), .ck(clk), .q(
        column[139]) );
  dp_1 \STAGE_1/M9/result_reg[12]  ( .ip(\STAGE_1/M9/sum [12]), .ck(clk), .q(
        column[140]) );
  dp_1 \STAGE_1/M9/result_reg[13]  ( .ip(\STAGE_1/M9/sum [13]), .ck(clk), .q(
        column[141]) );
  dp_1 \STAGE_1/M9/result_reg[14]  ( .ip(\STAGE_1/M9/sum [14]), .ck(clk), .q(
        column[142]) );
  dp_1 \STAGE_1/M9/result_reg[15]  ( .ip(\STAGE_1/M9/sum [15]), .ck(clk), .q(
        column[143]) );
  dp_1 \STAGE_1/M10/result_reg[0]  ( .ip(\STAGE_1/M10/sum [0]), .ck(clk), .q(
        column[144]) );
  dp_1 \STAGE_1/M10/result_reg[1]  ( .ip(\STAGE_1/M10/sum [1]), .ck(clk), .q(
        column[145]) );
  dp_1 \STAGE_1/M10/result_reg[2]  ( .ip(\STAGE_1/M10/sum [2]), .ck(clk), .q(
        column[146]) );
  dp_1 \STAGE_1/M10/result_reg[3]  ( .ip(\STAGE_1/M10/sum [3]), .ck(clk), .q(
        column[147]) );
  dp_1 \STAGE_1/M10/result_reg[4]  ( .ip(\STAGE_1/M10/sum [4]), .ck(clk), .q(
        column[148]) );
  dp_1 \STAGE_1/M10/result_reg[5]  ( .ip(\STAGE_1/M10/sum [5]), .ck(clk), .q(
        column[149]) );
  dp_1 \STAGE_1/M10/result_reg[6]  ( .ip(\STAGE_1/M10/sum [6]), .ck(clk), .q(
        column[150]) );
  dp_1 \STAGE_1/M10/result_reg[7]  ( .ip(\STAGE_1/M10/sum [7]), .ck(clk), .q(
        column[151]) );
  dp_1 \STAGE_1/M10/result_reg[8]  ( .ip(\STAGE_1/M10/sum [8]), .ck(clk), .q(
        column[152]) );
  dp_1 \STAGE_1/M10/result_reg[9]  ( .ip(\STAGE_1/M10/sum [9]), .ck(clk), .q(
        column[153]) );
  dp_1 \STAGE_1/M10/result_reg[10]  ( .ip(\STAGE_1/M10/sum [10]), .ck(clk), 
        .q(column[154]) );
  dp_1 \STAGE_1/M10/result_reg[11]  ( .ip(\STAGE_1/M10/sum [11]), .ck(clk), 
        .q(column[155]) );
  dp_1 \STAGE_1/M10/result_reg[12]  ( .ip(\STAGE_1/M10/sum [12]), .ck(clk), 
        .q(column[156]) );
  dp_1 \STAGE_1/M10/result_reg[13]  ( .ip(\STAGE_1/M10/sum [13]), .ck(clk), 
        .q(column[157]) );
  dp_1 \STAGE_1/M10/result_reg[14]  ( .ip(\STAGE_1/M10/sum [14]), .ck(clk), 
        .q(column[158]) );
  dp_1 \STAGE_1/M10/result_reg[15]  ( .ip(\STAGE_1/M10/sum [15]), .ck(clk), 
        .q(column[159]) );
  dp_1 \INPUTSRAM/q_reg[0]  ( .ip(\INPUTSRAM/mem_i[0][0] ), .ck(clk), .q(
        m1Inputs[0]) );
  dp_1 \INPUTSRAM/q_reg[1]  ( .ip(\INPUTSRAM/mem_i[0][1] ), .ck(clk), .q(
        m1Inputs[1]) );
  dp_1 \INPUTSRAM/q_reg[14]  ( .ip(\INPUTSRAM/mem_i[0][14] ), .ck(clk), .q(
        m1Inputs[14]) );
  dp_1 \INPUTSRAM/q_reg[16]  ( .ip(\INPUTSRAM/mem_i[1][0] ), .ck(clk), .q(
        m1Inputs[16]) );
  dp_1 \INPUTSRAM/q_reg[17]  ( .ip(\INPUTSRAM/mem_i[1][1] ), .ck(clk), .q(
        m1Inputs[17]) );
  dp_1 \INPUTSRAM/q_reg[29]  ( .ip(\INPUTSRAM/mem_i[1][13] ), .ck(clk), .q(
        m1Inputs[29]) );
  dp_1 \INPUTSRAM/q_reg[30]  ( .ip(\INPUTSRAM/mem_i[1][14] ), .ck(clk), .q(
        m1Inputs[30]) );
  dp_1 \INPUTSRAM/q_reg[31]  ( .ip(\INPUTSRAM/mem_i[1][15] ), .ck(clk), .q(
        m1Inputs[31]) );
  dp_1 \INPUTSRAM/q_reg[32]  ( .ip(\INPUTSRAM/mem_i[2][0] ), .ck(clk), .q(
        m1Inputs[32]) );
  dp_1 \INPUTSRAM/q_reg[33]  ( .ip(\INPUTSRAM/mem_i[2][1] ), .ck(clk), .q(
        m1Inputs[33]) );
  dp_1 \INPUTSRAM/q_reg[48]  ( .ip(\INPUTSRAM/mem_i[3][0] ), .ck(clk), .q(
        m1Inputs[48]) );
  dp_1 \INPUTSRAM/q_reg[49]  ( .ip(\INPUTSRAM/mem_i[3][1] ), .ck(clk), .q(
        m1Inputs[49]) );
  dp_1 \INPUTSRAM/q_reg[63]  ( .ip(\INPUTSRAM/mem_i[3][15] ), .ck(clk), .q(
        m1Inputs[63]) );
  dp_1 \INPUTSRAM/q_reg[65]  ( .ip(\INPUTSRAM/mem_i[4][1] ), .ck(clk), .q(
        m1Inputs[65]) );
  dp_1 \INPUTSRAM/q_reg[78]  ( .ip(\INPUTSRAM/mem_i[4][14] ), .ck(clk), .q(
        m1Inputs[78]) );
  dp_1 \INPUTSRAM/q_reg[79]  ( .ip(\INPUTSRAM/mem_i[4][15] ), .ck(clk), .q(
        m1Inputs[79]) );
  dp_1 \INPUTSRAM/q_reg[81]  ( .ip(\INPUTSRAM/mem_i[5][1] ), .ck(clk), .q(
        m1Inputs[81]) );
  dp_1 \INPUTSRAM/q_reg[94]  ( .ip(\INPUTSRAM/mem_i[5][14] ), .ck(clk), .q(
        m1Inputs[94]) );
  dp_1 \INPUTSRAM/q_reg[95]  ( .ip(\INPUTSRAM/mem_i[5][15] ), .ck(clk), .q(
        m1Inputs[95]) );
  dp_1 \INPUTSRAM/q_reg[97]  ( .ip(\INPUTSRAM/mem_i[6][1] ), .ck(clk), .q(
        m1Inputs[97]) );
  dp_1 \INPUTSRAM/q_reg[109]  ( .ip(\INPUTSRAM/mem_i[6][13] ), .ck(clk), .q(
        m1Inputs[109]) );
  dp_1 \INPUTSRAM/q_reg[110]  ( .ip(\INPUTSRAM/mem_i[6][14] ), .ck(clk), .q(
        m1Inputs[110]) );
  dp_1 \INPUTSRAM/q_reg[111]  ( .ip(\INPUTSRAM/mem_i[6][15] ), .ck(clk), .q(
        m1Inputs[111]) );
  dp_1 \INPUTSRAM/q_reg[113]  ( .ip(\INPUTSRAM/mem_i[7][1] ), .ck(clk), .q(
        m1Inputs[113]) );
  dp_1 \INPUTSRAM/q_reg[125]  ( .ip(\INPUTSRAM/mem_i[7][13] ), .ck(clk), .q(
        m1Inputs[125]) );
  dp_1 \INPUTSRAM/q_reg[126]  ( .ip(\INPUTSRAM/mem_i[7][14] ), .ck(clk), .q(
        m1Inputs[126]) );
  dp_1 \INPUTSRAM/q_reg[127]  ( .ip(\INPUTSRAM/mem_i[7][15] ), .ck(clk), .q(
        m1Inputs[127]) );
  dp_1 \INPUTSRAM/q_reg[128]  ( .ip(\INPUTSRAM/mem_i[8][0] ), .ck(clk), .q(
        m1Inputs[128]) );
  dp_1 \INPUTSRAM/q_reg[129]  ( .ip(\INPUTSRAM/mem_i[8][1] ), .ck(clk), .q(
        m1Inputs[129]) );
  dp_1 \INPUTSRAM/q_reg[142]  ( .ip(\INPUTSRAM/mem_i[8][14] ), .ck(clk), .q(
        m1Inputs[142]) );
  dp_1 \INPUTSRAM/q_reg[143]  ( .ip(\INPUTSRAM/mem_i[8][15] ), .ck(clk), .q(
        m1Inputs[143]) );
  dp_1 \INPUTSRAM/q_reg[144]  ( .ip(\INPUTSRAM/mem_i[9][0] ), .ck(clk), .q(
        m1Inputs[144]) );
  dp_1 \INPUTSRAM/q_reg[145]  ( .ip(\INPUTSRAM/mem_i[9][1] ), .ck(clk), .q(
        m1Inputs[145]) );
  dp_1 \INPUTSRAM/q_reg[158]  ( .ip(\INPUTSRAM/mem_i[9][14] ), .ck(clk), .q(
        m1Inputs[158]) );
  dp_1 \INPUTSRAM/q_reg[159]  ( .ip(\INPUTSRAM/mem_i[9][15] ), .ck(clk), .q(
        m1Inputs[159]) );
  dp_1 \CNTRL/count_20Q_reg[4]  ( .ip(n4111), .ck(clk), .q(
        \CNTRL/count_20Q [4]) );
  dp_1 \CNTRL/count_10Q_reg[3]  ( .ip(n4095), .ck(clk), .q(
        \CNTRL/count_10Q [3]) );
  dp_1 \CNTRL/currentState_reg[0]  ( .ip(n4107), .ck(clk), .q(
        \CNTRL/currentState [0]) );
  dp_1 \CNTRL/count_layer1_200Q_reg[7]  ( .ip(n4087), .ck(clk), .q(
        \CNTRL/count_layer1_200Q [7]) );
  dp_1 \CNTRL/count_layer1_784Q_reg[9]  ( .ip(\CNTRL/N242 ), .ck(clk), .q(
        \CNTRL/count_layer1_784Q [9]) );
  dp_1 \CNTRL/currentState_reg[1]  ( .ip(n4108), .ck(clk), .q(
        \CNTRL/currentState [1]) );
  dp_1 \CNTRL/currentState_reg[2]  ( .ip(n4109), .ck(clk), .q(
        \CNTRL/currentState [2]) );
  dp_1 \CNTRL/count_20Q_reg[0]  ( .ip(n4106), .ck(clk), .q(
        \CNTRL/count_20Q [0]) );
  dp_1 \CNTRL/count_20Q_reg[1]  ( .ip(n4105), .ck(clk), .q(
        \CNTRL/count_20Q [1]) );
  dp_1 \CNTRL/count_20Q_reg[2]  ( .ip(n4104), .ck(clk), .q(
        \CNTRL/count_20Q [2]) );
  dp_1 \CNTRL/count_20Q_reg[3]  ( .ip(n4103), .ck(clk), .q(
        \CNTRL/count_20Q [3]) );
  dp_1 \CNTRL/count_10Q_reg[0]  ( .ip(n4098), .ck(clk), .q(
        \CNTRL/count_10Q [0]) );
  dp_1 \CNTRL/count_10Q_reg[1]  ( .ip(n4097), .ck(clk), .q(
        \CNTRL/count_10Q [1]) );
  dp_1 \CNTRL/count_10Q_reg[2]  ( .ip(n4096), .ck(clk), .q(
        \CNTRL/count_10Q [2]) );
  dp_1 \CNTRL/count_layer1_784Q_reg[0]  ( .ip(\CNTRL/N233 ), .ck(clk), .q(
        \CNTRL/count_layer1_784Q [0]) );
  dp_1 \CNTRL/count_layer1_784Q_reg[1]  ( .ip(\CNTRL/N234 ), .ck(clk), .q(
        \CNTRL/count_layer1_784Q [1]) );
  dp_1 \CNTRL/count_layer1_784Q_reg[2]  ( .ip(\CNTRL/N235 ), .ck(clk), .q(
        \CNTRL/count_layer1_784Q [2]) );
  dp_1 \CNTRL/count_layer1_784Q_reg[3]  ( .ip(\CNTRL/N236 ), .ck(clk), .q(
        \CNTRL/count_layer1_784Q [3]) );
  dp_1 \CNTRL/count_layer1_784Q_reg[4]  ( .ip(\CNTRL/N237 ), .ck(clk), .q(
        \CNTRL/count_layer1_784Q [4]) );
  dp_1 \CNTRL/count_layer1_784Q_reg[5]  ( .ip(\CNTRL/N238 ), .ck(clk), .q(
        \CNTRL/count_layer1_784Q [5]) );
  dp_1 \CNTRL/count_layer1_784Q_reg[6]  ( .ip(\CNTRL/N239 ), .ck(clk), .q(
        \CNTRL/count_layer1_784Q [6]) );
  dp_1 \CNTRL/count_layer1_784Q_reg[7]  ( .ip(\CNTRL/N240 ), .ck(clk), .q(
        \CNTRL/count_layer1_784Q [7]) );
  dp_1 \CNTRL/count_layer1_784Q_reg[8]  ( .ip(\CNTRL/N241 ), .ck(clk), .q(
        \CNTRL/count_layer1_784Q [8]) );
  dp_1 \CNTRL/count_layer1_200Q_reg[1]  ( .ip(n4094), .ck(clk), .q(
        \CNTRL/count_layer1_200Q [1]) );
  dp_1 \CNTRL/count_layer1_200Q_reg[0]  ( .ip(n4093), .ck(clk), .q(
        \CNTRL/count_layer1_200Q [0]) );
  dp_1 \CNTRL/count_layer1_200Q_reg[2]  ( .ip(n4092), .ck(clk), .q(
        \CNTRL/count_layer1_200Q [2]) );
  dp_1 \CNTRL/count_layer1_200Q_reg[3]  ( .ip(n4091), .ck(clk), .q(
        \CNTRL/count_layer1_200Q [3]) );
  dp_1 \CNTRL/count_layer1_200Q_reg[4]  ( .ip(n4090), .ck(clk), .q(
        \CNTRL/count_layer1_200Q [4]) );
  dp_1 \CNTRL/count_layer1_200Q_reg[5]  ( .ip(n4089), .ck(clk), .q(
        \CNTRL/count_layer1_200Q [5]) );
  dp_1 \CNTRL/count_layer1_200Q_reg[6]  ( .ip(n4088), .ck(clk), .q(
        \CNTRL/count_layer1_200Q [6]) );
  dp_1 \CNTRL/count_10_2Q_reg[0]  ( .ip(n4102), .ck(clk), .q(
        \CNTRL/count_10_2Q [0]) );
  dp_1 \CNTRL/count_10_2Q_reg[1]  ( .ip(n4101), .ck(clk), .q(
        \CNTRL/count_10_2Q [1]) );
  dp_1 \CNTRL/count_10_2Q_reg[2]  ( .ip(n4100), .ck(clk), .q(
        \CNTRL/count_10_2Q [2]) );
  dp_1 \CNTRL/count_10_2Q_reg[3]  ( .ip(n4099), .ck(clk), .q(
        \CNTRL/count_10_2Q [3]) );
  dp_1 \ROUTEDATA/DataToM2_reg[0]  ( .ip(n4086), .ck(clk), .q(m2DataIn[0]) );
  dp_1 \ROUTEDATA/DataToM2_reg[1]  ( .ip(n4085), .ck(clk), .q(m2DataIn[1]) );
  dp_1 \ROUTEDATA/DataToM2_reg[2]  ( .ip(n4084), .ck(clk), .q(m2DataIn[2]) );
  dp_1 \ROUTEDATA/DataToM2_reg[3]  ( .ip(n4083), .ck(clk), .q(m2DataIn[3]) );
  dp_1 \ROUTEDATA/DataToM2_reg[4]  ( .ip(n4082), .ck(clk), .q(m2DataIn[4]) );
  dp_1 \ROUTEDATA/DataToM2_reg[5]  ( .ip(n4081), .ck(clk), .q(m2DataIn[5]) );
  dp_1 \ROUTEDATA/DataToM2_reg[6]  ( .ip(n4080), .ck(clk), .q(m2DataIn[6]) );
  dp_1 \ROUTEDATA/DataToM2_reg[7]  ( .ip(n4079), .ck(clk), .q(m2DataIn[7]) );
  dp_1 \ROUTEDATA/DataToM2_reg[8]  ( .ip(n4078), .ck(clk), .q(m2DataIn[8]) );
  dp_1 \ROUTEDATA/DataToM2_reg[9]  ( .ip(n4077), .ck(clk), .q(m2DataIn[9]) );
  dp_1 \ROUTEDATA/DataToM2_reg[10]  ( .ip(n4076), .ck(clk), .q(m2DataIn[10])
         );
  dp_1 \ROUTEDATA/DataToM2_reg[11]  ( .ip(n4075), .ck(clk), .q(m2DataIn[11])
         );
  dp_1 \ROUTEDATA/DataToM2_reg[12]  ( .ip(n4074), .ck(clk), .q(m2DataIn[12])
         );
  dp_1 \ROUTEDATA/DataToM2_reg[13]  ( .ip(n4073), .ck(clk), .q(m2DataIn[13])
         );
  dp_1 \ROUTEDATA/DataToM2_reg[14]  ( .ip(n4072), .ck(clk), .q(m2DataIn[14])
         );
  dp_1 \ROUTEDATA/DataToM2_reg[15]  ( .ip(n4071), .ck(clk), .q(m2DataIn[15])
         );
  dp_1 \WEIGHT_2/mem_w2_reg[0][0]  ( .ip(n4070), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][0] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][1]  ( .ip(n4069), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][1] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][2]  ( .ip(n4068), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][2] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][3]  ( .ip(n4067), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][3] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][4]  ( .ip(n4066), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][4] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][5]  ( .ip(n4065), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][5] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][6]  ( .ip(n4064), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][6] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][7]  ( .ip(n4063), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][7] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][8]  ( .ip(n4062), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][8] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][9]  ( .ip(n4061), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][9] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][10]  ( .ip(n4060), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][10] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][11]  ( .ip(n4059), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][11] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][12]  ( .ip(n4058), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][12] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][13]  ( .ip(n4057), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][13] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][14]  ( .ip(n4056), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][14] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[0][15]  ( .ip(n4055), .ck(clk), .q(
        \WEIGHT_2/mem_w2[0][15] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][0]  ( .ip(n4054), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][0] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][1]  ( .ip(n4053), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][1] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][2]  ( .ip(n4052), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][2] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][3]  ( .ip(n4051), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][3] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][4]  ( .ip(n4050), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][4] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][5]  ( .ip(n4049), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][5] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][6]  ( .ip(n4048), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][6] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][7]  ( .ip(n4047), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][7] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][8]  ( .ip(n4046), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][8] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][9]  ( .ip(n4045), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][9] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][10]  ( .ip(n4044), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][10] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][11]  ( .ip(n4043), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][11] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][12]  ( .ip(n4042), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][12] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][13]  ( .ip(n4041), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][13] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][14]  ( .ip(n4040), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][14] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[1][15]  ( .ip(n4039), .ck(clk), .q(
        \WEIGHT_2/mem_w2[1][15] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][0]  ( .ip(n4038), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][0] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][1]  ( .ip(n4037), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][1] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][2]  ( .ip(n4036), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][2] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][3]  ( .ip(n4035), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][3] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][4]  ( .ip(n4034), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][4] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][5]  ( .ip(n4033), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][5] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][6]  ( .ip(n4032), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][6] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][7]  ( .ip(n4031), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][7] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][8]  ( .ip(n4030), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][8] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][9]  ( .ip(n4029), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][9] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][10]  ( .ip(n4028), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][10] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][11]  ( .ip(n4027), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][11] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][12]  ( .ip(n4026), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][12] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][13]  ( .ip(n4025), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][13] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][14]  ( .ip(n4024), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][14] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[2][15]  ( .ip(n4023), .ck(clk), .q(
        \WEIGHT_2/mem_w2[2][15] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][0]  ( .ip(n4022), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][0] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][1]  ( .ip(n4021), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][1] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][2]  ( .ip(n4020), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][2] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][3]  ( .ip(n4019), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][3] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][4]  ( .ip(n4018), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][4] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][5]  ( .ip(n4017), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][5] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][6]  ( .ip(n4016), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][6] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][7]  ( .ip(n4015), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][7] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][8]  ( .ip(n4014), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][8] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][9]  ( .ip(n4013), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][9] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][10]  ( .ip(n4012), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][10] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][11]  ( .ip(n4011), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][11] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][12]  ( .ip(n4010), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][12] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][13]  ( .ip(n4009), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][13] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][14]  ( .ip(n4008), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][14] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[3][15]  ( .ip(n4007), .ck(clk), .q(
        \WEIGHT_2/mem_w2[3][15] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][0]  ( .ip(n4006), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][0] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][1]  ( .ip(n4005), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][1] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][2]  ( .ip(n4004), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][2] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][3]  ( .ip(n4003), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][3] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][4]  ( .ip(n4002), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][4] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][5]  ( .ip(n4001), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][5] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][6]  ( .ip(n4000), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][6] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][7]  ( .ip(n3999), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][7] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][8]  ( .ip(n3998), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][8] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][9]  ( .ip(n3997), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][9] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][10]  ( .ip(n3996), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][10] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][11]  ( .ip(n3995), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][11] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][12]  ( .ip(n3994), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][12] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][13]  ( .ip(n3993), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][13] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][14]  ( .ip(n3992), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][14] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[4][15]  ( .ip(n3991), .ck(clk), .q(
        \WEIGHT_2/mem_w2[4][15] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][0]  ( .ip(n3990), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][0] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][1]  ( .ip(n3989), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][1] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][2]  ( .ip(n3988), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][2] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][3]  ( .ip(n3987), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][3] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][4]  ( .ip(n3986), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][4] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][5]  ( .ip(n3985), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][5] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][6]  ( .ip(n3984), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][6] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][7]  ( .ip(n3983), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][7] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][8]  ( .ip(n3982), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][8] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][9]  ( .ip(n3981), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][9] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][10]  ( .ip(n3980), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][10] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][11]  ( .ip(n3979), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][11] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][12]  ( .ip(n3978), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][12] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][13]  ( .ip(n3977), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][13] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][14]  ( .ip(n3976), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][14] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[5][15]  ( .ip(n3975), .ck(clk), .q(
        \WEIGHT_2/mem_w2[5][15] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][0]  ( .ip(n3974), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][0] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][1]  ( .ip(n3973), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][1] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][2]  ( .ip(n3972), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][2] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][3]  ( .ip(n3971), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][3] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][4]  ( .ip(n3970), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][4] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][5]  ( .ip(n3969), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][5] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][6]  ( .ip(n3968), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][6] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][7]  ( .ip(n3967), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][7] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][8]  ( .ip(n3966), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][8] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][9]  ( .ip(n3965), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][9] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][10]  ( .ip(n3964), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][10] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][11]  ( .ip(n3963), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][11] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][12]  ( .ip(n3962), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][12] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][13]  ( .ip(n3961), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][13] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][14]  ( .ip(n3960), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][14] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[6][15]  ( .ip(n3959), .ck(clk), .q(
        \WEIGHT_2/mem_w2[6][15] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][0]  ( .ip(n3958), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][0] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][1]  ( .ip(n3957), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][1] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][2]  ( .ip(n3956), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][2] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][3]  ( .ip(n3955), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][3] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][4]  ( .ip(n3954), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][4] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][5]  ( .ip(n3953), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][5] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][6]  ( .ip(n3952), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][6] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][7]  ( .ip(n3951), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][7] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][8]  ( .ip(n3950), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][8] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][9]  ( .ip(n3949), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][9] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][10]  ( .ip(n3948), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][10] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][11]  ( .ip(n3947), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][11] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][12]  ( .ip(n3946), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][12] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][13]  ( .ip(n3945), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][13] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][14]  ( .ip(n3944), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][14] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[7][15]  ( .ip(n3943), .ck(clk), .q(
        \WEIGHT_2/mem_w2[7][15] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][0]  ( .ip(n3942), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][0] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][1]  ( .ip(n3941), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][1] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][2]  ( .ip(n3940), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][2] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][3]  ( .ip(n3939), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][3] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][4]  ( .ip(n3938), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][4] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][5]  ( .ip(n3937), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][5] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][6]  ( .ip(n3936), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][6] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][7]  ( .ip(n3935), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][7] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][8]  ( .ip(n3934), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][8] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][9]  ( .ip(n3933), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][9] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][10]  ( .ip(n3932), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][10] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][11]  ( .ip(n3931), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][11] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][12]  ( .ip(n3930), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][12] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][13]  ( .ip(n3929), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][13] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][14]  ( .ip(n3928), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][14] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[8][15]  ( .ip(n3927), .ck(clk), .q(
        \WEIGHT_2/mem_w2[8][15] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][0]  ( .ip(n3926), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][0] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][1]  ( .ip(n3925), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][1] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][2]  ( .ip(n3924), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][2] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][3]  ( .ip(n3923), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][3] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][4]  ( .ip(n3922), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][4] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][5]  ( .ip(n3921), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][5] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][6]  ( .ip(n3920), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][6] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][7]  ( .ip(n3919), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][7] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][8]  ( .ip(n3918), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][8] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][9]  ( .ip(n3917), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][9] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][10]  ( .ip(n3916), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][10] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][11]  ( .ip(n3915), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][11] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][12]  ( .ip(n3914), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][12] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][13]  ( .ip(n3913), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][13] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][14]  ( .ip(n3912), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][14] ) );
  dp_1 \WEIGHT_2/mem_w2_reg[9][15]  ( .ip(n3911), .ck(clk), .q(
        \WEIGHT_2/mem_w2[9][15] ) );
  dp_1 \ANSWER/rdata_reg[0]  ( .ip(\ANSWER/N487 ), .ck(clk), .q(rdata[0]) );
  dp_1 \ANSWER/rdata_reg[1]  ( .ip(\ANSWER/N486 ), .ck(clk), .q(rdata[1]) );
  dp_1 \ANSWER/rdata_reg[2]  ( .ip(\ANSWER/N485 ), .ck(clk), .q(rdata[2]) );
  dp_1 \ANSWER/rdata_reg[3]  ( .ip(\ANSWER/N484 ), .ck(clk), .q(rdata[3]) );
  dp_1 \ANSWER/rdata_reg[4]  ( .ip(\ANSWER/N483 ), .ck(clk), .q(rdata[4]) );
  dp_1 \ANSWER/rdata_reg[5]  ( .ip(\ANSWER/N482 ), .ck(clk), .q(rdata[5]) );
  dp_1 \ANSWER/rdata_reg[6]  ( .ip(\ANSWER/N481 ), .ck(clk), .q(rdata[6]) );
  dp_1 \ANSWER/rdata_reg[7]  ( .ip(\ANSWER/N480 ), .ck(clk), .q(rdata[7]) );
  dp_1 \ANSWER/rdata_reg[8]  ( .ip(\ANSWER/N479 ), .ck(clk), .q(rdata[8]) );
  dp_1 \ANSWER/rdata_reg[9]  ( .ip(\ANSWER/N478 ), .ck(clk), .q(rdata[9]) );
  dp_1 \ANSWER/rdata_reg[10]  ( .ip(\ANSWER/N477 ), .ck(clk), .q(rdata[10]) );
  dp_1 \ANSWER/rdata_reg[11]  ( .ip(\ANSWER/N476 ), .ck(clk), .q(rdata[11]) );
  dp_1 \ANSWER/rdata_reg[12]  ( .ip(\ANSWER/N475 ), .ck(clk), .q(rdata[12]) );
  dp_1 \ANSWER/rdata_reg[13]  ( .ip(\ANSWER/N474 ), .ck(clk), .q(rdata[13]) );
  dp_1 \ANSWER/rdata_reg[14]  ( .ip(\ANSWER/N473 ), .ck(clk), .q(rdata[14]) );
  dp_1 \ANSWER/rdata_reg[15]  ( .ip(\ANSWER/N472 ), .ck(clk), .q(rdata[15]) );
  dp_1 \SIGMOID/sign_bit_reg  ( .ip(n18918), .ck(clk), .q(\SIGMOID/sign_bit )
         );
  dp_1 \ANSWER/mem_reg[0][0][8]  ( .ip(n3102), .ck(clk), .q(
        \ANSWER/mem[0][0][8] ) );
  dp_1 \ANSWER/mem_reg[0][1][8]  ( .ip(n3101), .ck(clk), .q(
        \ANSWER/mem[0][1][8] ) );
  dp_1 \ANSWER/mem_reg[0][2][8]  ( .ip(n3100), .ck(clk), .q(
        \ANSWER/mem[0][2][8] ) );
  dp_1 \ANSWER/mem_reg[0][3][8]  ( .ip(n3099), .ck(clk), .q(
        \ANSWER/mem[0][3][8] ) );
  dp_1 \ANSWER/mem_reg[0][4][8]  ( .ip(n3098), .ck(clk), .q(
        \ANSWER/mem[0][4][8] ) );
  dp_1 \ANSWER/mem_reg[0][5][8]  ( .ip(n3097), .ck(clk), .q(
        \ANSWER/mem[0][5][8] ) );
  dp_1 \ANSWER/mem_reg[0][6][8]  ( .ip(n3096), .ck(clk), .q(
        \ANSWER/mem[0][6][8] ) );
  dp_1 \ANSWER/mem_reg[0][7][8]  ( .ip(n3095), .ck(clk), .q(
        \ANSWER/mem[0][7][8] ) );
  dp_1 \ANSWER/mem_reg[0][8][8]  ( .ip(n3094), .ck(clk), .q(
        \ANSWER/mem[0][8][8] ) );
  dp_1 \ANSWER/mem_reg[0][9][8]  ( .ip(n3093), .ck(clk), .q(
        \ANSWER/mem[0][9][8] ) );
  dp_1 \ANSWER/mem_reg[1][0][8]  ( .ip(n3092), .ck(clk), .q(
        \ANSWER/mem[1][0][8] ) );
  dp_1 \ANSWER/mem_reg[1][1][8]  ( .ip(n3091), .ck(clk), .q(
        \ANSWER/mem[1][1][8] ) );
  dp_1 \ANSWER/mem_reg[1][2][8]  ( .ip(n3090), .ck(clk), .q(
        \ANSWER/mem[1][2][8] ) );
  dp_1 \ANSWER/mem_reg[1][3][8]  ( .ip(n3089), .ck(clk), .q(
        \ANSWER/mem[1][3][8] ) );
  dp_1 \ANSWER/mem_reg[1][4][8]  ( .ip(n3088), .ck(clk), .q(
        \ANSWER/mem[1][4][8] ) );
  dp_1 \ANSWER/mem_reg[1][5][8]  ( .ip(n3087), .ck(clk), .q(
        \ANSWER/mem[1][5][8] ) );
  dp_1 \ANSWER/mem_reg[1][6][8]  ( .ip(n3086), .ck(clk), .q(
        \ANSWER/mem[1][6][8] ) );
  dp_1 \ANSWER/mem_reg[1][7][8]  ( .ip(n3085), .ck(clk), .q(
        \ANSWER/mem[1][7][8] ) );
  dp_1 \ANSWER/mem_reg[1][8][8]  ( .ip(n3084), .ck(clk), .q(
        \ANSWER/mem[1][8][8] ) );
  dp_1 \ANSWER/mem_reg[1][9][8]  ( .ip(n3083), .ck(clk), .q(
        \ANSWER/mem[1][9][8] ) );
  dp_1 \ANSWER/mem_reg[2][0][8]  ( .ip(n3082), .ck(clk), .q(
        \ANSWER/mem[2][0][8] ) );
  dp_1 \ANSWER/mem_reg[2][1][8]  ( .ip(n3081), .ck(clk), .q(
        \ANSWER/mem[2][1][8] ) );
  dp_1 \ANSWER/mem_reg[2][2][8]  ( .ip(n3080), .ck(clk), .q(
        \ANSWER/mem[2][2][8] ) );
  dp_1 \ANSWER/mem_reg[2][3][8]  ( .ip(n3079), .ck(clk), .q(
        \ANSWER/mem[2][3][8] ) );
  dp_1 \ANSWER/mem_reg[2][4][8]  ( .ip(n3078), .ck(clk), .q(
        \ANSWER/mem[2][4][8] ) );
  dp_1 \ANSWER/mem_reg[2][5][8]  ( .ip(n3077), .ck(clk), .q(
        \ANSWER/mem[2][5][8] ) );
  dp_1 \ANSWER/mem_reg[2][6][8]  ( .ip(n3076), .ck(clk), .q(
        \ANSWER/mem[2][6][8] ) );
  dp_1 \ANSWER/mem_reg[2][7][8]  ( .ip(n3075), .ck(clk), .q(
        \ANSWER/mem[2][7][8] ) );
  dp_1 \ANSWER/mem_reg[2][8][8]  ( .ip(n3074), .ck(clk), .q(
        \ANSWER/mem[2][8][8] ) );
  dp_1 \ANSWER/mem_reg[2][9][8]  ( .ip(n3073), .ck(clk), .q(
        \ANSWER/mem[2][9][8] ) );
  dp_1 \ANSWER/mem_reg[3][0][8]  ( .ip(n3072), .ck(clk), .q(
        \ANSWER/mem[3][0][8] ) );
  dp_1 \ANSWER/mem_reg[3][1][8]  ( .ip(n3071), .ck(clk), .q(
        \ANSWER/mem[3][1][8] ) );
  dp_1 \ANSWER/mem_reg[3][2][8]  ( .ip(n3070), .ck(clk), .q(
        \ANSWER/mem[3][2][8] ) );
  dp_1 \ANSWER/mem_reg[3][3][8]  ( .ip(n3069), .ck(clk), .q(
        \ANSWER/mem[3][3][8] ) );
  dp_1 \ANSWER/mem_reg[3][4][8]  ( .ip(n3068), .ck(clk), .q(
        \ANSWER/mem[3][4][8] ) );
  dp_1 \ANSWER/mem_reg[3][5][8]  ( .ip(n3067), .ck(clk), .q(
        \ANSWER/mem[3][5][8] ) );
  dp_1 \ANSWER/mem_reg[3][6][8]  ( .ip(n3066), .ck(clk), .q(
        \ANSWER/mem[3][6][8] ) );
  dp_1 \ANSWER/mem_reg[3][7][8]  ( .ip(n3065), .ck(clk), .q(
        \ANSWER/mem[3][7][8] ) );
  dp_1 \ANSWER/mem_reg[3][8][8]  ( .ip(n3064), .ck(clk), .q(
        \ANSWER/mem[3][8][8] ) );
  dp_1 \ANSWER/mem_reg[3][9][8]  ( .ip(n3063), .ck(clk), .q(
        \ANSWER/mem[3][9][8] ) );
  dp_1 \ANSWER/mem_reg[4][0][8]  ( .ip(n3062), .ck(clk), .q(
        \ANSWER/mem[4][0][8] ) );
  dp_1 \ANSWER/mem_reg[4][1][8]  ( .ip(n3061), .ck(clk), .q(
        \ANSWER/mem[4][1][8] ) );
  dp_1 \ANSWER/mem_reg[4][2][8]  ( .ip(n3060), .ck(clk), .q(
        \ANSWER/mem[4][2][8] ) );
  dp_1 \ANSWER/mem_reg[4][3][8]  ( .ip(n3059), .ck(clk), .q(
        \ANSWER/mem[4][3][8] ) );
  dp_1 \ANSWER/mem_reg[4][4][8]  ( .ip(n3058), .ck(clk), .q(
        \ANSWER/mem[4][4][8] ) );
  dp_1 \ANSWER/mem_reg[4][5][8]  ( .ip(n3057), .ck(clk), .q(
        \ANSWER/mem[4][5][8] ) );
  dp_1 \ANSWER/mem_reg[4][6][8]  ( .ip(n3056), .ck(clk), .q(
        \ANSWER/mem[4][6][8] ) );
  dp_1 \ANSWER/mem_reg[4][7][8]  ( .ip(n3055), .ck(clk), .q(
        \ANSWER/mem[4][7][8] ) );
  dp_1 \ANSWER/mem_reg[4][8][8]  ( .ip(n3054), .ck(clk), .q(
        \ANSWER/mem[4][8][8] ) );
  dp_1 \ANSWER/mem_reg[4][9][8]  ( .ip(n3053), .ck(clk), .q(
        \ANSWER/mem[4][9][8] ) );
  dp_1 \ANSWER/mem_reg[5][0][8]  ( .ip(n3052), .ck(clk), .q(
        \ANSWER/mem[5][0][8] ) );
  dp_1 \ANSWER/mem_reg[5][1][8]  ( .ip(n3051), .ck(clk), .q(
        \ANSWER/mem[5][1][8] ) );
  dp_1 \ANSWER/mem_reg[5][2][8]  ( .ip(n3050), .ck(clk), .q(
        \ANSWER/mem[5][2][8] ) );
  dp_1 \ANSWER/mem_reg[5][3][8]  ( .ip(n3049), .ck(clk), .q(
        \ANSWER/mem[5][3][8] ) );
  dp_1 \ANSWER/mem_reg[5][4][8]  ( .ip(n3048), .ck(clk), .q(
        \ANSWER/mem[5][4][8] ) );
  dp_1 \ANSWER/mem_reg[5][5][8]  ( .ip(n3047), .ck(clk), .q(
        \ANSWER/mem[5][5][8] ) );
  dp_1 \ANSWER/mem_reg[5][6][8]  ( .ip(n3046), .ck(clk), .q(
        \ANSWER/mem[5][6][8] ) );
  dp_1 \ANSWER/mem_reg[5][7][8]  ( .ip(n3045), .ck(clk), .q(
        \ANSWER/mem[5][7][8] ) );
  dp_1 \ANSWER/mem_reg[5][8][8]  ( .ip(n3044), .ck(clk), .q(
        \ANSWER/mem[5][8][8] ) );
  dp_1 \ANSWER/mem_reg[5][9][8]  ( .ip(n3043), .ck(clk), .q(
        \ANSWER/mem[5][9][8] ) );
  dp_1 \ANSWER/mem_reg[6][0][8]  ( .ip(n3042), .ck(clk), .q(
        \ANSWER/mem[6][0][8] ) );
  dp_1 \ANSWER/mem_reg[6][1][8]  ( .ip(n3041), .ck(clk), .q(
        \ANSWER/mem[6][1][8] ) );
  dp_1 \ANSWER/mem_reg[6][2][8]  ( .ip(n3040), .ck(clk), .q(
        \ANSWER/mem[6][2][8] ) );
  dp_1 \ANSWER/mem_reg[6][3][8]  ( .ip(n3039), .ck(clk), .q(
        \ANSWER/mem[6][3][8] ) );
  dp_1 \ANSWER/mem_reg[6][4][8]  ( .ip(n3038), .ck(clk), .q(
        \ANSWER/mem[6][4][8] ) );
  dp_1 \ANSWER/mem_reg[6][5][8]  ( .ip(n3037), .ck(clk), .q(
        \ANSWER/mem[6][5][8] ) );
  dp_1 \ANSWER/mem_reg[6][6][8]  ( .ip(n3036), .ck(clk), .q(
        \ANSWER/mem[6][6][8] ) );
  dp_1 \ANSWER/mem_reg[6][7][8]  ( .ip(n3035), .ck(clk), .q(
        \ANSWER/mem[6][7][8] ) );
  dp_1 \ANSWER/mem_reg[6][8][8]  ( .ip(n3034), .ck(clk), .q(
        \ANSWER/mem[6][8][8] ) );
  dp_1 \ANSWER/mem_reg[6][9][8]  ( .ip(n3033), .ck(clk), .q(
        \ANSWER/mem[6][9][8] ) );
  dp_1 \ANSWER/mem_reg[7][0][8]  ( .ip(n3032), .ck(clk), .q(
        \ANSWER/mem[7][0][8] ) );
  dp_1 \ANSWER/mem_reg[7][1][8]  ( .ip(n3031), .ck(clk), .q(
        \ANSWER/mem[7][1][8] ) );
  dp_1 \ANSWER/mem_reg[7][2][8]  ( .ip(n3030), .ck(clk), .q(
        \ANSWER/mem[7][2][8] ) );
  dp_1 \ANSWER/mem_reg[7][3][8]  ( .ip(n3029), .ck(clk), .q(
        \ANSWER/mem[7][3][8] ) );
  dp_1 \ANSWER/mem_reg[7][4][8]  ( .ip(n3028), .ck(clk), .q(
        \ANSWER/mem[7][4][8] ) );
  dp_1 \ANSWER/mem_reg[7][5][8]  ( .ip(n3027), .ck(clk), .q(
        \ANSWER/mem[7][5][8] ) );
  dp_1 \ANSWER/mem_reg[7][6][8]  ( .ip(n3026), .ck(clk), .q(
        \ANSWER/mem[7][6][8] ) );
  dp_1 \ANSWER/mem_reg[7][7][8]  ( .ip(n3025), .ck(clk), .q(
        \ANSWER/mem[7][7][8] ) );
  dp_1 \ANSWER/mem_reg[7][8][8]  ( .ip(n3024), .ck(clk), .q(
        \ANSWER/mem[7][8][8] ) );
  dp_1 \ANSWER/mem_reg[7][9][8]  ( .ip(n3023), .ck(clk), .q(
        \ANSWER/mem[7][9][8] ) );
  dp_1 \ANSWER/mem_reg[8][0][8]  ( .ip(n3022), .ck(clk), .q(
        \ANSWER/mem[8][0][8] ) );
  dp_1 \ANSWER/mem_reg[8][1][8]  ( .ip(n3021), .ck(clk), .q(
        \ANSWER/mem[8][1][8] ) );
  dp_1 \ANSWER/mem_reg[8][2][8]  ( .ip(n3020), .ck(clk), .q(
        \ANSWER/mem[8][2][8] ) );
  dp_1 \ANSWER/mem_reg[8][3][8]  ( .ip(n3019), .ck(clk), .q(
        \ANSWER/mem[8][3][8] ) );
  dp_1 \ANSWER/mem_reg[8][4][8]  ( .ip(n3018), .ck(clk), .q(
        \ANSWER/mem[8][4][8] ) );
  dp_1 \ANSWER/mem_reg[8][5][8]  ( .ip(n3017), .ck(clk), .q(
        \ANSWER/mem[8][5][8] ) );
  dp_1 \ANSWER/mem_reg[8][6][8]  ( .ip(n3016), .ck(clk), .q(
        \ANSWER/mem[8][6][8] ) );
  dp_1 \ANSWER/mem_reg[8][7][8]  ( .ip(n3015), .ck(clk), .q(
        \ANSWER/mem[8][7][8] ) );
  dp_1 \ANSWER/mem_reg[8][8][8]  ( .ip(n3014), .ck(clk), .q(
        \ANSWER/mem[8][8][8] ) );
  dp_1 \ANSWER/mem_reg[8][9][8]  ( .ip(n3013), .ck(clk), .q(
        \ANSWER/mem[8][9][8] ) );
  dp_1 \ANSWER/mem_reg[9][0][8]  ( .ip(n3012), .ck(clk), .q(
        \ANSWER/mem[9][0][8] ) );
  dp_1 \ANSWER/mem_reg[9][1][8]  ( .ip(n3011), .ck(clk), .q(
        \ANSWER/mem[9][1][8] ) );
  dp_1 \ANSWER/mem_reg[9][2][8]  ( .ip(n3010), .ck(clk), .q(
        \ANSWER/mem[9][2][8] ) );
  dp_1 \ANSWER/mem_reg[9][3][8]  ( .ip(n3009), .ck(clk), .q(
        \ANSWER/mem[9][3][8] ) );
  dp_1 \ANSWER/mem_reg[9][4][8]  ( .ip(n3008), .ck(clk), .q(
        \ANSWER/mem[9][4][8] ) );
  dp_1 \ANSWER/mem_reg[9][5][8]  ( .ip(n3007), .ck(clk), .q(
        \ANSWER/mem[9][5][8] ) );
  dp_1 \ANSWER/mem_reg[9][6][8]  ( .ip(n3006), .ck(clk), .q(
        \ANSWER/mem[9][6][8] ) );
  dp_1 \ANSWER/mem_reg[9][7][8]  ( .ip(n3005), .ck(clk), .q(
        \ANSWER/mem[9][7][8] ) );
  dp_1 \ANSWER/mem_reg[9][8][8]  ( .ip(n3004), .ck(clk), .q(
        \ANSWER/mem[9][8][8] ) );
  dp_1 \ANSWER/mem_reg[9][9][8]  ( .ip(n3003), .ck(clk), .q(
        \ANSWER/mem[9][9][8] ) );
  dp_1 \ANSWER/mem_reg[0][0][9]  ( .ip(n3002), .ck(clk), .q(
        \ANSWER/mem[0][0][9] ) );
  dp_1 \ANSWER/mem_reg[0][1][9]  ( .ip(n3001), .ck(clk), .q(
        \ANSWER/mem[0][1][9] ) );
  dp_1 \ANSWER/mem_reg[0][2][9]  ( .ip(n3000), .ck(clk), .q(
        \ANSWER/mem[0][2][9] ) );
  dp_1 \ANSWER/mem_reg[0][3][9]  ( .ip(n2999), .ck(clk), .q(
        \ANSWER/mem[0][3][9] ) );
  dp_1 \ANSWER/mem_reg[0][4][9]  ( .ip(n2998), .ck(clk), .q(
        \ANSWER/mem[0][4][9] ) );
  dp_1 \ANSWER/mem_reg[0][5][9]  ( .ip(n2997), .ck(clk), .q(
        \ANSWER/mem[0][5][9] ) );
  dp_1 \ANSWER/mem_reg[0][6][9]  ( .ip(n2996), .ck(clk), .q(
        \ANSWER/mem[0][6][9] ) );
  dp_1 \ANSWER/mem_reg[0][7][9]  ( .ip(n2995), .ck(clk), .q(
        \ANSWER/mem[0][7][9] ) );
  dp_1 \ANSWER/mem_reg[0][8][9]  ( .ip(n2994), .ck(clk), .q(
        \ANSWER/mem[0][8][9] ) );
  dp_1 \ANSWER/mem_reg[0][9][9]  ( .ip(n2993), .ck(clk), .q(
        \ANSWER/mem[0][9][9] ) );
  dp_1 \ANSWER/mem_reg[1][0][9]  ( .ip(n2992), .ck(clk), .q(
        \ANSWER/mem[1][0][9] ) );
  dp_1 \ANSWER/mem_reg[1][1][9]  ( .ip(n2991), .ck(clk), .q(
        \ANSWER/mem[1][1][9] ) );
  dp_1 \ANSWER/mem_reg[1][2][9]  ( .ip(n2990), .ck(clk), .q(
        \ANSWER/mem[1][2][9] ) );
  dp_1 \ANSWER/mem_reg[1][3][9]  ( .ip(n2989), .ck(clk), .q(
        \ANSWER/mem[1][3][9] ) );
  dp_1 \ANSWER/mem_reg[1][4][9]  ( .ip(n2988), .ck(clk), .q(
        \ANSWER/mem[1][4][9] ) );
  dp_1 \ANSWER/mem_reg[1][5][9]  ( .ip(n2987), .ck(clk), .q(
        \ANSWER/mem[1][5][9] ) );
  dp_1 \ANSWER/mem_reg[1][6][9]  ( .ip(n2986), .ck(clk), .q(
        \ANSWER/mem[1][6][9] ) );
  dp_1 \ANSWER/mem_reg[1][7][9]  ( .ip(n2985), .ck(clk), .q(
        \ANSWER/mem[1][7][9] ) );
  dp_1 \ANSWER/mem_reg[1][8][9]  ( .ip(n2984), .ck(clk), .q(
        \ANSWER/mem[1][8][9] ) );
  dp_1 \ANSWER/mem_reg[1][9][9]  ( .ip(n2983), .ck(clk), .q(
        \ANSWER/mem[1][9][9] ) );
  dp_1 \ANSWER/mem_reg[2][0][9]  ( .ip(n2982), .ck(clk), .q(
        \ANSWER/mem[2][0][9] ) );
  dp_1 \ANSWER/mem_reg[2][1][9]  ( .ip(n2981), .ck(clk), .q(
        \ANSWER/mem[2][1][9] ) );
  dp_1 \ANSWER/mem_reg[2][2][9]  ( .ip(n2980), .ck(clk), .q(
        \ANSWER/mem[2][2][9] ) );
  dp_1 \ANSWER/mem_reg[2][3][9]  ( .ip(n2979), .ck(clk), .q(
        \ANSWER/mem[2][3][9] ) );
  dp_1 \ANSWER/mem_reg[2][4][9]  ( .ip(n2978), .ck(clk), .q(
        \ANSWER/mem[2][4][9] ) );
  dp_1 \ANSWER/mem_reg[2][5][9]  ( .ip(n2977), .ck(clk), .q(
        \ANSWER/mem[2][5][9] ) );
  dp_1 \ANSWER/mem_reg[2][6][9]  ( .ip(n2976), .ck(clk), .q(
        \ANSWER/mem[2][6][9] ) );
  dp_1 \ANSWER/mem_reg[2][7][9]  ( .ip(n2975), .ck(clk), .q(
        \ANSWER/mem[2][7][9] ) );
  dp_1 \ANSWER/mem_reg[2][8][9]  ( .ip(n2974), .ck(clk), .q(
        \ANSWER/mem[2][8][9] ) );
  dp_1 \ANSWER/mem_reg[2][9][9]  ( .ip(n2973), .ck(clk), .q(
        \ANSWER/mem[2][9][9] ) );
  dp_1 \ANSWER/mem_reg[3][0][9]  ( .ip(n2972), .ck(clk), .q(
        \ANSWER/mem[3][0][9] ) );
  dp_1 \ANSWER/mem_reg[3][1][9]  ( .ip(n2971), .ck(clk), .q(
        \ANSWER/mem[3][1][9] ) );
  dp_1 \ANSWER/mem_reg[3][2][9]  ( .ip(n2970), .ck(clk), .q(
        \ANSWER/mem[3][2][9] ) );
  dp_1 \ANSWER/mem_reg[3][3][9]  ( .ip(n2969), .ck(clk), .q(
        \ANSWER/mem[3][3][9] ) );
  dp_1 \ANSWER/mem_reg[3][4][9]  ( .ip(n2968), .ck(clk), .q(
        \ANSWER/mem[3][4][9] ) );
  dp_1 \ANSWER/mem_reg[3][5][9]  ( .ip(n2967), .ck(clk), .q(
        \ANSWER/mem[3][5][9] ) );
  dp_1 \ANSWER/mem_reg[3][6][9]  ( .ip(n2966), .ck(clk), .q(
        \ANSWER/mem[3][6][9] ) );
  dp_1 \ANSWER/mem_reg[3][7][9]  ( .ip(n2965), .ck(clk), .q(
        \ANSWER/mem[3][7][9] ) );
  dp_1 \ANSWER/mem_reg[3][8][9]  ( .ip(n2964), .ck(clk), .q(
        \ANSWER/mem[3][8][9] ) );
  dp_1 \ANSWER/mem_reg[3][9][9]  ( .ip(n2963), .ck(clk), .q(
        \ANSWER/mem[3][9][9] ) );
  dp_1 \ANSWER/mem_reg[4][0][9]  ( .ip(n2962), .ck(clk), .q(
        \ANSWER/mem[4][0][9] ) );
  dp_1 \ANSWER/mem_reg[4][1][9]  ( .ip(n2961), .ck(clk), .q(
        \ANSWER/mem[4][1][9] ) );
  dp_1 \ANSWER/mem_reg[4][2][9]  ( .ip(n2960), .ck(clk), .q(
        \ANSWER/mem[4][2][9] ) );
  dp_1 \ANSWER/mem_reg[4][3][9]  ( .ip(n2959), .ck(clk), .q(
        \ANSWER/mem[4][3][9] ) );
  dp_1 \ANSWER/mem_reg[4][4][9]  ( .ip(n2958), .ck(clk), .q(
        \ANSWER/mem[4][4][9] ) );
  dp_1 \ANSWER/mem_reg[4][5][9]  ( .ip(n2957), .ck(clk), .q(
        \ANSWER/mem[4][5][9] ) );
  dp_1 \ANSWER/mem_reg[4][6][9]  ( .ip(n2956), .ck(clk), .q(
        \ANSWER/mem[4][6][9] ) );
  dp_1 \ANSWER/mem_reg[4][7][9]  ( .ip(n2955), .ck(clk), .q(
        \ANSWER/mem[4][7][9] ) );
  dp_1 \ANSWER/mem_reg[4][8][9]  ( .ip(n2954), .ck(clk), .q(
        \ANSWER/mem[4][8][9] ) );
  dp_1 \ANSWER/mem_reg[4][9][9]  ( .ip(n2953), .ck(clk), .q(
        \ANSWER/mem[4][9][9] ) );
  dp_1 \ANSWER/mem_reg[5][0][9]  ( .ip(n2952), .ck(clk), .q(
        \ANSWER/mem[5][0][9] ) );
  dp_1 \ANSWER/mem_reg[5][1][9]  ( .ip(n2951), .ck(clk), .q(
        \ANSWER/mem[5][1][9] ) );
  dp_1 \ANSWER/mem_reg[5][2][9]  ( .ip(n2950), .ck(clk), .q(
        \ANSWER/mem[5][2][9] ) );
  dp_1 \ANSWER/mem_reg[5][3][9]  ( .ip(n2949), .ck(clk), .q(
        \ANSWER/mem[5][3][9] ) );
  dp_1 \ANSWER/mem_reg[5][4][9]  ( .ip(n2948), .ck(clk), .q(
        \ANSWER/mem[5][4][9] ) );
  dp_1 \ANSWER/mem_reg[5][5][9]  ( .ip(n2947), .ck(clk), .q(
        \ANSWER/mem[5][5][9] ) );
  dp_1 \ANSWER/mem_reg[5][6][9]  ( .ip(n2946), .ck(clk), .q(
        \ANSWER/mem[5][6][9] ) );
  dp_1 \ANSWER/mem_reg[5][7][9]  ( .ip(n2945), .ck(clk), .q(
        \ANSWER/mem[5][7][9] ) );
  dp_1 \ANSWER/mem_reg[5][8][9]  ( .ip(n2944), .ck(clk), .q(
        \ANSWER/mem[5][8][9] ) );
  dp_1 \ANSWER/mem_reg[5][9][9]  ( .ip(n2943), .ck(clk), .q(
        \ANSWER/mem[5][9][9] ) );
  dp_1 \ANSWER/mem_reg[6][0][9]  ( .ip(n2942), .ck(clk), .q(
        \ANSWER/mem[6][0][9] ) );
  dp_1 \ANSWER/mem_reg[6][1][9]  ( .ip(n2941), .ck(clk), .q(
        \ANSWER/mem[6][1][9] ) );
  dp_1 \ANSWER/mem_reg[6][2][9]  ( .ip(n2940), .ck(clk), .q(
        \ANSWER/mem[6][2][9] ) );
  dp_1 \ANSWER/mem_reg[6][3][9]  ( .ip(n2939), .ck(clk), .q(
        \ANSWER/mem[6][3][9] ) );
  dp_1 \ANSWER/mem_reg[6][4][9]  ( .ip(n2938), .ck(clk), .q(
        \ANSWER/mem[6][4][9] ) );
  dp_1 \ANSWER/mem_reg[6][5][9]  ( .ip(n2937), .ck(clk), .q(
        \ANSWER/mem[6][5][9] ) );
  dp_1 \ANSWER/mem_reg[6][6][9]  ( .ip(n2936), .ck(clk), .q(
        \ANSWER/mem[6][6][9] ) );
  dp_1 \ANSWER/mem_reg[6][7][9]  ( .ip(n2935), .ck(clk), .q(
        \ANSWER/mem[6][7][9] ) );
  dp_1 \ANSWER/mem_reg[6][8][9]  ( .ip(n2934), .ck(clk), .q(
        \ANSWER/mem[6][8][9] ) );
  dp_1 \ANSWER/mem_reg[6][9][9]  ( .ip(n2933), .ck(clk), .q(
        \ANSWER/mem[6][9][9] ) );
  dp_1 \ANSWER/mem_reg[7][0][9]  ( .ip(n2932), .ck(clk), .q(
        \ANSWER/mem[7][0][9] ) );
  dp_1 \ANSWER/mem_reg[7][1][9]  ( .ip(n2931), .ck(clk), .q(
        \ANSWER/mem[7][1][9] ) );
  dp_1 \ANSWER/mem_reg[7][2][9]  ( .ip(n2930), .ck(clk), .q(
        \ANSWER/mem[7][2][9] ) );
  dp_1 \ANSWER/mem_reg[7][3][9]  ( .ip(n2929), .ck(clk), .q(
        \ANSWER/mem[7][3][9] ) );
  dp_1 \ANSWER/mem_reg[7][4][9]  ( .ip(n2928), .ck(clk), .q(
        \ANSWER/mem[7][4][9] ) );
  dp_1 \ANSWER/mem_reg[7][5][9]  ( .ip(n2927), .ck(clk), .q(
        \ANSWER/mem[7][5][9] ) );
  dp_1 \ANSWER/mem_reg[7][6][9]  ( .ip(n2926), .ck(clk), .q(
        \ANSWER/mem[7][6][9] ) );
  dp_1 \ANSWER/mem_reg[7][7][9]  ( .ip(n2925), .ck(clk), .q(
        \ANSWER/mem[7][7][9] ) );
  dp_1 \ANSWER/mem_reg[7][8][9]  ( .ip(n2924), .ck(clk), .q(
        \ANSWER/mem[7][8][9] ) );
  dp_1 \ANSWER/mem_reg[7][9][9]  ( .ip(n2923), .ck(clk), .q(
        \ANSWER/mem[7][9][9] ) );
  dp_1 \ANSWER/mem_reg[8][0][9]  ( .ip(n2922), .ck(clk), .q(
        \ANSWER/mem[8][0][9] ) );
  dp_1 \ANSWER/mem_reg[8][1][9]  ( .ip(n2921), .ck(clk), .q(
        \ANSWER/mem[8][1][9] ) );
  dp_1 \ANSWER/mem_reg[8][2][9]  ( .ip(n2920), .ck(clk), .q(
        \ANSWER/mem[8][2][9] ) );
  dp_1 \ANSWER/mem_reg[8][3][9]  ( .ip(n2919), .ck(clk), .q(
        \ANSWER/mem[8][3][9] ) );
  dp_1 \ANSWER/mem_reg[8][4][9]  ( .ip(n2918), .ck(clk), .q(
        \ANSWER/mem[8][4][9] ) );
  dp_1 \ANSWER/mem_reg[8][5][9]  ( .ip(n2917), .ck(clk), .q(
        \ANSWER/mem[8][5][9] ) );
  dp_1 \ANSWER/mem_reg[8][6][9]  ( .ip(n2916), .ck(clk), .q(
        \ANSWER/mem[8][6][9] ) );
  dp_1 \ANSWER/mem_reg[8][7][9]  ( .ip(n2915), .ck(clk), .q(
        \ANSWER/mem[8][7][9] ) );
  dp_1 \ANSWER/mem_reg[8][8][9]  ( .ip(n2914), .ck(clk), .q(
        \ANSWER/mem[8][8][9] ) );
  dp_1 \ANSWER/mem_reg[8][9][9]  ( .ip(n2913), .ck(clk), .q(
        \ANSWER/mem[8][9][9] ) );
  dp_1 \ANSWER/mem_reg[9][0][9]  ( .ip(n2912), .ck(clk), .q(
        \ANSWER/mem[9][0][9] ) );
  dp_1 \ANSWER/mem_reg[9][1][9]  ( .ip(n2911), .ck(clk), .q(
        \ANSWER/mem[9][1][9] ) );
  dp_1 \ANSWER/mem_reg[9][2][9]  ( .ip(n2910), .ck(clk), .q(
        \ANSWER/mem[9][2][9] ) );
  dp_1 \ANSWER/mem_reg[9][3][9]  ( .ip(n2909), .ck(clk), .q(
        \ANSWER/mem[9][3][9] ) );
  dp_1 \ANSWER/mem_reg[9][4][9]  ( .ip(n2908), .ck(clk), .q(
        \ANSWER/mem[9][4][9] ) );
  dp_1 \ANSWER/mem_reg[9][5][9]  ( .ip(n2907), .ck(clk), .q(
        \ANSWER/mem[9][5][9] ) );
  dp_1 \ANSWER/mem_reg[9][6][9]  ( .ip(n2906), .ck(clk), .q(
        \ANSWER/mem[9][6][9] ) );
  dp_1 \ANSWER/mem_reg[9][7][9]  ( .ip(n2905), .ck(clk), .q(
        \ANSWER/mem[9][7][9] ) );
  dp_1 \ANSWER/mem_reg[9][8][9]  ( .ip(n2904), .ck(clk), .q(
        \ANSWER/mem[9][8][9] ) );
  dp_1 \ANSWER/mem_reg[9][9][9]  ( .ip(n2903), .ck(clk), .q(
        \ANSWER/mem[9][9][9] ) );
  dp_1 \ANSWER/mem_reg[0][0][10]  ( .ip(n2902), .ck(clk), .q(
        \ANSWER/mem[0][0][10] ) );
  dp_1 \ANSWER/mem_reg[0][1][10]  ( .ip(n2901), .ck(clk), .q(
        \ANSWER/mem[0][1][10] ) );
  dp_1 \ANSWER/mem_reg[0][2][10]  ( .ip(n2900), .ck(clk), .q(
        \ANSWER/mem[0][2][10] ) );
  dp_1 \ANSWER/mem_reg[0][3][10]  ( .ip(n2899), .ck(clk), .q(
        \ANSWER/mem[0][3][10] ) );
  dp_1 \ANSWER/mem_reg[0][4][10]  ( .ip(n2898), .ck(clk), .q(
        \ANSWER/mem[0][4][10] ) );
  dp_1 \ANSWER/mem_reg[0][5][10]  ( .ip(n2897), .ck(clk), .q(
        \ANSWER/mem[0][5][10] ) );
  dp_1 \ANSWER/mem_reg[0][6][10]  ( .ip(n2896), .ck(clk), .q(
        \ANSWER/mem[0][6][10] ) );
  dp_1 \ANSWER/mem_reg[0][7][10]  ( .ip(n2895), .ck(clk), .q(
        \ANSWER/mem[0][7][10] ) );
  dp_1 \ANSWER/mem_reg[0][8][10]  ( .ip(n2894), .ck(clk), .q(
        \ANSWER/mem[0][8][10] ) );
  dp_1 \ANSWER/mem_reg[0][9][10]  ( .ip(n2893), .ck(clk), .q(
        \ANSWER/mem[0][9][10] ) );
  dp_1 \ANSWER/mem_reg[1][0][10]  ( .ip(n2892), .ck(clk), .q(
        \ANSWER/mem[1][0][10] ) );
  dp_1 \ANSWER/mem_reg[1][1][10]  ( .ip(n2891), .ck(clk), .q(
        \ANSWER/mem[1][1][10] ) );
  dp_1 \ANSWER/mem_reg[1][2][10]  ( .ip(n2890), .ck(clk), .q(
        \ANSWER/mem[1][2][10] ) );
  dp_1 \ANSWER/mem_reg[1][3][10]  ( .ip(n2889), .ck(clk), .q(
        \ANSWER/mem[1][3][10] ) );
  dp_1 \ANSWER/mem_reg[1][4][10]  ( .ip(n2888), .ck(clk), .q(
        \ANSWER/mem[1][4][10] ) );
  dp_1 \ANSWER/mem_reg[1][5][10]  ( .ip(n2887), .ck(clk), .q(
        \ANSWER/mem[1][5][10] ) );
  dp_1 \ANSWER/mem_reg[1][6][10]  ( .ip(n2886), .ck(clk), .q(
        \ANSWER/mem[1][6][10] ) );
  dp_1 \ANSWER/mem_reg[1][7][10]  ( .ip(n2885), .ck(clk), .q(
        \ANSWER/mem[1][7][10] ) );
  dp_1 \ANSWER/mem_reg[1][8][10]  ( .ip(n2884), .ck(clk), .q(
        \ANSWER/mem[1][8][10] ) );
  dp_1 \ANSWER/mem_reg[1][9][10]  ( .ip(n2883), .ck(clk), .q(
        \ANSWER/mem[1][9][10] ) );
  dp_1 \ANSWER/mem_reg[2][0][10]  ( .ip(n2882), .ck(clk), .q(
        \ANSWER/mem[2][0][10] ) );
  dp_1 \ANSWER/mem_reg[2][1][10]  ( .ip(n2881), .ck(clk), .q(
        \ANSWER/mem[2][1][10] ) );
  dp_1 \ANSWER/mem_reg[2][2][10]  ( .ip(n2880), .ck(clk), .q(
        \ANSWER/mem[2][2][10] ) );
  dp_1 \ANSWER/mem_reg[2][3][10]  ( .ip(n2879), .ck(clk), .q(
        \ANSWER/mem[2][3][10] ) );
  dp_1 \ANSWER/mem_reg[2][4][10]  ( .ip(n2878), .ck(clk), .q(
        \ANSWER/mem[2][4][10] ) );
  dp_1 \ANSWER/mem_reg[2][5][10]  ( .ip(n2877), .ck(clk), .q(
        \ANSWER/mem[2][5][10] ) );
  dp_1 \ANSWER/mem_reg[2][6][10]  ( .ip(n2876), .ck(clk), .q(
        \ANSWER/mem[2][6][10] ) );
  dp_1 \ANSWER/mem_reg[2][7][10]  ( .ip(n2875), .ck(clk), .q(
        \ANSWER/mem[2][7][10] ) );
  dp_1 \ANSWER/mem_reg[2][8][10]  ( .ip(n2874), .ck(clk), .q(
        \ANSWER/mem[2][8][10] ) );
  dp_1 \ANSWER/mem_reg[2][9][10]  ( .ip(n2873), .ck(clk), .q(
        \ANSWER/mem[2][9][10] ) );
  dp_1 \ANSWER/mem_reg[3][0][10]  ( .ip(n2872), .ck(clk), .q(
        \ANSWER/mem[3][0][10] ) );
  dp_1 \ANSWER/mem_reg[3][1][10]  ( .ip(n2871), .ck(clk), .q(
        \ANSWER/mem[3][1][10] ) );
  dp_1 \ANSWER/mem_reg[3][2][10]  ( .ip(n2870), .ck(clk), .q(
        \ANSWER/mem[3][2][10] ) );
  dp_1 \ANSWER/mem_reg[3][3][10]  ( .ip(n2869), .ck(clk), .q(
        \ANSWER/mem[3][3][10] ) );
  dp_1 \ANSWER/mem_reg[3][4][10]  ( .ip(n2868), .ck(clk), .q(
        \ANSWER/mem[3][4][10] ) );
  dp_1 \ANSWER/mem_reg[3][5][10]  ( .ip(n2867), .ck(clk), .q(
        \ANSWER/mem[3][5][10] ) );
  dp_1 \ANSWER/mem_reg[3][6][10]  ( .ip(n2866), .ck(clk), .q(
        \ANSWER/mem[3][6][10] ) );
  dp_1 \ANSWER/mem_reg[3][7][10]  ( .ip(n2865), .ck(clk), .q(
        \ANSWER/mem[3][7][10] ) );
  dp_1 \ANSWER/mem_reg[3][8][10]  ( .ip(n2864), .ck(clk), .q(
        \ANSWER/mem[3][8][10] ) );
  dp_1 \ANSWER/mem_reg[3][9][10]  ( .ip(n2863), .ck(clk), .q(
        \ANSWER/mem[3][9][10] ) );
  dp_1 \ANSWER/mem_reg[4][0][10]  ( .ip(n2862), .ck(clk), .q(
        \ANSWER/mem[4][0][10] ) );
  dp_1 \ANSWER/mem_reg[4][1][10]  ( .ip(n2861), .ck(clk), .q(
        \ANSWER/mem[4][1][10] ) );
  dp_1 \ANSWER/mem_reg[4][2][10]  ( .ip(n2860), .ck(clk), .q(
        \ANSWER/mem[4][2][10] ) );
  dp_1 \ANSWER/mem_reg[4][3][10]  ( .ip(n2859), .ck(clk), .q(
        \ANSWER/mem[4][3][10] ) );
  dp_1 \ANSWER/mem_reg[4][4][10]  ( .ip(n2858), .ck(clk), .q(
        \ANSWER/mem[4][4][10] ) );
  dp_1 \ANSWER/mem_reg[4][5][10]  ( .ip(n2857), .ck(clk), .q(
        \ANSWER/mem[4][5][10] ) );
  dp_1 \ANSWER/mem_reg[4][6][10]  ( .ip(n2856), .ck(clk), .q(
        \ANSWER/mem[4][6][10] ) );
  dp_1 \ANSWER/mem_reg[4][7][10]  ( .ip(n2855), .ck(clk), .q(
        \ANSWER/mem[4][7][10] ) );
  dp_1 \ANSWER/mem_reg[4][8][10]  ( .ip(n2854), .ck(clk), .q(
        \ANSWER/mem[4][8][10] ) );
  dp_1 \ANSWER/mem_reg[4][9][10]  ( .ip(n2853), .ck(clk), .q(
        \ANSWER/mem[4][9][10] ) );
  dp_1 \ANSWER/mem_reg[5][0][10]  ( .ip(n2852), .ck(clk), .q(
        \ANSWER/mem[5][0][10] ) );
  dp_1 \ANSWER/mem_reg[5][1][10]  ( .ip(n2851), .ck(clk), .q(
        \ANSWER/mem[5][1][10] ) );
  dp_1 \ANSWER/mem_reg[5][2][10]  ( .ip(n2850), .ck(clk), .q(
        \ANSWER/mem[5][2][10] ) );
  dp_1 \ANSWER/mem_reg[5][3][10]  ( .ip(n2849), .ck(clk), .q(
        \ANSWER/mem[5][3][10] ) );
  dp_1 \ANSWER/mem_reg[5][4][10]  ( .ip(n2848), .ck(clk), .q(
        \ANSWER/mem[5][4][10] ) );
  dp_1 \ANSWER/mem_reg[5][5][10]  ( .ip(n2847), .ck(clk), .q(
        \ANSWER/mem[5][5][10] ) );
  dp_1 \ANSWER/mem_reg[5][6][10]  ( .ip(n2846), .ck(clk), .q(
        \ANSWER/mem[5][6][10] ) );
  dp_1 \ANSWER/mem_reg[5][7][10]  ( .ip(n2845), .ck(clk), .q(
        \ANSWER/mem[5][7][10] ) );
  dp_1 \ANSWER/mem_reg[5][8][10]  ( .ip(n2844), .ck(clk), .q(
        \ANSWER/mem[5][8][10] ) );
  dp_1 \ANSWER/mem_reg[5][9][10]  ( .ip(n2843), .ck(clk), .q(
        \ANSWER/mem[5][9][10] ) );
  dp_1 \ANSWER/mem_reg[6][0][10]  ( .ip(n2842), .ck(clk), .q(
        \ANSWER/mem[6][0][10] ) );
  dp_1 \ANSWER/mem_reg[6][1][10]  ( .ip(n2841), .ck(clk), .q(
        \ANSWER/mem[6][1][10] ) );
  dp_1 \ANSWER/mem_reg[6][2][10]  ( .ip(n2840), .ck(clk), .q(
        \ANSWER/mem[6][2][10] ) );
  dp_1 \ANSWER/mem_reg[6][3][10]  ( .ip(n2839), .ck(clk), .q(
        \ANSWER/mem[6][3][10] ) );
  dp_1 \ANSWER/mem_reg[6][4][10]  ( .ip(n2838), .ck(clk), .q(
        \ANSWER/mem[6][4][10] ) );
  dp_1 \ANSWER/mem_reg[6][5][10]  ( .ip(n2837), .ck(clk), .q(
        \ANSWER/mem[6][5][10] ) );
  dp_1 \ANSWER/mem_reg[6][6][10]  ( .ip(n2836), .ck(clk), .q(
        \ANSWER/mem[6][6][10] ) );
  dp_1 \ANSWER/mem_reg[6][7][10]  ( .ip(n2835), .ck(clk), .q(
        \ANSWER/mem[6][7][10] ) );
  dp_1 \ANSWER/mem_reg[6][8][10]  ( .ip(n2834), .ck(clk), .q(
        \ANSWER/mem[6][8][10] ) );
  dp_1 \ANSWER/mem_reg[6][9][10]  ( .ip(n2833), .ck(clk), .q(
        \ANSWER/mem[6][9][10] ) );
  dp_1 \ANSWER/mem_reg[7][0][10]  ( .ip(n2832), .ck(clk), .q(
        \ANSWER/mem[7][0][10] ) );
  dp_1 \ANSWER/mem_reg[7][1][10]  ( .ip(n2831), .ck(clk), .q(
        \ANSWER/mem[7][1][10] ) );
  dp_1 \ANSWER/mem_reg[7][2][10]  ( .ip(n2830), .ck(clk), .q(
        \ANSWER/mem[7][2][10] ) );
  dp_1 \ANSWER/mem_reg[7][3][10]  ( .ip(n2829), .ck(clk), .q(
        \ANSWER/mem[7][3][10] ) );
  dp_1 \ANSWER/mem_reg[7][4][10]  ( .ip(n2828), .ck(clk), .q(
        \ANSWER/mem[7][4][10] ) );
  dp_1 \ANSWER/mem_reg[7][5][10]  ( .ip(n2827), .ck(clk), .q(
        \ANSWER/mem[7][5][10] ) );
  dp_1 \ANSWER/mem_reg[7][6][10]  ( .ip(n2826), .ck(clk), .q(
        \ANSWER/mem[7][6][10] ) );
  dp_1 \ANSWER/mem_reg[7][7][10]  ( .ip(n2825), .ck(clk), .q(
        \ANSWER/mem[7][7][10] ) );
  dp_1 \ANSWER/mem_reg[7][8][10]  ( .ip(n2824), .ck(clk), .q(
        \ANSWER/mem[7][8][10] ) );
  dp_1 \ANSWER/mem_reg[7][9][10]  ( .ip(n2823), .ck(clk), .q(
        \ANSWER/mem[7][9][10] ) );
  dp_1 \ANSWER/mem_reg[8][0][10]  ( .ip(n2822), .ck(clk), .q(
        \ANSWER/mem[8][0][10] ) );
  dp_1 \ANSWER/mem_reg[8][1][10]  ( .ip(n2821), .ck(clk), .q(
        \ANSWER/mem[8][1][10] ) );
  dp_1 \ANSWER/mem_reg[8][2][10]  ( .ip(n2820), .ck(clk), .q(
        \ANSWER/mem[8][2][10] ) );
  dp_1 \ANSWER/mem_reg[8][3][10]  ( .ip(n2819), .ck(clk), .q(
        \ANSWER/mem[8][3][10] ) );
  dp_1 \ANSWER/mem_reg[8][4][10]  ( .ip(n2818), .ck(clk), .q(
        \ANSWER/mem[8][4][10] ) );
  dp_1 \ANSWER/mem_reg[8][5][10]  ( .ip(n2817), .ck(clk), .q(
        \ANSWER/mem[8][5][10] ) );
  dp_1 \ANSWER/mem_reg[8][6][10]  ( .ip(n2816), .ck(clk), .q(
        \ANSWER/mem[8][6][10] ) );
  dp_1 \ANSWER/mem_reg[8][7][10]  ( .ip(n2815), .ck(clk), .q(
        \ANSWER/mem[8][7][10] ) );
  dp_1 \ANSWER/mem_reg[8][8][10]  ( .ip(n2814), .ck(clk), .q(
        \ANSWER/mem[8][8][10] ) );
  dp_1 \ANSWER/mem_reg[8][9][10]  ( .ip(n2813), .ck(clk), .q(
        \ANSWER/mem[8][9][10] ) );
  dp_1 \ANSWER/mem_reg[9][0][10]  ( .ip(n2812), .ck(clk), .q(
        \ANSWER/mem[9][0][10] ) );
  dp_1 \ANSWER/mem_reg[9][1][10]  ( .ip(n2811), .ck(clk), .q(
        \ANSWER/mem[9][1][10] ) );
  dp_1 \ANSWER/mem_reg[9][2][10]  ( .ip(n2810), .ck(clk), .q(
        \ANSWER/mem[9][2][10] ) );
  dp_1 \ANSWER/mem_reg[9][3][10]  ( .ip(n2809), .ck(clk), .q(
        \ANSWER/mem[9][3][10] ) );
  dp_1 \ANSWER/mem_reg[9][4][10]  ( .ip(n2808), .ck(clk), .q(
        \ANSWER/mem[9][4][10] ) );
  dp_1 \ANSWER/mem_reg[9][5][10]  ( .ip(n2807), .ck(clk), .q(
        \ANSWER/mem[9][5][10] ) );
  dp_1 \ANSWER/mem_reg[9][6][10]  ( .ip(n2806), .ck(clk), .q(
        \ANSWER/mem[9][6][10] ) );
  dp_1 \ANSWER/mem_reg[9][7][10]  ( .ip(n2805), .ck(clk), .q(
        \ANSWER/mem[9][7][10] ) );
  dp_1 \ANSWER/mem_reg[9][8][10]  ( .ip(n2804), .ck(clk), .q(
        \ANSWER/mem[9][8][10] ) );
  dp_1 \ANSWER/mem_reg[9][9][10]  ( .ip(n2803), .ck(clk), .q(
        \ANSWER/mem[9][9][10] ) );
  dp_1 \ANSWER/mem_reg[0][0][11]  ( .ip(n2802), .ck(clk), .q(
        \ANSWER/mem[0][0][11] ) );
  dp_1 \ANSWER/mem_reg[0][1][11]  ( .ip(n2801), .ck(clk), .q(
        \ANSWER/mem[0][1][11] ) );
  dp_1 \ANSWER/mem_reg[0][2][11]  ( .ip(n2800), .ck(clk), .q(
        \ANSWER/mem[0][2][11] ) );
  dp_1 \ANSWER/mem_reg[0][3][11]  ( .ip(n2799), .ck(clk), .q(
        \ANSWER/mem[0][3][11] ) );
  dp_1 \ANSWER/mem_reg[0][4][11]  ( .ip(n2798), .ck(clk), .q(
        \ANSWER/mem[0][4][11] ) );
  dp_1 \ANSWER/mem_reg[0][5][11]  ( .ip(n2797), .ck(clk), .q(
        \ANSWER/mem[0][5][11] ) );
  dp_1 \ANSWER/mem_reg[0][6][11]  ( .ip(n2796), .ck(clk), .q(
        \ANSWER/mem[0][6][11] ) );
  dp_1 \ANSWER/mem_reg[0][7][11]  ( .ip(n2795), .ck(clk), .q(
        \ANSWER/mem[0][7][11] ) );
  dp_1 \ANSWER/mem_reg[0][8][11]  ( .ip(n2794), .ck(clk), .q(
        \ANSWER/mem[0][8][11] ) );
  dp_1 \ANSWER/mem_reg[0][9][11]  ( .ip(n2793), .ck(clk), .q(
        \ANSWER/mem[0][9][11] ) );
  dp_1 \ANSWER/mem_reg[1][0][11]  ( .ip(n2792), .ck(clk), .q(
        \ANSWER/mem[1][0][11] ) );
  dp_1 \ANSWER/mem_reg[1][1][11]  ( .ip(n2791), .ck(clk), .q(
        \ANSWER/mem[1][1][11] ) );
  dp_1 \ANSWER/mem_reg[1][2][11]  ( .ip(n2790), .ck(clk), .q(
        \ANSWER/mem[1][2][11] ) );
  dp_1 \ANSWER/mem_reg[1][3][11]  ( .ip(n2789), .ck(clk), .q(
        \ANSWER/mem[1][3][11] ) );
  dp_1 \ANSWER/mem_reg[1][4][11]  ( .ip(n2788), .ck(clk), .q(
        \ANSWER/mem[1][4][11] ) );
  dp_1 \ANSWER/mem_reg[1][5][11]  ( .ip(n2787), .ck(clk), .q(
        \ANSWER/mem[1][5][11] ) );
  dp_1 \ANSWER/mem_reg[1][6][11]  ( .ip(n2786), .ck(clk), .q(
        \ANSWER/mem[1][6][11] ) );
  dp_1 \ANSWER/mem_reg[1][7][11]  ( .ip(n2785), .ck(clk), .q(
        \ANSWER/mem[1][7][11] ) );
  dp_1 \ANSWER/mem_reg[1][8][11]  ( .ip(n2784), .ck(clk), .q(
        \ANSWER/mem[1][8][11] ) );
  dp_1 \ANSWER/mem_reg[1][9][11]  ( .ip(n2783), .ck(clk), .q(
        \ANSWER/mem[1][9][11] ) );
  dp_1 \ANSWER/mem_reg[2][0][11]  ( .ip(n2782), .ck(clk), .q(
        \ANSWER/mem[2][0][11] ) );
  dp_1 \ANSWER/mem_reg[2][1][11]  ( .ip(n2781), .ck(clk), .q(
        \ANSWER/mem[2][1][11] ) );
  dp_1 \ANSWER/mem_reg[2][2][11]  ( .ip(n2780), .ck(clk), .q(
        \ANSWER/mem[2][2][11] ) );
  dp_1 \ANSWER/mem_reg[2][3][11]  ( .ip(n2779), .ck(clk), .q(
        \ANSWER/mem[2][3][11] ) );
  dp_1 \ANSWER/mem_reg[2][4][11]  ( .ip(n2778), .ck(clk), .q(
        \ANSWER/mem[2][4][11] ) );
  dp_1 \ANSWER/mem_reg[2][5][11]  ( .ip(n2777), .ck(clk), .q(
        \ANSWER/mem[2][5][11] ) );
  dp_1 \ANSWER/mem_reg[2][6][11]  ( .ip(n2776), .ck(clk), .q(
        \ANSWER/mem[2][6][11] ) );
  dp_1 \ANSWER/mem_reg[2][7][11]  ( .ip(n2775), .ck(clk), .q(
        \ANSWER/mem[2][7][11] ) );
  dp_1 \ANSWER/mem_reg[2][8][11]  ( .ip(n2774), .ck(clk), .q(
        \ANSWER/mem[2][8][11] ) );
  dp_1 \ANSWER/mem_reg[2][9][11]  ( .ip(n2773), .ck(clk), .q(
        \ANSWER/mem[2][9][11] ) );
  dp_1 \ANSWER/mem_reg[3][0][11]  ( .ip(n2772), .ck(clk), .q(
        \ANSWER/mem[3][0][11] ) );
  dp_1 \ANSWER/mem_reg[3][1][11]  ( .ip(n2771), .ck(clk), .q(
        \ANSWER/mem[3][1][11] ) );
  dp_1 \ANSWER/mem_reg[3][2][11]  ( .ip(n2770), .ck(clk), .q(
        \ANSWER/mem[3][2][11] ) );
  dp_1 \ANSWER/mem_reg[3][3][11]  ( .ip(n2769), .ck(clk), .q(
        \ANSWER/mem[3][3][11] ) );
  dp_1 \ANSWER/mem_reg[3][4][11]  ( .ip(n2768), .ck(clk), .q(
        \ANSWER/mem[3][4][11] ) );
  dp_1 \ANSWER/mem_reg[3][5][11]  ( .ip(n2767), .ck(clk), .q(
        \ANSWER/mem[3][5][11] ) );
  dp_1 \ANSWER/mem_reg[3][6][11]  ( .ip(n2766), .ck(clk), .q(
        \ANSWER/mem[3][6][11] ) );
  dp_1 \ANSWER/mem_reg[3][7][11]  ( .ip(n2765), .ck(clk), .q(
        \ANSWER/mem[3][7][11] ) );
  dp_1 \ANSWER/mem_reg[3][8][11]  ( .ip(n2764), .ck(clk), .q(
        \ANSWER/mem[3][8][11] ) );
  dp_1 \ANSWER/mem_reg[3][9][11]  ( .ip(n2763), .ck(clk), .q(
        \ANSWER/mem[3][9][11] ) );
  dp_1 \ANSWER/mem_reg[4][0][11]  ( .ip(n2762), .ck(clk), .q(
        \ANSWER/mem[4][0][11] ) );
  dp_1 \ANSWER/mem_reg[4][1][11]  ( .ip(n2761), .ck(clk), .q(
        \ANSWER/mem[4][1][11] ) );
  dp_1 \ANSWER/mem_reg[4][2][11]  ( .ip(n2760), .ck(clk), .q(
        \ANSWER/mem[4][2][11] ) );
  dp_1 \ANSWER/mem_reg[4][3][11]  ( .ip(n2759), .ck(clk), .q(
        \ANSWER/mem[4][3][11] ) );
  dp_1 \ANSWER/mem_reg[4][4][11]  ( .ip(n2758), .ck(clk), .q(
        \ANSWER/mem[4][4][11] ) );
  dp_1 \ANSWER/mem_reg[4][5][11]  ( .ip(n2757), .ck(clk), .q(
        \ANSWER/mem[4][5][11] ) );
  dp_1 \ANSWER/mem_reg[4][6][11]  ( .ip(n2756), .ck(clk), .q(
        \ANSWER/mem[4][6][11] ) );
  dp_1 \ANSWER/mem_reg[4][7][11]  ( .ip(n2755), .ck(clk), .q(
        \ANSWER/mem[4][7][11] ) );
  dp_1 \ANSWER/mem_reg[4][8][11]  ( .ip(n2754), .ck(clk), .q(
        \ANSWER/mem[4][8][11] ) );
  dp_1 \ANSWER/mem_reg[4][9][11]  ( .ip(n2753), .ck(clk), .q(
        \ANSWER/mem[4][9][11] ) );
  dp_1 \ANSWER/mem_reg[5][0][11]  ( .ip(n2752), .ck(clk), .q(
        \ANSWER/mem[5][0][11] ) );
  dp_1 \ANSWER/mem_reg[5][1][11]  ( .ip(n2751), .ck(clk), .q(
        \ANSWER/mem[5][1][11] ) );
  dp_1 \ANSWER/mem_reg[5][2][11]  ( .ip(n2750), .ck(clk), .q(
        \ANSWER/mem[5][2][11] ) );
  dp_1 \ANSWER/mem_reg[5][3][11]  ( .ip(n2749), .ck(clk), .q(
        \ANSWER/mem[5][3][11] ) );
  dp_1 \ANSWER/mem_reg[5][4][11]  ( .ip(n2748), .ck(clk), .q(
        \ANSWER/mem[5][4][11] ) );
  dp_1 \ANSWER/mem_reg[5][5][11]  ( .ip(n2747), .ck(clk), .q(
        \ANSWER/mem[5][5][11] ) );
  dp_1 \ANSWER/mem_reg[5][6][11]  ( .ip(n2746), .ck(clk), .q(
        \ANSWER/mem[5][6][11] ) );
  dp_1 \ANSWER/mem_reg[5][7][11]  ( .ip(n2745), .ck(clk), .q(
        \ANSWER/mem[5][7][11] ) );
  dp_1 \ANSWER/mem_reg[5][8][11]  ( .ip(n2744), .ck(clk), .q(
        \ANSWER/mem[5][8][11] ) );
  dp_1 \ANSWER/mem_reg[5][9][11]  ( .ip(n2743), .ck(clk), .q(
        \ANSWER/mem[5][9][11] ) );
  dp_1 \ANSWER/mem_reg[6][0][11]  ( .ip(n2742), .ck(clk), .q(
        \ANSWER/mem[6][0][11] ) );
  dp_1 \ANSWER/mem_reg[6][1][11]  ( .ip(n2741), .ck(clk), .q(
        \ANSWER/mem[6][1][11] ) );
  dp_1 \ANSWER/mem_reg[6][2][11]  ( .ip(n2740), .ck(clk), .q(
        \ANSWER/mem[6][2][11] ) );
  dp_1 \ANSWER/mem_reg[6][3][11]  ( .ip(n2739), .ck(clk), .q(
        \ANSWER/mem[6][3][11] ) );
  dp_1 \ANSWER/mem_reg[6][4][11]  ( .ip(n2738), .ck(clk), .q(
        \ANSWER/mem[6][4][11] ) );
  dp_1 \ANSWER/mem_reg[6][5][11]  ( .ip(n2737), .ck(clk), .q(
        \ANSWER/mem[6][5][11] ) );
  dp_1 \ANSWER/mem_reg[6][6][11]  ( .ip(n2736), .ck(clk), .q(
        \ANSWER/mem[6][6][11] ) );
  dp_1 \ANSWER/mem_reg[6][7][11]  ( .ip(n2735), .ck(clk), .q(
        \ANSWER/mem[6][7][11] ) );
  dp_1 \ANSWER/mem_reg[6][8][11]  ( .ip(n2734), .ck(clk), .q(
        \ANSWER/mem[6][8][11] ) );
  dp_1 \ANSWER/mem_reg[6][9][11]  ( .ip(n2733), .ck(clk), .q(
        \ANSWER/mem[6][9][11] ) );
  dp_1 \ANSWER/mem_reg[7][0][11]  ( .ip(n2732), .ck(clk), .q(
        \ANSWER/mem[7][0][11] ) );
  dp_1 \ANSWER/mem_reg[7][1][11]  ( .ip(n2731), .ck(clk), .q(
        \ANSWER/mem[7][1][11] ) );
  dp_1 \ANSWER/mem_reg[7][2][11]  ( .ip(n2730), .ck(clk), .q(
        \ANSWER/mem[7][2][11] ) );
  dp_1 \ANSWER/mem_reg[7][3][11]  ( .ip(n2729), .ck(clk), .q(
        \ANSWER/mem[7][3][11] ) );
  dp_1 \ANSWER/mem_reg[7][4][11]  ( .ip(n2728), .ck(clk), .q(
        \ANSWER/mem[7][4][11] ) );
  dp_1 \ANSWER/mem_reg[7][5][11]  ( .ip(n2727), .ck(clk), .q(
        \ANSWER/mem[7][5][11] ) );
  dp_1 \ANSWER/mem_reg[7][6][11]  ( .ip(n2726), .ck(clk), .q(
        \ANSWER/mem[7][6][11] ) );
  dp_1 \ANSWER/mem_reg[7][7][11]  ( .ip(n2725), .ck(clk), .q(
        \ANSWER/mem[7][7][11] ) );
  dp_1 \ANSWER/mem_reg[7][8][11]  ( .ip(n2724), .ck(clk), .q(
        \ANSWER/mem[7][8][11] ) );
  dp_1 \ANSWER/mem_reg[7][9][11]  ( .ip(n2723), .ck(clk), .q(
        \ANSWER/mem[7][9][11] ) );
  dp_1 \ANSWER/mem_reg[8][0][11]  ( .ip(n2722), .ck(clk), .q(
        \ANSWER/mem[8][0][11] ) );
  dp_1 \ANSWER/mem_reg[8][1][11]  ( .ip(n2721), .ck(clk), .q(
        \ANSWER/mem[8][1][11] ) );
  dp_1 \ANSWER/mem_reg[8][2][11]  ( .ip(n2720), .ck(clk), .q(
        \ANSWER/mem[8][2][11] ) );
  dp_1 \ANSWER/mem_reg[8][3][11]  ( .ip(n2719), .ck(clk), .q(
        \ANSWER/mem[8][3][11] ) );
  dp_1 \ANSWER/mem_reg[8][4][11]  ( .ip(n2718), .ck(clk), .q(
        \ANSWER/mem[8][4][11] ) );
  dp_1 \ANSWER/mem_reg[8][5][11]  ( .ip(n2717), .ck(clk), .q(
        \ANSWER/mem[8][5][11] ) );
  dp_1 \ANSWER/mem_reg[8][6][11]  ( .ip(n2716), .ck(clk), .q(
        \ANSWER/mem[8][6][11] ) );
  dp_1 \ANSWER/mem_reg[8][7][11]  ( .ip(n2715), .ck(clk), .q(
        \ANSWER/mem[8][7][11] ) );
  dp_1 \ANSWER/mem_reg[8][8][11]  ( .ip(n2714), .ck(clk), .q(
        \ANSWER/mem[8][8][11] ) );
  dp_1 \ANSWER/mem_reg[8][9][11]  ( .ip(n2713), .ck(clk), .q(
        \ANSWER/mem[8][9][11] ) );
  dp_1 \ANSWER/mem_reg[9][0][11]  ( .ip(n2712), .ck(clk), .q(
        \ANSWER/mem[9][0][11] ) );
  dp_1 \ANSWER/mem_reg[9][1][11]  ( .ip(n2711), .ck(clk), .q(
        \ANSWER/mem[9][1][11] ) );
  dp_1 \ANSWER/mem_reg[9][2][11]  ( .ip(n2710), .ck(clk), .q(
        \ANSWER/mem[9][2][11] ) );
  dp_1 \ANSWER/mem_reg[9][3][11]  ( .ip(n2709), .ck(clk), .q(
        \ANSWER/mem[9][3][11] ) );
  dp_1 \ANSWER/mem_reg[9][4][11]  ( .ip(n2708), .ck(clk), .q(
        \ANSWER/mem[9][4][11] ) );
  dp_1 \ANSWER/mem_reg[9][5][11]  ( .ip(n2707), .ck(clk), .q(
        \ANSWER/mem[9][5][11] ) );
  dp_1 \ANSWER/mem_reg[9][6][11]  ( .ip(n2706), .ck(clk), .q(
        \ANSWER/mem[9][6][11] ) );
  dp_1 \ANSWER/mem_reg[9][7][11]  ( .ip(n2705), .ck(clk), .q(
        \ANSWER/mem[9][7][11] ) );
  dp_1 \ANSWER/mem_reg[9][8][11]  ( .ip(n2704), .ck(clk), .q(
        \ANSWER/mem[9][8][11] ) );
  dp_1 \ANSWER/mem_reg[9][9][11]  ( .ip(n2703), .ck(clk), .q(
        \ANSWER/mem[9][9][11] ) );
  dp_1 \ANSWER/mem_reg[0][0][12]  ( .ip(n2702), .ck(clk), .q(
        \ANSWER/mem[0][0][12] ) );
  dp_1 \ANSWER/mem_reg[0][1][12]  ( .ip(n2701), .ck(clk), .q(
        \ANSWER/mem[0][1][12] ) );
  dp_1 \ANSWER/mem_reg[0][2][12]  ( .ip(n2700), .ck(clk), .q(
        \ANSWER/mem[0][2][12] ) );
  dp_1 \ANSWER/mem_reg[0][3][12]  ( .ip(n2699), .ck(clk), .q(
        \ANSWER/mem[0][3][12] ) );
  dp_1 \ANSWER/mem_reg[0][4][12]  ( .ip(n2698), .ck(clk), .q(
        \ANSWER/mem[0][4][12] ) );
  dp_1 \ANSWER/mem_reg[0][5][12]  ( .ip(n2697), .ck(clk), .q(
        \ANSWER/mem[0][5][12] ) );
  dp_1 \ANSWER/mem_reg[0][6][12]  ( .ip(n2696), .ck(clk), .q(
        \ANSWER/mem[0][6][12] ) );
  dp_1 \ANSWER/mem_reg[0][7][12]  ( .ip(n2695), .ck(clk), .q(
        \ANSWER/mem[0][7][12] ) );
  dp_1 \ANSWER/mem_reg[0][8][12]  ( .ip(n2694), .ck(clk), .q(
        \ANSWER/mem[0][8][12] ) );
  dp_1 \ANSWER/mem_reg[0][9][12]  ( .ip(n2693), .ck(clk), .q(
        \ANSWER/mem[0][9][12] ) );
  dp_1 \ANSWER/mem_reg[1][0][12]  ( .ip(n2692), .ck(clk), .q(
        \ANSWER/mem[1][0][12] ) );
  dp_1 \ANSWER/mem_reg[1][1][12]  ( .ip(n2691), .ck(clk), .q(
        \ANSWER/mem[1][1][12] ) );
  dp_1 \ANSWER/mem_reg[1][2][12]  ( .ip(n2690), .ck(clk), .q(
        \ANSWER/mem[1][2][12] ) );
  dp_1 \ANSWER/mem_reg[1][3][12]  ( .ip(n2689), .ck(clk), .q(
        \ANSWER/mem[1][3][12] ) );
  dp_1 \ANSWER/mem_reg[1][4][12]  ( .ip(n2688), .ck(clk), .q(
        \ANSWER/mem[1][4][12] ) );
  dp_1 \ANSWER/mem_reg[1][5][12]  ( .ip(n2687), .ck(clk), .q(
        \ANSWER/mem[1][5][12] ) );
  dp_1 \ANSWER/mem_reg[1][6][12]  ( .ip(n2686), .ck(clk), .q(
        \ANSWER/mem[1][6][12] ) );
  dp_1 \ANSWER/mem_reg[1][7][12]  ( .ip(n2685), .ck(clk), .q(
        \ANSWER/mem[1][7][12] ) );
  dp_1 \ANSWER/mem_reg[1][8][12]  ( .ip(n2684), .ck(clk), .q(
        \ANSWER/mem[1][8][12] ) );
  dp_1 \ANSWER/mem_reg[1][9][12]  ( .ip(n2683), .ck(clk), .q(
        \ANSWER/mem[1][9][12] ) );
  dp_1 \ANSWER/mem_reg[2][0][12]  ( .ip(n2682), .ck(clk), .q(
        \ANSWER/mem[2][0][12] ) );
  dp_1 \ANSWER/mem_reg[2][1][12]  ( .ip(n2681), .ck(clk), .q(
        \ANSWER/mem[2][1][12] ) );
  dp_1 \ANSWER/mem_reg[2][2][12]  ( .ip(n2680), .ck(clk), .q(
        \ANSWER/mem[2][2][12] ) );
  dp_1 \ANSWER/mem_reg[2][3][12]  ( .ip(n2679), .ck(clk), .q(
        \ANSWER/mem[2][3][12] ) );
  dp_1 \ANSWER/mem_reg[2][4][12]  ( .ip(n2678), .ck(clk), .q(
        \ANSWER/mem[2][4][12] ) );
  dp_1 \ANSWER/mem_reg[2][5][12]  ( .ip(n2677), .ck(clk), .q(
        \ANSWER/mem[2][5][12] ) );
  dp_1 \ANSWER/mem_reg[2][6][12]  ( .ip(n2676), .ck(clk), .q(
        \ANSWER/mem[2][6][12] ) );
  dp_1 \ANSWER/mem_reg[2][7][12]  ( .ip(n2675), .ck(clk), .q(
        \ANSWER/mem[2][7][12] ) );
  dp_1 \ANSWER/mem_reg[2][8][12]  ( .ip(n2674), .ck(clk), .q(
        \ANSWER/mem[2][8][12] ) );
  dp_1 \ANSWER/mem_reg[2][9][12]  ( .ip(n2673), .ck(clk), .q(
        \ANSWER/mem[2][9][12] ) );
  dp_1 \ANSWER/mem_reg[3][0][12]  ( .ip(n2672), .ck(clk), .q(
        \ANSWER/mem[3][0][12] ) );
  dp_1 \ANSWER/mem_reg[3][1][12]  ( .ip(n2671), .ck(clk), .q(
        \ANSWER/mem[3][1][12] ) );
  dp_1 \ANSWER/mem_reg[3][2][12]  ( .ip(n2670), .ck(clk), .q(
        \ANSWER/mem[3][2][12] ) );
  dp_1 \ANSWER/mem_reg[3][3][12]  ( .ip(n2669), .ck(clk), .q(
        \ANSWER/mem[3][3][12] ) );
  dp_1 \ANSWER/mem_reg[3][4][12]  ( .ip(n2668), .ck(clk), .q(
        \ANSWER/mem[3][4][12] ) );
  dp_1 \ANSWER/mem_reg[3][5][12]  ( .ip(n2667), .ck(clk), .q(
        \ANSWER/mem[3][5][12] ) );
  dp_1 \ANSWER/mem_reg[3][6][12]  ( .ip(n2666), .ck(clk), .q(
        \ANSWER/mem[3][6][12] ) );
  dp_1 \ANSWER/mem_reg[3][7][12]  ( .ip(n2665), .ck(clk), .q(
        \ANSWER/mem[3][7][12] ) );
  dp_1 \ANSWER/mem_reg[3][8][12]  ( .ip(n2664), .ck(clk), .q(
        \ANSWER/mem[3][8][12] ) );
  dp_1 \ANSWER/mem_reg[3][9][12]  ( .ip(n2663), .ck(clk), .q(
        \ANSWER/mem[3][9][12] ) );
  dp_1 \ANSWER/mem_reg[4][0][12]  ( .ip(n2662), .ck(clk), .q(
        \ANSWER/mem[4][0][12] ) );
  dp_1 \ANSWER/mem_reg[4][1][12]  ( .ip(n2661), .ck(clk), .q(
        \ANSWER/mem[4][1][12] ) );
  dp_1 \ANSWER/mem_reg[4][2][12]  ( .ip(n2660), .ck(clk), .q(
        \ANSWER/mem[4][2][12] ) );
  dp_1 \ANSWER/mem_reg[4][3][12]  ( .ip(n2659), .ck(clk), .q(
        \ANSWER/mem[4][3][12] ) );
  dp_1 \ANSWER/mem_reg[4][4][12]  ( .ip(n2658), .ck(clk), .q(
        \ANSWER/mem[4][4][12] ) );
  dp_1 \ANSWER/mem_reg[4][5][12]  ( .ip(n2657), .ck(clk), .q(
        \ANSWER/mem[4][5][12] ) );
  dp_1 \ANSWER/mem_reg[4][6][12]  ( .ip(n2656), .ck(clk), .q(
        \ANSWER/mem[4][6][12] ) );
  dp_1 \ANSWER/mem_reg[4][7][12]  ( .ip(n2655), .ck(clk), .q(
        \ANSWER/mem[4][7][12] ) );
  dp_1 \ANSWER/mem_reg[4][8][12]  ( .ip(n2654), .ck(clk), .q(
        \ANSWER/mem[4][8][12] ) );
  dp_1 \ANSWER/mem_reg[4][9][12]  ( .ip(n2653), .ck(clk), .q(
        \ANSWER/mem[4][9][12] ) );
  dp_1 \ANSWER/mem_reg[5][0][12]  ( .ip(n2652), .ck(clk), .q(
        \ANSWER/mem[5][0][12] ) );
  dp_1 \ANSWER/mem_reg[5][1][12]  ( .ip(n2651), .ck(clk), .q(
        \ANSWER/mem[5][1][12] ) );
  dp_1 \ANSWER/mem_reg[5][2][12]  ( .ip(n2650), .ck(clk), .q(
        \ANSWER/mem[5][2][12] ) );
  dp_1 \ANSWER/mem_reg[5][3][12]  ( .ip(n2649), .ck(clk), .q(
        \ANSWER/mem[5][3][12] ) );
  dp_1 \ANSWER/mem_reg[5][4][12]  ( .ip(n2648), .ck(clk), .q(
        \ANSWER/mem[5][4][12] ) );
  dp_1 \ANSWER/mem_reg[5][5][12]  ( .ip(n2647), .ck(clk), .q(
        \ANSWER/mem[5][5][12] ) );
  dp_1 \ANSWER/mem_reg[5][6][12]  ( .ip(n2646), .ck(clk), .q(
        \ANSWER/mem[5][6][12] ) );
  dp_1 \ANSWER/mem_reg[5][7][12]  ( .ip(n2645), .ck(clk), .q(
        \ANSWER/mem[5][7][12] ) );
  dp_1 \ANSWER/mem_reg[5][8][12]  ( .ip(n2644), .ck(clk), .q(
        \ANSWER/mem[5][8][12] ) );
  dp_1 \ANSWER/mem_reg[5][9][12]  ( .ip(n2643), .ck(clk), .q(
        \ANSWER/mem[5][9][12] ) );
  dp_1 \ANSWER/mem_reg[6][0][12]  ( .ip(n2642), .ck(clk), .q(
        \ANSWER/mem[6][0][12] ) );
  dp_1 \ANSWER/mem_reg[6][1][12]  ( .ip(n2641), .ck(clk), .q(
        \ANSWER/mem[6][1][12] ) );
  dp_1 \ANSWER/mem_reg[6][2][12]  ( .ip(n2640), .ck(clk), .q(
        \ANSWER/mem[6][2][12] ) );
  dp_1 \ANSWER/mem_reg[6][3][12]  ( .ip(n2639), .ck(clk), .q(
        \ANSWER/mem[6][3][12] ) );
  dp_1 \ANSWER/mem_reg[6][4][12]  ( .ip(n2638), .ck(clk), .q(
        \ANSWER/mem[6][4][12] ) );
  dp_1 \ANSWER/mem_reg[6][5][12]  ( .ip(n2637), .ck(clk), .q(
        \ANSWER/mem[6][5][12] ) );
  dp_1 \ANSWER/mem_reg[6][6][12]  ( .ip(n2636), .ck(clk), .q(
        \ANSWER/mem[6][6][12] ) );
  dp_1 \ANSWER/mem_reg[6][7][12]  ( .ip(n2635), .ck(clk), .q(
        \ANSWER/mem[6][7][12] ) );
  dp_1 \ANSWER/mem_reg[6][8][12]  ( .ip(n2634), .ck(clk), .q(
        \ANSWER/mem[6][8][12] ) );
  dp_1 \ANSWER/mem_reg[6][9][12]  ( .ip(n2633), .ck(clk), .q(
        \ANSWER/mem[6][9][12] ) );
  dp_1 \ANSWER/mem_reg[7][0][12]  ( .ip(n2632), .ck(clk), .q(
        \ANSWER/mem[7][0][12] ) );
  dp_1 \ANSWER/mem_reg[7][1][12]  ( .ip(n2631), .ck(clk), .q(
        \ANSWER/mem[7][1][12] ) );
  dp_1 \ANSWER/mem_reg[7][2][12]  ( .ip(n2630), .ck(clk), .q(
        \ANSWER/mem[7][2][12] ) );
  dp_1 \ANSWER/mem_reg[7][3][12]  ( .ip(n2629), .ck(clk), .q(
        \ANSWER/mem[7][3][12] ) );
  dp_1 \ANSWER/mem_reg[7][4][12]  ( .ip(n2628), .ck(clk), .q(
        \ANSWER/mem[7][4][12] ) );
  dp_1 \ANSWER/mem_reg[7][5][12]  ( .ip(n2627), .ck(clk), .q(
        \ANSWER/mem[7][5][12] ) );
  dp_1 \ANSWER/mem_reg[7][6][12]  ( .ip(n2626), .ck(clk), .q(
        \ANSWER/mem[7][6][12] ) );
  dp_1 \ANSWER/mem_reg[7][7][12]  ( .ip(n2625), .ck(clk), .q(
        \ANSWER/mem[7][7][12] ) );
  dp_1 \ANSWER/mem_reg[7][8][12]  ( .ip(n2624), .ck(clk), .q(
        \ANSWER/mem[7][8][12] ) );
  dp_1 \ANSWER/mem_reg[7][9][12]  ( .ip(n2623), .ck(clk), .q(
        \ANSWER/mem[7][9][12] ) );
  dp_1 \ANSWER/mem_reg[8][0][12]  ( .ip(n2622), .ck(clk), .q(
        \ANSWER/mem[8][0][12] ) );
  dp_1 \ANSWER/mem_reg[8][1][12]  ( .ip(n2621), .ck(clk), .q(
        \ANSWER/mem[8][1][12] ) );
  dp_1 \ANSWER/mem_reg[8][2][12]  ( .ip(n2620), .ck(clk), .q(
        \ANSWER/mem[8][2][12] ) );
  dp_1 \ANSWER/mem_reg[8][3][12]  ( .ip(n2619), .ck(clk), .q(
        \ANSWER/mem[8][3][12] ) );
  dp_1 \ANSWER/mem_reg[8][4][12]  ( .ip(n2618), .ck(clk), .q(
        \ANSWER/mem[8][4][12] ) );
  dp_1 \ANSWER/mem_reg[8][5][12]  ( .ip(n2617), .ck(clk), .q(
        \ANSWER/mem[8][5][12] ) );
  dp_1 \ANSWER/mem_reg[8][6][12]  ( .ip(n2616), .ck(clk), .q(
        \ANSWER/mem[8][6][12] ) );
  dp_1 \ANSWER/mem_reg[8][7][12]  ( .ip(n2615), .ck(clk), .q(
        \ANSWER/mem[8][7][12] ) );
  dp_1 \ANSWER/mem_reg[8][8][12]  ( .ip(n2614), .ck(clk), .q(
        \ANSWER/mem[8][8][12] ) );
  dp_1 \ANSWER/mem_reg[8][9][12]  ( .ip(n2613), .ck(clk), .q(
        \ANSWER/mem[8][9][12] ) );
  dp_1 \ANSWER/mem_reg[9][0][12]  ( .ip(n2612), .ck(clk), .q(
        \ANSWER/mem[9][0][12] ) );
  dp_1 \ANSWER/mem_reg[9][1][12]  ( .ip(n2611), .ck(clk), .q(
        \ANSWER/mem[9][1][12] ) );
  dp_1 \ANSWER/mem_reg[9][2][12]  ( .ip(n2610), .ck(clk), .q(
        \ANSWER/mem[9][2][12] ) );
  dp_1 \ANSWER/mem_reg[9][3][12]  ( .ip(n2609), .ck(clk), .q(
        \ANSWER/mem[9][3][12] ) );
  dp_1 \ANSWER/mem_reg[9][4][12]  ( .ip(n2608), .ck(clk), .q(
        \ANSWER/mem[9][4][12] ) );
  dp_1 \ANSWER/mem_reg[9][5][12]  ( .ip(n2607), .ck(clk), .q(
        \ANSWER/mem[9][5][12] ) );
  dp_1 \ANSWER/mem_reg[9][6][12]  ( .ip(n2606), .ck(clk), .q(
        \ANSWER/mem[9][6][12] ) );
  dp_1 \ANSWER/mem_reg[9][7][12]  ( .ip(n2605), .ck(clk), .q(
        \ANSWER/mem[9][7][12] ) );
  dp_1 \ANSWER/mem_reg[9][8][12]  ( .ip(n2604), .ck(clk), .q(
        \ANSWER/mem[9][8][12] ) );
  dp_1 \ANSWER/mem_reg[9][9][12]  ( .ip(n2603), .ck(clk), .q(
        \ANSWER/mem[9][9][12] ) );
  dp_1 \ANSWER/mem_reg[0][0][13]  ( .ip(n2602), .ck(clk), .q(
        \ANSWER/mem[0][0][13] ) );
  dp_1 \ANSWER/mem_reg[0][1][13]  ( .ip(n2601), .ck(clk), .q(
        \ANSWER/mem[0][1][13] ) );
  dp_1 \ANSWER/mem_reg[0][2][13]  ( .ip(n2600), .ck(clk), .q(
        \ANSWER/mem[0][2][13] ) );
  dp_1 \ANSWER/mem_reg[0][3][13]  ( .ip(n2599), .ck(clk), .q(
        \ANSWER/mem[0][3][13] ) );
  dp_1 \ANSWER/mem_reg[0][4][13]  ( .ip(n2598), .ck(clk), .q(
        \ANSWER/mem[0][4][13] ) );
  dp_1 \ANSWER/mem_reg[0][5][13]  ( .ip(n2597), .ck(clk), .q(
        \ANSWER/mem[0][5][13] ) );
  dp_1 \ANSWER/mem_reg[0][6][13]  ( .ip(n2596), .ck(clk), .q(
        \ANSWER/mem[0][6][13] ) );
  dp_1 \ANSWER/mem_reg[0][7][13]  ( .ip(n2595), .ck(clk), .q(
        \ANSWER/mem[0][7][13] ) );
  dp_1 \ANSWER/mem_reg[0][8][13]  ( .ip(n2594), .ck(clk), .q(
        \ANSWER/mem[0][8][13] ) );
  dp_1 \ANSWER/mem_reg[0][9][13]  ( .ip(n2593), .ck(clk), .q(
        \ANSWER/mem[0][9][13] ) );
  dp_1 \ANSWER/mem_reg[1][0][13]  ( .ip(n2592), .ck(clk), .q(
        \ANSWER/mem[1][0][13] ) );
  dp_1 \ANSWER/mem_reg[1][1][13]  ( .ip(n2591), .ck(clk), .q(
        \ANSWER/mem[1][1][13] ) );
  dp_1 \ANSWER/mem_reg[1][2][13]  ( .ip(n2590), .ck(clk), .q(
        \ANSWER/mem[1][2][13] ) );
  dp_1 \ANSWER/mem_reg[1][3][13]  ( .ip(n2589), .ck(clk), .q(
        \ANSWER/mem[1][3][13] ) );
  dp_1 \ANSWER/mem_reg[1][4][13]  ( .ip(n2588), .ck(clk), .q(
        \ANSWER/mem[1][4][13] ) );
  dp_1 \ANSWER/mem_reg[1][5][13]  ( .ip(n2587), .ck(clk), .q(
        \ANSWER/mem[1][5][13] ) );
  dp_1 \ANSWER/mem_reg[1][6][13]  ( .ip(n2586), .ck(clk), .q(
        \ANSWER/mem[1][6][13] ) );
  dp_1 \ANSWER/mem_reg[1][7][13]  ( .ip(n2585), .ck(clk), .q(
        \ANSWER/mem[1][7][13] ) );
  dp_1 \ANSWER/mem_reg[1][8][13]  ( .ip(n2584), .ck(clk), .q(
        \ANSWER/mem[1][8][13] ) );
  dp_1 \ANSWER/mem_reg[1][9][13]  ( .ip(n2583), .ck(clk), .q(
        \ANSWER/mem[1][9][13] ) );
  dp_1 \ANSWER/mem_reg[2][0][13]  ( .ip(n2582), .ck(clk), .q(
        \ANSWER/mem[2][0][13] ) );
  dp_1 \ANSWER/mem_reg[2][1][13]  ( .ip(n2581), .ck(clk), .q(
        \ANSWER/mem[2][1][13] ) );
  dp_1 \ANSWER/mem_reg[2][2][13]  ( .ip(n2580), .ck(clk), .q(
        \ANSWER/mem[2][2][13] ) );
  dp_1 \ANSWER/mem_reg[2][3][13]  ( .ip(n2579), .ck(clk), .q(
        \ANSWER/mem[2][3][13] ) );
  dp_1 \ANSWER/mem_reg[2][4][13]  ( .ip(n2578), .ck(clk), .q(
        \ANSWER/mem[2][4][13] ) );
  dp_1 \ANSWER/mem_reg[2][5][13]  ( .ip(n2577), .ck(clk), .q(
        \ANSWER/mem[2][5][13] ) );
  dp_1 \ANSWER/mem_reg[2][6][13]  ( .ip(n2576), .ck(clk), .q(
        \ANSWER/mem[2][6][13] ) );
  dp_1 \ANSWER/mem_reg[2][7][13]  ( .ip(n2575), .ck(clk), .q(
        \ANSWER/mem[2][7][13] ) );
  dp_1 \ANSWER/mem_reg[2][8][13]  ( .ip(n2574), .ck(clk), .q(
        \ANSWER/mem[2][8][13] ) );
  dp_1 \ANSWER/mem_reg[2][9][13]  ( .ip(n2573), .ck(clk), .q(
        \ANSWER/mem[2][9][13] ) );
  dp_1 \ANSWER/mem_reg[3][0][13]  ( .ip(n2572), .ck(clk), .q(
        \ANSWER/mem[3][0][13] ) );
  dp_1 \ANSWER/mem_reg[3][1][13]  ( .ip(n2571), .ck(clk), .q(
        \ANSWER/mem[3][1][13] ) );
  dp_1 \ANSWER/mem_reg[3][2][13]  ( .ip(n2570), .ck(clk), .q(
        \ANSWER/mem[3][2][13] ) );
  dp_1 \ANSWER/mem_reg[3][3][13]  ( .ip(n2569), .ck(clk), .q(
        \ANSWER/mem[3][3][13] ) );
  dp_1 \ANSWER/mem_reg[3][4][13]  ( .ip(n2568), .ck(clk), .q(
        \ANSWER/mem[3][4][13] ) );
  dp_1 \ANSWER/mem_reg[3][5][13]  ( .ip(n2567), .ck(clk), .q(
        \ANSWER/mem[3][5][13] ) );
  dp_1 \ANSWER/mem_reg[3][6][13]  ( .ip(n2566), .ck(clk), .q(
        \ANSWER/mem[3][6][13] ) );
  dp_1 \ANSWER/mem_reg[3][7][13]  ( .ip(n2565), .ck(clk), .q(
        \ANSWER/mem[3][7][13] ) );
  dp_1 \ANSWER/mem_reg[3][8][13]  ( .ip(n2564), .ck(clk), .q(
        \ANSWER/mem[3][8][13] ) );
  dp_1 \ANSWER/mem_reg[3][9][13]  ( .ip(n2563), .ck(clk), .q(
        \ANSWER/mem[3][9][13] ) );
  dp_1 \ANSWER/mem_reg[4][0][13]  ( .ip(n2562), .ck(clk), .q(
        \ANSWER/mem[4][0][13] ) );
  dp_1 \ANSWER/mem_reg[4][1][13]  ( .ip(n2561), .ck(clk), .q(
        \ANSWER/mem[4][1][13] ) );
  dp_1 \ANSWER/mem_reg[4][2][13]  ( .ip(n2560), .ck(clk), .q(
        \ANSWER/mem[4][2][13] ) );
  dp_1 \ANSWER/mem_reg[4][3][13]  ( .ip(n2559), .ck(clk), .q(
        \ANSWER/mem[4][3][13] ) );
  dp_1 \ANSWER/mem_reg[4][4][13]  ( .ip(n2558), .ck(clk), .q(
        \ANSWER/mem[4][4][13] ) );
  dp_1 \ANSWER/mem_reg[4][5][13]  ( .ip(n2557), .ck(clk), .q(
        \ANSWER/mem[4][5][13] ) );
  dp_1 \ANSWER/mem_reg[4][6][13]  ( .ip(n2556), .ck(clk), .q(
        \ANSWER/mem[4][6][13] ) );
  dp_1 \ANSWER/mem_reg[4][7][13]  ( .ip(n2555), .ck(clk), .q(
        \ANSWER/mem[4][7][13] ) );
  dp_1 \ANSWER/mem_reg[4][8][13]  ( .ip(n2554), .ck(clk), .q(
        \ANSWER/mem[4][8][13] ) );
  dp_1 \ANSWER/mem_reg[4][9][13]  ( .ip(n2553), .ck(clk), .q(
        \ANSWER/mem[4][9][13] ) );
  dp_1 \ANSWER/mem_reg[5][0][13]  ( .ip(n2552), .ck(clk), .q(
        \ANSWER/mem[5][0][13] ) );
  dp_1 \ANSWER/mem_reg[5][1][13]  ( .ip(n2551), .ck(clk), .q(
        \ANSWER/mem[5][1][13] ) );
  dp_1 \ANSWER/mem_reg[5][2][13]  ( .ip(n2550), .ck(clk), .q(
        \ANSWER/mem[5][2][13] ) );
  dp_1 \ANSWER/mem_reg[5][3][13]  ( .ip(n2549), .ck(clk), .q(
        \ANSWER/mem[5][3][13] ) );
  dp_1 \ANSWER/mem_reg[5][4][13]  ( .ip(n2548), .ck(clk), .q(
        \ANSWER/mem[5][4][13] ) );
  dp_1 \ANSWER/mem_reg[5][5][13]  ( .ip(n2547), .ck(clk), .q(
        \ANSWER/mem[5][5][13] ) );
  dp_1 \ANSWER/mem_reg[5][6][13]  ( .ip(n2546), .ck(clk), .q(
        \ANSWER/mem[5][6][13] ) );
  dp_1 \ANSWER/mem_reg[5][7][13]  ( .ip(n2545), .ck(clk), .q(
        \ANSWER/mem[5][7][13] ) );
  dp_1 \ANSWER/mem_reg[5][8][13]  ( .ip(n2544), .ck(clk), .q(
        \ANSWER/mem[5][8][13] ) );
  dp_1 \ANSWER/mem_reg[5][9][13]  ( .ip(n2543), .ck(clk), .q(
        \ANSWER/mem[5][9][13] ) );
  dp_1 \ANSWER/mem_reg[6][0][13]  ( .ip(n2542), .ck(clk), .q(
        \ANSWER/mem[6][0][13] ) );
  dp_1 \ANSWER/mem_reg[6][1][13]  ( .ip(n2541), .ck(clk), .q(
        \ANSWER/mem[6][1][13] ) );
  dp_1 \ANSWER/mem_reg[6][2][13]  ( .ip(n2540), .ck(clk), .q(
        \ANSWER/mem[6][2][13] ) );
  dp_1 \ANSWER/mem_reg[6][3][13]  ( .ip(n2539), .ck(clk), .q(
        \ANSWER/mem[6][3][13] ) );
  dp_1 \ANSWER/mem_reg[6][4][13]  ( .ip(n2538), .ck(clk), .q(
        \ANSWER/mem[6][4][13] ) );
  dp_1 \ANSWER/mem_reg[6][5][13]  ( .ip(n2537), .ck(clk), .q(
        \ANSWER/mem[6][5][13] ) );
  dp_1 \ANSWER/mem_reg[6][6][13]  ( .ip(n2536), .ck(clk), .q(
        \ANSWER/mem[6][6][13] ) );
  dp_1 \ANSWER/mem_reg[6][7][13]  ( .ip(n2535), .ck(clk), .q(
        \ANSWER/mem[6][7][13] ) );
  dp_1 \ANSWER/mem_reg[6][8][13]  ( .ip(n2534), .ck(clk), .q(
        \ANSWER/mem[6][8][13] ) );
  dp_1 \ANSWER/mem_reg[6][9][13]  ( .ip(n2533), .ck(clk), .q(
        \ANSWER/mem[6][9][13] ) );
  dp_1 \ANSWER/mem_reg[7][0][13]  ( .ip(n2532), .ck(clk), .q(
        \ANSWER/mem[7][0][13] ) );
  dp_1 \ANSWER/mem_reg[7][1][13]  ( .ip(n2531), .ck(clk), .q(
        \ANSWER/mem[7][1][13] ) );
  dp_1 \ANSWER/mem_reg[7][2][13]  ( .ip(n2530), .ck(clk), .q(
        \ANSWER/mem[7][2][13] ) );
  dp_1 \ANSWER/mem_reg[7][3][13]  ( .ip(n2529), .ck(clk), .q(
        \ANSWER/mem[7][3][13] ) );
  dp_1 \ANSWER/mem_reg[7][4][13]  ( .ip(n2528), .ck(clk), .q(
        \ANSWER/mem[7][4][13] ) );
  dp_1 \ANSWER/mem_reg[7][5][13]  ( .ip(n2527), .ck(clk), .q(
        \ANSWER/mem[7][5][13] ) );
  dp_1 \ANSWER/mem_reg[7][6][13]  ( .ip(n2526), .ck(clk), .q(
        \ANSWER/mem[7][6][13] ) );
  dp_1 \ANSWER/mem_reg[7][7][13]  ( .ip(n2525), .ck(clk), .q(
        \ANSWER/mem[7][7][13] ) );
  dp_1 \ANSWER/mem_reg[7][8][13]  ( .ip(n2524), .ck(clk), .q(
        \ANSWER/mem[7][8][13] ) );
  dp_1 \ANSWER/mem_reg[7][9][13]  ( .ip(n2523), .ck(clk), .q(
        \ANSWER/mem[7][9][13] ) );
  dp_1 \ANSWER/mem_reg[8][0][13]  ( .ip(n2522), .ck(clk), .q(
        \ANSWER/mem[8][0][13] ) );
  dp_1 \ANSWER/mem_reg[8][1][13]  ( .ip(n2521), .ck(clk), .q(
        \ANSWER/mem[8][1][13] ) );
  dp_1 \ANSWER/mem_reg[8][2][13]  ( .ip(n2520), .ck(clk), .q(
        \ANSWER/mem[8][2][13] ) );
  dp_1 \ANSWER/mem_reg[8][3][13]  ( .ip(n2519), .ck(clk), .q(
        \ANSWER/mem[8][3][13] ) );
  dp_1 \ANSWER/mem_reg[8][4][13]  ( .ip(n2518), .ck(clk), .q(
        \ANSWER/mem[8][4][13] ) );
  dp_1 \ANSWER/mem_reg[8][5][13]  ( .ip(n2517), .ck(clk), .q(
        \ANSWER/mem[8][5][13] ) );
  dp_1 \ANSWER/mem_reg[8][6][13]  ( .ip(n2516), .ck(clk), .q(
        \ANSWER/mem[8][6][13] ) );
  dp_1 \ANSWER/mem_reg[8][7][13]  ( .ip(n2515), .ck(clk), .q(
        \ANSWER/mem[8][7][13] ) );
  dp_1 \ANSWER/mem_reg[8][8][13]  ( .ip(n2514), .ck(clk), .q(
        \ANSWER/mem[8][8][13] ) );
  dp_1 \ANSWER/mem_reg[8][9][13]  ( .ip(n2513), .ck(clk), .q(
        \ANSWER/mem[8][9][13] ) );
  dp_1 \ANSWER/mem_reg[9][0][13]  ( .ip(n2512), .ck(clk), .q(
        \ANSWER/mem[9][0][13] ) );
  dp_1 \ANSWER/mem_reg[9][1][13]  ( .ip(n2511), .ck(clk), .q(
        \ANSWER/mem[9][1][13] ) );
  dp_1 \ANSWER/mem_reg[9][2][13]  ( .ip(n2510), .ck(clk), .q(
        \ANSWER/mem[9][2][13] ) );
  dp_1 \ANSWER/mem_reg[9][3][13]  ( .ip(n2509), .ck(clk), .q(
        \ANSWER/mem[9][3][13] ) );
  dp_1 \ANSWER/mem_reg[9][4][13]  ( .ip(n2508), .ck(clk), .q(
        \ANSWER/mem[9][4][13] ) );
  dp_1 \ANSWER/mem_reg[9][5][13]  ( .ip(n2507), .ck(clk), .q(
        \ANSWER/mem[9][5][13] ) );
  dp_1 \ANSWER/mem_reg[9][6][13]  ( .ip(n2506), .ck(clk), .q(
        \ANSWER/mem[9][6][13] ) );
  dp_1 \ANSWER/mem_reg[9][7][13]  ( .ip(n2505), .ck(clk), .q(
        \ANSWER/mem[9][7][13] ) );
  dp_1 \ANSWER/mem_reg[9][8][13]  ( .ip(n2504), .ck(clk), .q(
        \ANSWER/mem[9][8][13] ) );
  dp_1 \ANSWER/mem_reg[9][9][13]  ( .ip(n2503), .ck(clk), .q(
        \ANSWER/mem[9][9][13] ) );
  dp_1 \ANSWER/mem_reg[0][0][14]  ( .ip(n2502), .ck(clk), .q(
        \ANSWER/mem[0][0][14] ) );
  dp_1 \ANSWER/mem_reg[0][1][14]  ( .ip(n2501), .ck(clk), .q(
        \ANSWER/mem[0][1][14] ) );
  dp_1 \ANSWER/mem_reg[0][2][14]  ( .ip(n2500), .ck(clk), .q(
        \ANSWER/mem[0][2][14] ) );
  dp_1 \ANSWER/mem_reg[0][3][14]  ( .ip(n2499), .ck(clk), .q(
        \ANSWER/mem[0][3][14] ) );
  dp_1 \ANSWER/mem_reg[0][4][14]  ( .ip(n2498), .ck(clk), .q(
        \ANSWER/mem[0][4][14] ) );
  dp_1 \ANSWER/mem_reg[0][5][14]  ( .ip(n2497), .ck(clk), .q(
        \ANSWER/mem[0][5][14] ) );
  dp_1 \ANSWER/mem_reg[0][6][14]  ( .ip(n2496), .ck(clk), .q(
        \ANSWER/mem[0][6][14] ) );
  dp_1 \ANSWER/mem_reg[0][7][14]  ( .ip(n2495), .ck(clk), .q(
        \ANSWER/mem[0][7][14] ) );
  dp_1 \ANSWER/mem_reg[0][8][14]  ( .ip(n2494), .ck(clk), .q(
        \ANSWER/mem[0][8][14] ) );
  dp_1 \ANSWER/mem_reg[0][9][14]  ( .ip(n2493), .ck(clk), .q(
        \ANSWER/mem[0][9][14] ) );
  dp_1 \ANSWER/mem_reg[1][0][14]  ( .ip(n2492), .ck(clk), .q(
        \ANSWER/mem[1][0][14] ) );
  dp_1 \ANSWER/mem_reg[1][1][14]  ( .ip(n2491), .ck(clk), .q(
        \ANSWER/mem[1][1][14] ) );
  dp_1 \ANSWER/mem_reg[1][2][14]  ( .ip(n2490), .ck(clk), .q(
        \ANSWER/mem[1][2][14] ) );
  dp_1 \ANSWER/mem_reg[1][3][14]  ( .ip(n2489), .ck(clk), .q(
        \ANSWER/mem[1][3][14] ) );
  dp_1 \ANSWER/mem_reg[1][4][14]  ( .ip(n2488), .ck(clk), .q(
        \ANSWER/mem[1][4][14] ) );
  dp_1 \ANSWER/mem_reg[1][5][14]  ( .ip(n2487), .ck(clk), .q(
        \ANSWER/mem[1][5][14] ) );
  dp_1 \ANSWER/mem_reg[1][6][14]  ( .ip(n2486), .ck(clk), .q(
        \ANSWER/mem[1][6][14] ) );
  dp_1 \ANSWER/mem_reg[1][7][14]  ( .ip(n2485), .ck(clk), .q(
        \ANSWER/mem[1][7][14] ) );
  dp_1 \ANSWER/mem_reg[1][8][14]  ( .ip(n2484), .ck(clk), .q(
        \ANSWER/mem[1][8][14] ) );
  dp_1 \ANSWER/mem_reg[1][9][14]  ( .ip(n2483), .ck(clk), .q(
        \ANSWER/mem[1][9][14] ) );
  dp_1 \ANSWER/mem_reg[2][0][14]  ( .ip(n2482), .ck(clk), .q(
        \ANSWER/mem[2][0][14] ) );
  dp_1 \ANSWER/mem_reg[2][1][14]  ( .ip(n2481), .ck(clk), .q(
        \ANSWER/mem[2][1][14] ) );
  dp_1 \ANSWER/mem_reg[2][2][14]  ( .ip(n2480), .ck(clk), .q(
        \ANSWER/mem[2][2][14] ) );
  dp_1 \ANSWER/mem_reg[2][3][14]  ( .ip(n2479), .ck(clk), .q(
        \ANSWER/mem[2][3][14] ) );
  dp_1 \ANSWER/mem_reg[2][4][14]  ( .ip(n2478), .ck(clk), .q(
        \ANSWER/mem[2][4][14] ) );
  dp_1 \ANSWER/mem_reg[2][5][14]  ( .ip(n2477), .ck(clk), .q(
        \ANSWER/mem[2][5][14] ) );
  dp_1 \ANSWER/mem_reg[2][6][14]  ( .ip(n2476), .ck(clk), .q(
        \ANSWER/mem[2][6][14] ) );
  dp_1 \ANSWER/mem_reg[2][7][14]  ( .ip(n2475), .ck(clk), .q(
        \ANSWER/mem[2][7][14] ) );
  dp_1 \ANSWER/mem_reg[2][8][14]  ( .ip(n2474), .ck(clk), .q(
        \ANSWER/mem[2][8][14] ) );
  dp_1 \ANSWER/mem_reg[2][9][14]  ( .ip(n2473), .ck(clk), .q(
        \ANSWER/mem[2][9][14] ) );
  dp_1 \ANSWER/mem_reg[3][0][14]  ( .ip(n2472), .ck(clk), .q(
        \ANSWER/mem[3][0][14] ) );
  dp_1 \ANSWER/mem_reg[3][1][14]  ( .ip(n2471), .ck(clk), .q(
        \ANSWER/mem[3][1][14] ) );
  dp_1 \ANSWER/mem_reg[3][2][14]  ( .ip(n2470), .ck(clk), .q(
        \ANSWER/mem[3][2][14] ) );
  dp_1 \ANSWER/mem_reg[3][3][14]  ( .ip(n2469), .ck(clk), .q(
        \ANSWER/mem[3][3][14] ) );
  dp_1 \ANSWER/mem_reg[3][4][14]  ( .ip(n2468), .ck(clk), .q(
        \ANSWER/mem[3][4][14] ) );
  dp_1 \ANSWER/mem_reg[3][5][14]  ( .ip(n2467), .ck(clk), .q(
        \ANSWER/mem[3][5][14] ) );
  dp_1 \ANSWER/mem_reg[3][6][14]  ( .ip(n2466), .ck(clk), .q(
        \ANSWER/mem[3][6][14] ) );
  dp_1 \ANSWER/mem_reg[3][7][14]  ( .ip(n2465), .ck(clk), .q(
        \ANSWER/mem[3][7][14] ) );
  dp_1 \ANSWER/mem_reg[3][8][14]  ( .ip(n2464), .ck(clk), .q(
        \ANSWER/mem[3][8][14] ) );
  dp_1 \ANSWER/mem_reg[3][9][14]  ( .ip(n2463), .ck(clk), .q(
        \ANSWER/mem[3][9][14] ) );
  dp_1 \ANSWER/mem_reg[4][0][14]  ( .ip(n2462), .ck(clk), .q(
        \ANSWER/mem[4][0][14] ) );
  dp_1 \ANSWER/mem_reg[4][1][14]  ( .ip(n2461), .ck(clk), .q(
        \ANSWER/mem[4][1][14] ) );
  dp_1 \ANSWER/mem_reg[4][2][14]  ( .ip(n2460), .ck(clk), .q(
        \ANSWER/mem[4][2][14] ) );
  dp_1 \ANSWER/mem_reg[4][3][14]  ( .ip(n2459), .ck(clk), .q(
        \ANSWER/mem[4][3][14] ) );
  dp_1 \ANSWER/mem_reg[4][4][14]  ( .ip(n2458), .ck(clk), .q(
        \ANSWER/mem[4][4][14] ) );
  dp_1 \ANSWER/mem_reg[4][5][14]  ( .ip(n2457), .ck(clk), .q(
        \ANSWER/mem[4][5][14] ) );
  dp_1 \ANSWER/mem_reg[4][6][14]  ( .ip(n2456), .ck(clk), .q(
        \ANSWER/mem[4][6][14] ) );
  dp_1 \ANSWER/mem_reg[4][7][14]  ( .ip(n2455), .ck(clk), .q(
        \ANSWER/mem[4][7][14] ) );
  dp_1 \ANSWER/mem_reg[4][8][14]  ( .ip(n2454), .ck(clk), .q(
        \ANSWER/mem[4][8][14] ) );
  dp_1 \ANSWER/mem_reg[4][9][14]  ( .ip(n2453), .ck(clk), .q(
        \ANSWER/mem[4][9][14] ) );
  dp_1 \ANSWER/mem_reg[5][0][14]  ( .ip(n2452), .ck(clk), .q(
        \ANSWER/mem[5][0][14] ) );
  dp_1 \ANSWER/mem_reg[5][1][14]  ( .ip(n2451), .ck(clk), .q(
        \ANSWER/mem[5][1][14] ) );
  dp_1 \ANSWER/mem_reg[5][2][14]  ( .ip(n2450), .ck(clk), .q(
        \ANSWER/mem[5][2][14] ) );
  dp_1 \ANSWER/mem_reg[5][3][14]  ( .ip(n2449), .ck(clk), .q(
        \ANSWER/mem[5][3][14] ) );
  dp_1 \ANSWER/mem_reg[5][4][14]  ( .ip(n2448), .ck(clk), .q(
        \ANSWER/mem[5][4][14] ) );
  dp_1 \ANSWER/mem_reg[5][5][14]  ( .ip(n2447), .ck(clk), .q(
        \ANSWER/mem[5][5][14] ) );
  dp_1 \ANSWER/mem_reg[5][6][14]  ( .ip(n2446), .ck(clk), .q(
        \ANSWER/mem[5][6][14] ) );
  dp_1 \ANSWER/mem_reg[5][7][14]  ( .ip(n2445), .ck(clk), .q(
        \ANSWER/mem[5][7][14] ) );
  dp_1 \ANSWER/mem_reg[5][8][14]  ( .ip(n2444), .ck(clk), .q(
        \ANSWER/mem[5][8][14] ) );
  dp_1 \ANSWER/mem_reg[5][9][14]  ( .ip(n2443), .ck(clk), .q(
        \ANSWER/mem[5][9][14] ) );
  dp_1 \ANSWER/mem_reg[6][0][14]  ( .ip(n2442), .ck(clk), .q(
        \ANSWER/mem[6][0][14] ) );
  dp_1 \ANSWER/mem_reg[6][1][14]  ( .ip(n2441), .ck(clk), .q(
        \ANSWER/mem[6][1][14] ) );
  dp_1 \ANSWER/mem_reg[6][2][14]  ( .ip(n2440), .ck(clk), .q(
        \ANSWER/mem[6][2][14] ) );
  dp_1 \ANSWER/mem_reg[6][3][14]  ( .ip(n2439), .ck(clk), .q(
        \ANSWER/mem[6][3][14] ) );
  dp_1 \ANSWER/mem_reg[6][4][14]  ( .ip(n2438), .ck(clk), .q(
        \ANSWER/mem[6][4][14] ) );
  dp_1 \ANSWER/mem_reg[6][5][14]  ( .ip(n2437), .ck(clk), .q(
        \ANSWER/mem[6][5][14] ) );
  dp_1 \ANSWER/mem_reg[6][6][14]  ( .ip(n2436), .ck(clk), .q(
        \ANSWER/mem[6][6][14] ) );
  dp_1 \ANSWER/mem_reg[6][7][14]  ( .ip(n2435), .ck(clk), .q(
        \ANSWER/mem[6][7][14] ) );
  dp_1 \ANSWER/mem_reg[6][8][14]  ( .ip(n2434), .ck(clk), .q(
        \ANSWER/mem[6][8][14] ) );
  dp_1 \ANSWER/mem_reg[6][9][14]  ( .ip(n2433), .ck(clk), .q(
        \ANSWER/mem[6][9][14] ) );
  dp_1 \ANSWER/mem_reg[7][0][14]  ( .ip(n2432), .ck(clk), .q(
        \ANSWER/mem[7][0][14] ) );
  dp_1 \ANSWER/mem_reg[7][1][14]  ( .ip(n2431), .ck(clk), .q(
        \ANSWER/mem[7][1][14] ) );
  dp_1 \ANSWER/mem_reg[7][2][14]  ( .ip(n2430), .ck(clk), .q(
        \ANSWER/mem[7][2][14] ) );
  dp_1 \ANSWER/mem_reg[7][3][14]  ( .ip(n2429), .ck(clk), .q(
        \ANSWER/mem[7][3][14] ) );
  dp_1 \ANSWER/mem_reg[7][4][14]  ( .ip(n2428), .ck(clk), .q(
        \ANSWER/mem[7][4][14] ) );
  dp_1 \ANSWER/mem_reg[7][5][14]  ( .ip(n2427), .ck(clk), .q(
        \ANSWER/mem[7][5][14] ) );
  dp_1 \ANSWER/mem_reg[7][6][14]  ( .ip(n2426), .ck(clk), .q(
        \ANSWER/mem[7][6][14] ) );
  dp_1 \ANSWER/mem_reg[7][7][14]  ( .ip(n2425), .ck(clk), .q(
        \ANSWER/mem[7][7][14] ) );
  dp_1 \ANSWER/mem_reg[7][8][14]  ( .ip(n2424), .ck(clk), .q(
        \ANSWER/mem[7][8][14] ) );
  dp_1 \ANSWER/mem_reg[7][9][14]  ( .ip(n2423), .ck(clk), .q(
        \ANSWER/mem[7][9][14] ) );
  dp_1 \ANSWER/mem_reg[8][0][14]  ( .ip(n2422), .ck(clk), .q(
        \ANSWER/mem[8][0][14] ) );
  dp_1 \ANSWER/mem_reg[8][1][14]  ( .ip(n2421), .ck(clk), .q(
        \ANSWER/mem[8][1][14] ) );
  dp_1 \ANSWER/mem_reg[8][2][14]  ( .ip(n2420), .ck(clk), .q(
        \ANSWER/mem[8][2][14] ) );
  dp_1 \ANSWER/mem_reg[8][3][14]  ( .ip(n2419), .ck(clk), .q(
        \ANSWER/mem[8][3][14] ) );
  dp_1 \ANSWER/mem_reg[8][4][14]  ( .ip(n2418), .ck(clk), .q(
        \ANSWER/mem[8][4][14] ) );
  dp_1 \ANSWER/mem_reg[8][5][14]  ( .ip(n2417), .ck(clk), .q(
        \ANSWER/mem[8][5][14] ) );
  dp_1 \ANSWER/mem_reg[8][6][14]  ( .ip(n2416), .ck(clk), .q(
        \ANSWER/mem[8][6][14] ) );
  dp_1 \ANSWER/mem_reg[8][7][14]  ( .ip(n2415), .ck(clk), .q(
        \ANSWER/mem[8][7][14] ) );
  dp_1 \ANSWER/mem_reg[8][8][14]  ( .ip(n2414), .ck(clk), .q(
        \ANSWER/mem[8][8][14] ) );
  dp_1 \ANSWER/mem_reg[8][9][14]  ( .ip(n2413), .ck(clk), .q(
        \ANSWER/mem[8][9][14] ) );
  dp_1 \ANSWER/mem_reg[9][0][14]  ( .ip(n2412), .ck(clk), .q(
        \ANSWER/mem[9][0][14] ) );
  dp_1 \ANSWER/mem_reg[9][1][14]  ( .ip(n2411), .ck(clk), .q(
        \ANSWER/mem[9][1][14] ) );
  dp_1 \ANSWER/mem_reg[9][2][14]  ( .ip(n2410), .ck(clk), .q(
        \ANSWER/mem[9][2][14] ) );
  dp_1 \ANSWER/mem_reg[9][3][14]  ( .ip(n2409), .ck(clk), .q(
        \ANSWER/mem[9][3][14] ) );
  dp_1 \ANSWER/mem_reg[9][4][14]  ( .ip(n2408), .ck(clk), .q(
        \ANSWER/mem[9][4][14] ) );
  dp_1 \ANSWER/mem_reg[9][5][14]  ( .ip(n2407), .ck(clk), .q(
        \ANSWER/mem[9][5][14] ) );
  dp_1 \ANSWER/mem_reg[9][6][14]  ( .ip(n2406), .ck(clk), .q(
        \ANSWER/mem[9][6][14] ) );
  dp_1 \ANSWER/mem_reg[9][7][14]  ( .ip(n2405), .ck(clk), .q(
        \ANSWER/mem[9][7][14] ) );
  dp_1 \ANSWER/mem_reg[9][8][14]  ( .ip(n2404), .ck(clk), .q(
        \ANSWER/mem[9][8][14] ) );
  dp_1 \ANSWER/mem_reg[9][9][14]  ( .ip(n2403), .ck(clk), .q(
        \ANSWER/mem[9][9][14] ) );
  dp_1 \ANSWER/mem_reg[0][0][15]  ( .ip(n2402), .ck(clk), .q(
        \ANSWER/mem[0][0][15] ) );
  dp_1 \ANSWER/mem_reg[0][1][15]  ( .ip(n2401), .ck(clk), .q(
        \ANSWER/mem[0][1][15] ) );
  dp_1 \ANSWER/mem_reg[0][2][15]  ( .ip(n2400), .ck(clk), .q(
        \ANSWER/mem[0][2][15] ) );
  dp_1 \ANSWER/mem_reg[0][3][15]  ( .ip(n2399), .ck(clk), .q(
        \ANSWER/mem[0][3][15] ) );
  dp_1 \ANSWER/mem_reg[0][4][15]  ( .ip(n2398), .ck(clk), .q(
        \ANSWER/mem[0][4][15] ) );
  dp_1 \ANSWER/mem_reg[0][5][15]  ( .ip(n2397), .ck(clk), .q(
        \ANSWER/mem[0][5][15] ) );
  dp_1 \ANSWER/mem_reg[0][6][15]  ( .ip(n2396), .ck(clk), .q(
        \ANSWER/mem[0][6][15] ) );
  dp_1 \ANSWER/mem_reg[0][7][15]  ( .ip(n2395), .ck(clk), .q(
        \ANSWER/mem[0][7][15] ) );
  dp_1 \ANSWER/mem_reg[0][8][15]  ( .ip(n2394), .ck(clk), .q(
        \ANSWER/mem[0][8][15] ) );
  dp_1 \ANSWER/mem_reg[0][9][15]  ( .ip(n2393), .ck(clk), .q(
        \ANSWER/mem[0][9][15] ) );
  dp_1 \ANSWER/mem_reg[1][0][15]  ( .ip(n2392), .ck(clk), .q(
        \ANSWER/mem[1][0][15] ) );
  dp_1 \ANSWER/mem_reg[1][1][15]  ( .ip(n2391), .ck(clk), .q(
        \ANSWER/mem[1][1][15] ) );
  dp_1 \ANSWER/mem_reg[1][2][15]  ( .ip(n2390), .ck(clk), .q(
        \ANSWER/mem[1][2][15] ) );
  dp_1 \ANSWER/mem_reg[1][3][15]  ( .ip(n2389), .ck(clk), .q(
        \ANSWER/mem[1][3][15] ) );
  dp_1 \ANSWER/mem_reg[1][4][15]  ( .ip(n2388), .ck(clk), .q(
        \ANSWER/mem[1][4][15] ) );
  dp_1 \ANSWER/mem_reg[1][5][15]  ( .ip(n2387), .ck(clk), .q(
        \ANSWER/mem[1][5][15] ) );
  dp_1 \ANSWER/mem_reg[1][6][15]  ( .ip(n2386), .ck(clk), .q(
        \ANSWER/mem[1][6][15] ) );
  dp_1 \ANSWER/mem_reg[1][7][15]  ( .ip(n2385), .ck(clk), .q(
        \ANSWER/mem[1][7][15] ) );
  dp_1 \ANSWER/mem_reg[1][8][15]  ( .ip(n2384), .ck(clk), .q(
        \ANSWER/mem[1][8][15] ) );
  dp_1 \ANSWER/mem_reg[1][9][15]  ( .ip(n2383), .ck(clk), .q(
        \ANSWER/mem[1][9][15] ) );
  dp_1 \ANSWER/mem_reg[2][0][15]  ( .ip(n2382), .ck(clk), .q(
        \ANSWER/mem[2][0][15] ) );
  dp_1 \ANSWER/mem_reg[2][1][15]  ( .ip(n2381), .ck(clk), .q(
        \ANSWER/mem[2][1][15] ) );
  dp_1 \ANSWER/mem_reg[2][2][15]  ( .ip(n2380), .ck(clk), .q(
        \ANSWER/mem[2][2][15] ) );
  dp_1 \ANSWER/mem_reg[2][3][15]  ( .ip(n2379), .ck(clk), .q(
        \ANSWER/mem[2][3][15] ) );
  dp_1 \ANSWER/mem_reg[2][4][15]  ( .ip(n2378), .ck(clk), .q(
        \ANSWER/mem[2][4][15] ) );
  dp_1 \ANSWER/mem_reg[2][5][15]  ( .ip(n2377), .ck(clk), .q(
        \ANSWER/mem[2][5][15] ) );
  dp_1 \ANSWER/mem_reg[2][6][15]  ( .ip(n2376), .ck(clk), .q(
        \ANSWER/mem[2][6][15] ) );
  dp_1 \ANSWER/mem_reg[2][7][15]  ( .ip(n2375), .ck(clk), .q(
        \ANSWER/mem[2][7][15] ) );
  dp_1 \ANSWER/mem_reg[2][8][15]  ( .ip(n2374), .ck(clk), .q(
        \ANSWER/mem[2][8][15] ) );
  dp_1 \ANSWER/mem_reg[2][9][15]  ( .ip(n2373), .ck(clk), .q(
        \ANSWER/mem[2][9][15] ) );
  dp_1 \ANSWER/mem_reg[3][0][15]  ( .ip(n2372), .ck(clk), .q(
        \ANSWER/mem[3][0][15] ) );
  dp_1 \ANSWER/mem_reg[3][1][15]  ( .ip(n2371), .ck(clk), .q(
        \ANSWER/mem[3][1][15] ) );
  dp_1 \ANSWER/mem_reg[3][2][15]  ( .ip(n2370), .ck(clk), .q(
        \ANSWER/mem[3][2][15] ) );
  dp_1 \ANSWER/mem_reg[3][3][15]  ( .ip(n2369), .ck(clk), .q(
        \ANSWER/mem[3][3][15] ) );
  dp_1 \ANSWER/mem_reg[3][4][15]  ( .ip(n2368), .ck(clk), .q(
        \ANSWER/mem[3][4][15] ) );
  dp_1 \ANSWER/mem_reg[3][5][15]  ( .ip(n2367), .ck(clk), .q(
        \ANSWER/mem[3][5][15] ) );
  dp_1 \ANSWER/mem_reg[3][6][15]  ( .ip(n2366), .ck(clk), .q(
        \ANSWER/mem[3][6][15] ) );
  dp_1 \ANSWER/mem_reg[3][7][15]  ( .ip(n2365), .ck(clk), .q(
        \ANSWER/mem[3][7][15] ) );
  dp_1 \ANSWER/mem_reg[3][8][15]  ( .ip(n2364), .ck(clk), .q(
        \ANSWER/mem[3][8][15] ) );
  dp_1 \ANSWER/mem_reg[3][9][15]  ( .ip(n2363), .ck(clk), .q(
        \ANSWER/mem[3][9][15] ) );
  dp_1 \ANSWER/mem_reg[4][0][15]  ( .ip(n2362), .ck(clk), .q(
        \ANSWER/mem[4][0][15] ) );
  dp_1 \ANSWER/mem_reg[4][1][15]  ( .ip(n2361), .ck(clk), .q(
        \ANSWER/mem[4][1][15] ) );
  dp_1 \ANSWER/mem_reg[4][2][15]  ( .ip(n2360), .ck(clk), .q(
        \ANSWER/mem[4][2][15] ) );
  dp_1 \ANSWER/mem_reg[4][3][15]  ( .ip(n2359), .ck(clk), .q(
        \ANSWER/mem[4][3][15] ) );
  dp_1 \ANSWER/mem_reg[4][4][15]  ( .ip(n2358), .ck(clk), .q(
        \ANSWER/mem[4][4][15] ) );
  dp_1 \ANSWER/mem_reg[4][5][15]  ( .ip(n2357), .ck(clk), .q(
        \ANSWER/mem[4][5][15] ) );
  dp_1 \ANSWER/mem_reg[4][6][15]  ( .ip(n2356), .ck(clk), .q(
        \ANSWER/mem[4][6][15] ) );
  dp_1 \ANSWER/mem_reg[4][7][15]  ( .ip(n2355), .ck(clk), .q(
        \ANSWER/mem[4][7][15] ) );
  dp_1 \ANSWER/mem_reg[4][8][15]  ( .ip(n2354), .ck(clk), .q(
        \ANSWER/mem[4][8][15] ) );
  dp_1 \ANSWER/mem_reg[4][9][15]  ( .ip(n2353), .ck(clk), .q(
        \ANSWER/mem[4][9][15] ) );
  dp_1 \ANSWER/mem_reg[5][0][15]  ( .ip(n2352), .ck(clk), .q(
        \ANSWER/mem[5][0][15] ) );
  dp_1 \ANSWER/mem_reg[5][1][15]  ( .ip(n2351), .ck(clk), .q(
        \ANSWER/mem[5][1][15] ) );
  dp_1 \ANSWER/mem_reg[5][2][15]  ( .ip(n2350), .ck(clk), .q(
        \ANSWER/mem[5][2][15] ) );
  dp_1 \ANSWER/mem_reg[5][3][15]  ( .ip(n2349), .ck(clk), .q(
        \ANSWER/mem[5][3][15] ) );
  dp_1 \ANSWER/mem_reg[5][4][15]  ( .ip(n2348), .ck(clk), .q(
        \ANSWER/mem[5][4][15] ) );
  dp_1 \ANSWER/mem_reg[5][5][15]  ( .ip(n2347), .ck(clk), .q(
        \ANSWER/mem[5][5][15] ) );
  dp_1 \ANSWER/mem_reg[5][6][15]  ( .ip(n2346), .ck(clk), .q(
        \ANSWER/mem[5][6][15] ) );
  dp_1 \ANSWER/mem_reg[5][7][15]  ( .ip(n2345), .ck(clk), .q(
        \ANSWER/mem[5][7][15] ) );
  dp_1 \ANSWER/mem_reg[5][8][15]  ( .ip(n2344), .ck(clk), .q(
        \ANSWER/mem[5][8][15] ) );
  dp_1 \ANSWER/mem_reg[5][9][15]  ( .ip(n2343), .ck(clk), .q(
        \ANSWER/mem[5][9][15] ) );
  dp_1 \ANSWER/mem_reg[6][0][15]  ( .ip(n2342), .ck(clk), .q(
        \ANSWER/mem[6][0][15] ) );
  dp_1 \ANSWER/mem_reg[6][1][15]  ( .ip(n2341), .ck(clk), .q(
        \ANSWER/mem[6][1][15] ) );
  dp_1 \ANSWER/mem_reg[6][2][15]  ( .ip(n2340), .ck(clk), .q(
        \ANSWER/mem[6][2][15] ) );
  dp_1 \ANSWER/mem_reg[6][3][15]  ( .ip(n2339), .ck(clk), .q(
        \ANSWER/mem[6][3][15] ) );
  dp_1 \ANSWER/mem_reg[6][4][15]  ( .ip(n2338), .ck(clk), .q(
        \ANSWER/mem[6][4][15] ) );
  dp_1 \ANSWER/mem_reg[6][5][15]  ( .ip(n2337), .ck(clk), .q(
        \ANSWER/mem[6][5][15] ) );
  dp_1 \ANSWER/mem_reg[6][6][15]  ( .ip(n2336), .ck(clk), .q(
        \ANSWER/mem[6][6][15] ) );
  dp_1 \ANSWER/mem_reg[6][7][15]  ( .ip(n2335), .ck(clk), .q(
        \ANSWER/mem[6][7][15] ) );
  dp_1 \ANSWER/mem_reg[6][8][15]  ( .ip(n2334), .ck(clk), .q(
        \ANSWER/mem[6][8][15] ) );
  dp_1 \ANSWER/mem_reg[6][9][15]  ( .ip(n2333), .ck(clk), .q(
        \ANSWER/mem[6][9][15] ) );
  dp_1 \ANSWER/mem_reg[7][0][15]  ( .ip(n2332), .ck(clk), .q(
        \ANSWER/mem[7][0][15] ) );
  dp_1 \ANSWER/mem_reg[7][1][15]  ( .ip(n2331), .ck(clk), .q(
        \ANSWER/mem[7][1][15] ) );
  dp_1 \ANSWER/mem_reg[7][2][15]  ( .ip(n2330), .ck(clk), .q(
        \ANSWER/mem[7][2][15] ) );
  dp_1 \ANSWER/mem_reg[7][3][15]  ( .ip(n2329), .ck(clk), .q(
        \ANSWER/mem[7][3][15] ) );
  dp_1 \ANSWER/mem_reg[7][4][15]  ( .ip(n2328), .ck(clk), .q(
        \ANSWER/mem[7][4][15] ) );
  dp_1 \ANSWER/mem_reg[7][5][15]  ( .ip(n2327), .ck(clk), .q(
        \ANSWER/mem[7][5][15] ) );
  dp_1 \ANSWER/mem_reg[7][6][15]  ( .ip(n2326), .ck(clk), .q(
        \ANSWER/mem[7][6][15] ) );
  dp_1 \ANSWER/mem_reg[7][7][15]  ( .ip(n2325), .ck(clk), .q(
        \ANSWER/mem[7][7][15] ) );
  dp_1 \ANSWER/mem_reg[7][8][15]  ( .ip(n2324), .ck(clk), .q(
        \ANSWER/mem[7][8][15] ) );
  dp_1 \ANSWER/mem_reg[7][9][15]  ( .ip(n2323), .ck(clk), .q(
        \ANSWER/mem[7][9][15] ) );
  dp_1 \ANSWER/mem_reg[8][0][15]  ( .ip(n2322), .ck(clk), .q(
        \ANSWER/mem[8][0][15] ) );
  dp_1 \ANSWER/mem_reg[8][1][15]  ( .ip(n2321), .ck(clk), .q(
        \ANSWER/mem[8][1][15] ) );
  dp_1 \ANSWER/mem_reg[8][2][15]  ( .ip(n2320), .ck(clk), .q(
        \ANSWER/mem[8][2][15] ) );
  dp_1 \ANSWER/mem_reg[8][3][15]  ( .ip(n2319), .ck(clk), .q(
        \ANSWER/mem[8][3][15] ) );
  dp_1 \ANSWER/mem_reg[8][4][15]  ( .ip(n2318), .ck(clk), .q(
        \ANSWER/mem[8][4][15] ) );
  dp_1 \ANSWER/mem_reg[8][5][15]  ( .ip(n2317), .ck(clk), .q(
        \ANSWER/mem[8][5][15] ) );
  dp_1 \ANSWER/mem_reg[8][6][15]  ( .ip(n2316), .ck(clk), .q(
        \ANSWER/mem[8][6][15] ) );
  dp_1 \ANSWER/mem_reg[8][7][15]  ( .ip(n2315), .ck(clk), .q(
        \ANSWER/mem[8][7][15] ) );
  dp_1 \ANSWER/mem_reg[8][8][15]  ( .ip(n2314), .ck(clk), .q(
        \ANSWER/mem[8][8][15] ) );
  dp_1 \ANSWER/mem_reg[8][9][15]  ( .ip(n2313), .ck(clk), .q(
        \ANSWER/mem[8][9][15] ) );
  dp_1 \ANSWER/mem_reg[9][0][15]  ( .ip(n2312), .ck(clk), .q(
        \ANSWER/mem[9][0][15] ) );
  dp_1 \ANSWER/mem_reg[9][1][15]  ( .ip(n2311), .ck(clk), .q(
        \ANSWER/mem[9][1][15] ) );
  dp_1 \ANSWER/mem_reg[9][2][15]  ( .ip(n2310), .ck(clk), .q(
        \ANSWER/mem[9][2][15] ) );
  dp_1 \ANSWER/mem_reg[9][3][15]  ( .ip(n2309), .ck(clk), .q(
        \ANSWER/mem[9][3][15] ) );
  dp_1 \ANSWER/mem_reg[9][4][15]  ( .ip(n2308), .ck(clk), .q(
        \ANSWER/mem[9][4][15] ) );
  dp_1 \ANSWER/mem_reg[9][5][15]  ( .ip(n2307), .ck(clk), .q(
        \ANSWER/mem[9][5][15] ) );
  dp_1 \ANSWER/mem_reg[9][6][15]  ( .ip(n2306), .ck(clk), .q(
        \ANSWER/mem[9][6][15] ) );
  dp_1 \ANSWER/mem_reg[9][7][15]  ( .ip(n2305), .ck(clk), .q(
        \ANSWER/mem[9][7][15] ) );
  dp_1 \ANSWER/mem_reg[9][8][15]  ( .ip(n2304), .ck(clk), .q(
        \ANSWER/mem[9][8][15] ) );
  dp_1 \ANSWER/mem_reg[9][9][15]  ( .ip(n2303), .ck(clk), .q(
        \ANSWER/mem[9][9][15] ) );
  dp_1 \SIGMOID/lut_out_reg[0]  ( .ip(n3910), .ck(clk), .q(\SIGMOID/N64 ) );
  dp_1 \ANSWER/mem_reg[0][0][0]  ( .ip(n3902), .ck(clk), .q(
        \ANSWER/mem[0][0][0] ) );
  dp_1 \ANSWER/mem_reg[0][1][0]  ( .ip(n3901), .ck(clk), .q(
        \ANSWER/mem[0][1][0] ) );
  dp_1 \ANSWER/mem_reg[0][2][0]  ( .ip(n3900), .ck(clk), .q(
        \ANSWER/mem[0][2][0] ) );
  dp_1 \ANSWER/mem_reg[0][3][0]  ( .ip(n3899), .ck(clk), .q(
        \ANSWER/mem[0][3][0] ) );
  dp_1 \ANSWER/mem_reg[0][4][0]  ( .ip(n3898), .ck(clk), .q(
        \ANSWER/mem[0][4][0] ) );
  dp_1 \ANSWER/mem_reg[0][5][0]  ( .ip(n3897), .ck(clk), .q(
        \ANSWER/mem[0][5][0] ) );
  dp_1 \ANSWER/mem_reg[0][6][0]  ( .ip(n3896), .ck(clk), .q(
        \ANSWER/mem[0][6][0] ) );
  dp_1 \ANSWER/mem_reg[0][7][0]  ( .ip(n3895), .ck(clk), .q(
        \ANSWER/mem[0][7][0] ) );
  dp_1 \ANSWER/mem_reg[0][8][0]  ( .ip(n3894), .ck(clk), .q(
        \ANSWER/mem[0][8][0] ) );
  dp_1 \ANSWER/mem_reg[0][9][0]  ( .ip(n3893), .ck(clk), .q(
        \ANSWER/mem[0][9][0] ) );
  dp_1 \ANSWER/mem_reg[1][0][0]  ( .ip(n3892), .ck(clk), .q(
        \ANSWER/mem[1][0][0] ) );
  dp_1 \ANSWER/mem_reg[1][1][0]  ( .ip(n3891), .ck(clk), .q(
        \ANSWER/mem[1][1][0] ) );
  dp_1 \ANSWER/mem_reg[1][2][0]  ( .ip(n3890), .ck(clk), .q(
        \ANSWER/mem[1][2][0] ) );
  dp_1 \ANSWER/mem_reg[1][3][0]  ( .ip(n3889), .ck(clk), .q(
        \ANSWER/mem[1][3][0] ) );
  dp_1 \ANSWER/mem_reg[1][4][0]  ( .ip(n3888), .ck(clk), .q(
        \ANSWER/mem[1][4][0] ) );
  dp_1 \ANSWER/mem_reg[1][5][0]  ( .ip(n3887), .ck(clk), .q(
        \ANSWER/mem[1][5][0] ) );
  dp_1 \ANSWER/mem_reg[1][6][0]  ( .ip(n3886), .ck(clk), .q(
        \ANSWER/mem[1][6][0] ) );
  dp_1 \ANSWER/mem_reg[1][7][0]  ( .ip(n3885), .ck(clk), .q(
        \ANSWER/mem[1][7][0] ) );
  dp_1 \ANSWER/mem_reg[1][8][0]  ( .ip(n3884), .ck(clk), .q(
        \ANSWER/mem[1][8][0] ) );
  dp_1 \ANSWER/mem_reg[1][9][0]  ( .ip(n3883), .ck(clk), .q(
        \ANSWER/mem[1][9][0] ) );
  dp_1 \ANSWER/mem_reg[2][0][0]  ( .ip(n3882), .ck(clk), .q(
        \ANSWER/mem[2][0][0] ) );
  dp_1 \ANSWER/mem_reg[2][1][0]  ( .ip(n3881), .ck(clk), .q(
        \ANSWER/mem[2][1][0] ) );
  dp_1 \ANSWER/mem_reg[2][2][0]  ( .ip(n3880), .ck(clk), .q(
        \ANSWER/mem[2][2][0] ) );
  dp_1 \ANSWER/mem_reg[2][3][0]  ( .ip(n3879), .ck(clk), .q(
        \ANSWER/mem[2][3][0] ) );
  dp_1 \ANSWER/mem_reg[2][4][0]  ( .ip(n3878), .ck(clk), .q(
        \ANSWER/mem[2][4][0] ) );
  dp_1 \ANSWER/mem_reg[2][5][0]  ( .ip(n3877), .ck(clk), .q(
        \ANSWER/mem[2][5][0] ) );
  dp_1 \ANSWER/mem_reg[2][6][0]  ( .ip(n3876), .ck(clk), .q(
        \ANSWER/mem[2][6][0] ) );
  dp_1 \ANSWER/mem_reg[2][7][0]  ( .ip(n3875), .ck(clk), .q(
        \ANSWER/mem[2][7][0] ) );
  dp_1 \ANSWER/mem_reg[2][8][0]  ( .ip(n3874), .ck(clk), .q(
        \ANSWER/mem[2][8][0] ) );
  dp_1 \ANSWER/mem_reg[2][9][0]  ( .ip(n3873), .ck(clk), .q(
        \ANSWER/mem[2][9][0] ) );
  dp_1 \ANSWER/mem_reg[3][0][0]  ( .ip(n3872), .ck(clk), .q(
        \ANSWER/mem[3][0][0] ) );
  dp_1 \ANSWER/mem_reg[3][1][0]  ( .ip(n3871), .ck(clk), .q(
        \ANSWER/mem[3][1][0] ) );
  dp_1 \ANSWER/mem_reg[3][2][0]  ( .ip(n3870), .ck(clk), .q(
        \ANSWER/mem[3][2][0] ) );
  dp_1 \ANSWER/mem_reg[3][3][0]  ( .ip(n3869), .ck(clk), .q(
        \ANSWER/mem[3][3][0] ) );
  dp_1 \ANSWER/mem_reg[3][4][0]  ( .ip(n3868), .ck(clk), .q(
        \ANSWER/mem[3][4][0] ) );
  dp_1 \ANSWER/mem_reg[3][5][0]  ( .ip(n3867), .ck(clk), .q(
        \ANSWER/mem[3][5][0] ) );
  dp_1 \ANSWER/mem_reg[3][6][0]  ( .ip(n3866), .ck(clk), .q(
        \ANSWER/mem[3][6][0] ) );
  dp_1 \ANSWER/mem_reg[3][7][0]  ( .ip(n3865), .ck(clk), .q(
        \ANSWER/mem[3][7][0] ) );
  dp_1 \ANSWER/mem_reg[3][8][0]  ( .ip(n3864), .ck(clk), .q(
        \ANSWER/mem[3][8][0] ) );
  dp_1 \ANSWER/mem_reg[3][9][0]  ( .ip(n3863), .ck(clk), .q(
        \ANSWER/mem[3][9][0] ) );
  dp_1 \ANSWER/mem_reg[4][0][0]  ( .ip(n3862), .ck(clk), .q(
        \ANSWER/mem[4][0][0] ) );
  dp_1 \ANSWER/mem_reg[4][1][0]  ( .ip(n3861), .ck(clk), .q(
        \ANSWER/mem[4][1][0] ) );
  dp_1 \ANSWER/mem_reg[4][2][0]  ( .ip(n3860), .ck(clk), .q(
        \ANSWER/mem[4][2][0] ) );
  dp_1 \ANSWER/mem_reg[4][3][0]  ( .ip(n3859), .ck(clk), .q(
        \ANSWER/mem[4][3][0] ) );
  dp_1 \ANSWER/mem_reg[4][4][0]  ( .ip(n3858), .ck(clk), .q(
        \ANSWER/mem[4][4][0] ) );
  dp_1 \ANSWER/mem_reg[4][5][0]  ( .ip(n3857), .ck(clk), .q(
        \ANSWER/mem[4][5][0] ) );
  dp_1 \ANSWER/mem_reg[4][6][0]  ( .ip(n3856), .ck(clk), .q(
        \ANSWER/mem[4][6][0] ) );
  dp_1 \ANSWER/mem_reg[4][7][0]  ( .ip(n3855), .ck(clk), .q(
        \ANSWER/mem[4][7][0] ) );
  dp_1 \ANSWER/mem_reg[4][8][0]  ( .ip(n3854), .ck(clk), .q(
        \ANSWER/mem[4][8][0] ) );
  dp_1 \ANSWER/mem_reg[4][9][0]  ( .ip(n3853), .ck(clk), .q(
        \ANSWER/mem[4][9][0] ) );
  dp_1 \ANSWER/mem_reg[5][0][0]  ( .ip(n3852), .ck(clk), .q(
        \ANSWER/mem[5][0][0] ) );
  dp_1 \ANSWER/mem_reg[5][1][0]  ( .ip(n3851), .ck(clk), .q(
        \ANSWER/mem[5][1][0] ) );
  dp_1 \ANSWER/mem_reg[5][2][0]  ( .ip(n3850), .ck(clk), .q(
        \ANSWER/mem[5][2][0] ) );
  dp_1 \ANSWER/mem_reg[5][3][0]  ( .ip(n3849), .ck(clk), .q(
        \ANSWER/mem[5][3][0] ) );
  dp_1 \ANSWER/mem_reg[5][4][0]  ( .ip(n3848), .ck(clk), .q(
        \ANSWER/mem[5][4][0] ) );
  dp_1 \ANSWER/mem_reg[5][5][0]  ( .ip(n3847), .ck(clk), .q(
        \ANSWER/mem[5][5][0] ) );
  dp_1 \ANSWER/mem_reg[5][6][0]  ( .ip(n3846), .ck(clk), .q(
        \ANSWER/mem[5][6][0] ) );
  dp_1 \ANSWER/mem_reg[5][7][0]  ( .ip(n3845), .ck(clk), .q(
        \ANSWER/mem[5][7][0] ) );
  dp_1 \ANSWER/mem_reg[5][8][0]  ( .ip(n3844), .ck(clk), .q(
        \ANSWER/mem[5][8][0] ) );
  dp_1 \ANSWER/mem_reg[5][9][0]  ( .ip(n3843), .ck(clk), .q(
        \ANSWER/mem[5][9][0] ) );
  dp_1 \ANSWER/mem_reg[6][0][0]  ( .ip(n3842), .ck(clk), .q(
        \ANSWER/mem[6][0][0] ) );
  dp_1 \ANSWER/mem_reg[6][1][0]  ( .ip(n3841), .ck(clk), .q(
        \ANSWER/mem[6][1][0] ) );
  dp_1 \ANSWER/mem_reg[6][2][0]  ( .ip(n3840), .ck(clk), .q(
        \ANSWER/mem[6][2][0] ) );
  dp_1 \ANSWER/mem_reg[6][3][0]  ( .ip(n3839), .ck(clk), .q(
        \ANSWER/mem[6][3][0] ) );
  dp_1 \ANSWER/mem_reg[6][4][0]  ( .ip(n3838), .ck(clk), .q(
        \ANSWER/mem[6][4][0] ) );
  dp_1 \ANSWER/mem_reg[6][5][0]  ( .ip(n3837), .ck(clk), .q(
        \ANSWER/mem[6][5][0] ) );
  dp_1 \ANSWER/mem_reg[6][6][0]  ( .ip(n3836), .ck(clk), .q(
        \ANSWER/mem[6][6][0] ) );
  dp_1 \ANSWER/mem_reg[6][7][0]  ( .ip(n3835), .ck(clk), .q(
        \ANSWER/mem[6][7][0] ) );
  dp_1 \ANSWER/mem_reg[6][8][0]  ( .ip(n3834), .ck(clk), .q(
        \ANSWER/mem[6][8][0] ) );
  dp_1 \ANSWER/mem_reg[6][9][0]  ( .ip(n3833), .ck(clk), .q(
        \ANSWER/mem[6][9][0] ) );
  dp_1 \ANSWER/mem_reg[7][0][0]  ( .ip(n3832), .ck(clk), .q(
        \ANSWER/mem[7][0][0] ) );
  dp_1 \ANSWER/mem_reg[7][1][0]  ( .ip(n3831), .ck(clk), .q(
        \ANSWER/mem[7][1][0] ) );
  dp_1 \ANSWER/mem_reg[7][2][0]  ( .ip(n3830), .ck(clk), .q(
        \ANSWER/mem[7][2][0] ) );
  dp_1 \ANSWER/mem_reg[7][3][0]  ( .ip(n3829), .ck(clk), .q(
        \ANSWER/mem[7][3][0] ) );
  dp_1 \ANSWER/mem_reg[7][4][0]  ( .ip(n3828), .ck(clk), .q(
        \ANSWER/mem[7][4][0] ) );
  dp_1 \ANSWER/mem_reg[7][5][0]  ( .ip(n3827), .ck(clk), .q(
        \ANSWER/mem[7][5][0] ) );
  dp_1 \ANSWER/mem_reg[7][6][0]  ( .ip(n3826), .ck(clk), .q(
        \ANSWER/mem[7][6][0] ) );
  dp_1 \ANSWER/mem_reg[7][7][0]  ( .ip(n3825), .ck(clk), .q(
        \ANSWER/mem[7][7][0] ) );
  dp_1 \ANSWER/mem_reg[7][8][0]  ( .ip(n3824), .ck(clk), .q(
        \ANSWER/mem[7][8][0] ) );
  dp_1 \ANSWER/mem_reg[7][9][0]  ( .ip(n3823), .ck(clk), .q(
        \ANSWER/mem[7][9][0] ) );
  dp_1 \ANSWER/mem_reg[8][0][0]  ( .ip(n3822), .ck(clk), .q(
        \ANSWER/mem[8][0][0] ) );
  dp_1 \ANSWER/mem_reg[8][1][0]  ( .ip(n3821), .ck(clk), .q(
        \ANSWER/mem[8][1][0] ) );
  dp_1 \ANSWER/mem_reg[8][2][0]  ( .ip(n3820), .ck(clk), .q(
        \ANSWER/mem[8][2][0] ) );
  dp_1 \ANSWER/mem_reg[8][3][0]  ( .ip(n3819), .ck(clk), .q(
        \ANSWER/mem[8][3][0] ) );
  dp_1 \ANSWER/mem_reg[8][4][0]  ( .ip(n3818), .ck(clk), .q(
        \ANSWER/mem[8][4][0] ) );
  dp_1 \ANSWER/mem_reg[8][5][0]  ( .ip(n3817), .ck(clk), .q(
        \ANSWER/mem[8][5][0] ) );
  dp_1 \ANSWER/mem_reg[8][6][0]  ( .ip(n3816), .ck(clk), .q(
        \ANSWER/mem[8][6][0] ) );
  dp_1 \ANSWER/mem_reg[8][7][0]  ( .ip(n3815), .ck(clk), .q(
        \ANSWER/mem[8][7][0] ) );
  dp_1 \ANSWER/mem_reg[8][8][0]  ( .ip(n3814), .ck(clk), .q(
        \ANSWER/mem[8][8][0] ) );
  dp_1 \ANSWER/mem_reg[8][9][0]  ( .ip(n3813), .ck(clk), .q(
        \ANSWER/mem[8][9][0] ) );
  dp_1 \ANSWER/mem_reg[9][0][0]  ( .ip(n3812), .ck(clk), .q(
        \ANSWER/mem[9][0][0] ) );
  dp_1 \ANSWER/mem_reg[9][1][0]  ( .ip(n3811), .ck(clk), .q(
        \ANSWER/mem[9][1][0] ) );
  dp_1 \ANSWER/mem_reg[9][2][0]  ( .ip(n3810), .ck(clk), .q(
        \ANSWER/mem[9][2][0] ) );
  dp_1 \ANSWER/mem_reg[9][3][0]  ( .ip(n3809), .ck(clk), .q(
        \ANSWER/mem[9][3][0] ) );
  dp_1 \ANSWER/mem_reg[9][4][0]  ( .ip(n3808), .ck(clk), .q(
        \ANSWER/mem[9][4][0] ) );
  dp_1 \ANSWER/mem_reg[9][5][0]  ( .ip(n3807), .ck(clk), .q(
        \ANSWER/mem[9][5][0] ) );
  dp_1 \ANSWER/mem_reg[9][6][0]  ( .ip(n3806), .ck(clk), .q(
        \ANSWER/mem[9][6][0] ) );
  dp_1 \ANSWER/mem_reg[9][7][0]  ( .ip(n3805), .ck(clk), .q(
        \ANSWER/mem[9][7][0] ) );
  dp_1 \ANSWER/mem_reg[9][8][0]  ( .ip(n3804), .ck(clk), .q(
        \ANSWER/mem[9][8][0] ) );
  dp_1 \ANSWER/mem_reg[9][9][0]  ( .ip(n3803), .ck(clk), .q(
        \ANSWER/mem[9][9][0] ) );
  dp_1 \SIGMOID/lut_out_reg[1]  ( .ip(n3909), .ck(clk), .q(
        \SIGMOID/lut_out [1]) );
  dp_1 \ANSWER/mem_reg[0][0][1]  ( .ip(n3802), .ck(clk), .q(
        \ANSWER/mem[0][0][1] ) );
  dp_1 \ANSWER/mem_reg[0][1][1]  ( .ip(n3801), .ck(clk), .q(
        \ANSWER/mem[0][1][1] ) );
  dp_1 \ANSWER/mem_reg[0][2][1]  ( .ip(n3800), .ck(clk), .q(
        \ANSWER/mem[0][2][1] ) );
  dp_1 \ANSWER/mem_reg[0][3][1]  ( .ip(n3799), .ck(clk), .q(
        \ANSWER/mem[0][3][1] ) );
  dp_1 \ANSWER/mem_reg[0][4][1]  ( .ip(n3798), .ck(clk), .q(
        \ANSWER/mem[0][4][1] ) );
  dp_1 \ANSWER/mem_reg[0][5][1]  ( .ip(n3797), .ck(clk), .q(
        \ANSWER/mem[0][5][1] ) );
  dp_1 \ANSWER/mem_reg[0][6][1]  ( .ip(n3796), .ck(clk), .q(
        \ANSWER/mem[0][6][1] ) );
  dp_1 \ANSWER/mem_reg[0][7][1]  ( .ip(n3795), .ck(clk), .q(
        \ANSWER/mem[0][7][1] ) );
  dp_1 \ANSWER/mem_reg[0][8][1]  ( .ip(n3794), .ck(clk), .q(
        \ANSWER/mem[0][8][1] ) );
  dp_1 \ANSWER/mem_reg[0][9][1]  ( .ip(n3793), .ck(clk), .q(
        \ANSWER/mem[0][9][1] ) );
  dp_1 \ANSWER/mem_reg[1][0][1]  ( .ip(n3792), .ck(clk), .q(
        \ANSWER/mem[1][0][1] ) );
  dp_1 \ANSWER/mem_reg[1][1][1]  ( .ip(n3791), .ck(clk), .q(
        \ANSWER/mem[1][1][1] ) );
  dp_1 \ANSWER/mem_reg[1][2][1]  ( .ip(n3790), .ck(clk), .q(
        \ANSWER/mem[1][2][1] ) );
  dp_1 \ANSWER/mem_reg[1][3][1]  ( .ip(n3789), .ck(clk), .q(
        \ANSWER/mem[1][3][1] ) );
  dp_1 \ANSWER/mem_reg[1][4][1]  ( .ip(n3788), .ck(clk), .q(
        \ANSWER/mem[1][4][1] ) );
  dp_1 \ANSWER/mem_reg[1][5][1]  ( .ip(n3787), .ck(clk), .q(
        \ANSWER/mem[1][5][1] ) );
  dp_1 \ANSWER/mem_reg[1][6][1]  ( .ip(n3786), .ck(clk), .q(
        \ANSWER/mem[1][6][1] ) );
  dp_1 \ANSWER/mem_reg[1][7][1]  ( .ip(n3785), .ck(clk), .q(
        \ANSWER/mem[1][7][1] ) );
  dp_1 \ANSWER/mem_reg[1][8][1]  ( .ip(n3784), .ck(clk), .q(
        \ANSWER/mem[1][8][1] ) );
  dp_1 \ANSWER/mem_reg[1][9][1]  ( .ip(n3783), .ck(clk), .q(
        \ANSWER/mem[1][9][1] ) );
  dp_1 \ANSWER/mem_reg[2][0][1]  ( .ip(n3782), .ck(clk), .q(
        \ANSWER/mem[2][0][1] ) );
  dp_1 \ANSWER/mem_reg[2][1][1]  ( .ip(n3781), .ck(clk), .q(
        \ANSWER/mem[2][1][1] ) );
  dp_1 \ANSWER/mem_reg[2][2][1]  ( .ip(n3780), .ck(clk), .q(
        \ANSWER/mem[2][2][1] ) );
  dp_1 \ANSWER/mem_reg[2][3][1]  ( .ip(n3779), .ck(clk), .q(
        \ANSWER/mem[2][3][1] ) );
  dp_1 \ANSWER/mem_reg[2][4][1]  ( .ip(n3778), .ck(clk), .q(
        \ANSWER/mem[2][4][1] ) );
  dp_1 \ANSWER/mem_reg[2][5][1]  ( .ip(n3777), .ck(clk), .q(
        \ANSWER/mem[2][5][1] ) );
  dp_1 \ANSWER/mem_reg[2][6][1]  ( .ip(n3776), .ck(clk), .q(
        \ANSWER/mem[2][6][1] ) );
  dp_1 \ANSWER/mem_reg[2][7][1]  ( .ip(n3775), .ck(clk), .q(
        \ANSWER/mem[2][7][1] ) );
  dp_1 \ANSWER/mem_reg[2][8][1]  ( .ip(n3774), .ck(clk), .q(
        \ANSWER/mem[2][8][1] ) );
  dp_1 \ANSWER/mem_reg[2][9][1]  ( .ip(n3773), .ck(clk), .q(
        \ANSWER/mem[2][9][1] ) );
  dp_1 \ANSWER/mem_reg[3][0][1]  ( .ip(n3772), .ck(clk), .q(
        \ANSWER/mem[3][0][1] ) );
  dp_1 \ANSWER/mem_reg[3][1][1]  ( .ip(n3771), .ck(clk), .q(
        \ANSWER/mem[3][1][1] ) );
  dp_1 \ANSWER/mem_reg[3][2][1]  ( .ip(n3770), .ck(clk), .q(
        \ANSWER/mem[3][2][1] ) );
  dp_1 \ANSWER/mem_reg[3][3][1]  ( .ip(n3769), .ck(clk), .q(
        \ANSWER/mem[3][3][1] ) );
  dp_1 \ANSWER/mem_reg[3][4][1]  ( .ip(n3768), .ck(clk), .q(
        \ANSWER/mem[3][4][1] ) );
  dp_1 \ANSWER/mem_reg[3][5][1]  ( .ip(n3767), .ck(clk), .q(
        \ANSWER/mem[3][5][1] ) );
  dp_1 \ANSWER/mem_reg[3][6][1]  ( .ip(n3766), .ck(clk), .q(
        \ANSWER/mem[3][6][1] ) );
  dp_1 \ANSWER/mem_reg[3][7][1]  ( .ip(n3765), .ck(clk), .q(
        \ANSWER/mem[3][7][1] ) );
  dp_1 \ANSWER/mem_reg[3][8][1]  ( .ip(n3764), .ck(clk), .q(
        \ANSWER/mem[3][8][1] ) );
  dp_1 \ANSWER/mem_reg[3][9][1]  ( .ip(n3763), .ck(clk), .q(
        \ANSWER/mem[3][9][1] ) );
  dp_1 \ANSWER/mem_reg[4][0][1]  ( .ip(n3762), .ck(clk), .q(
        \ANSWER/mem[4][0][1] ) );
  dp_1 \ANSWER/mem_reg[4][1][1]  ( .ip(n3761), .ck(clk), .q(
        \ANSWER/mem[4][1][1] ) );
  dp_1 \ANSWER/mem_reg[4][2][1]  ( .ip(n3760), .ck(clk), .q(
        \ANSWER/mem[4][2][1] ) );
  dp_1 \ANSWER/mem_reg[4][3][1]  ( .ip(n3759), .ck(clk), .q(
        \ANSWER/mem[4][3][1] ) );
  dp_1 \ANSWER/mem_reg[4][4][1]  ( .ip(n3758), .ck(clk), .q(
        \ANSWER/mem[4][4][1] ) );
  dp_1 \ANSWER/mem_reg[4][5][1]  ( .ip(n3757), .ck(clk), .q(
        \ANSWER/mem[4][5][1] ) );
  dp_1 \ANSWER/mem_reg[4][6][1]  ( .ip(n3756), .ck(clk), .q(
        \ANSWER/mem[4][6][1] ) );
  dp_1 \ANSWER/mem_reg[4][7][1]  ( .ip(n3755), .ck(clk), .q(
        \ANSWER/mem[4][7][1] ) );
  dp_1 \ANSWER/mem_reg[4][8][1]  ( .ip(n3754), .ck(clk), .q(
        \ANSWER/mem[4][8][1] ) );
  dp_1 \ANSWER/mem_reg[4][9][1]  ( .ip(n3753), .ck(clk), .q(
        \ANSWER/mem[4][9][1] ) );
  dp_1 \ANSWER/mem_reg[5][0][1]  ( .ip(n3752), .ck(clk), .q(
        \ANSWER/mem[5][0][1] ) );
  dp_1 \ANSWER/mem_reg[5][1][1]  ( .ip(n3751), .ck(clk), .q(
        \ANSWER/mem[5][1][1] ) );
  dp_1 \ANSWER/mem_reg[5][2][1]  ( .ip(n3750), .ck(clk), .q(
        \ANSWER/mem[5][2][1] ) );
  dp_1 \ANSWER/mem_reg[5][3][1]  ( .ip(n3749), .ck(clk), .q(
        \ANSWER/mem[5][3][1] ) );
  dp_1 \ANSWER/mem_reg[5][4][1]  ( .ip(n3748), .ck(clk), .q(
        \ANSWER/mem[5][4][1] ) );
  dp_1 \ANSWER/mem_reg[5][5][1]  ( .ip(n3747), .ck(clk), .q(
        \ANSWER/mem[5][5][1] ) );
  dp_1 \ANSWER/mem_reg[5][6][1]  ( .ip(n3746), .ck(clk), .q(
        \ANSWER/mem[5][6][1] ) );
  dp_1 \ANSWER/mem_reg[5][7][1]  ( .ip(n3745), .ck(clk), .q(
        \ANSWER/mem[5][7][1] ) );
  dp_1 \ANSWER/mem_reg[5][8][1]  ( .ip(n3744), .ck(clk), .q(
        \ANSWER/mem[5][8][1] ) );
  dp_1 \ANSWER/mem_reg[5][9][1]  ( .ip(n3743), .ck(clk), .q(
        \ANSWER/mem[5][9][1] ) );
  dp_1 \ANSWER/mem_reg[6][0][1]  ( .ip(n3742), .ck(clk), .q(
        \ANSWER/mem[6][0][1] ) );
  dp_1 \ANSWER/mem_reg[6][1][1]  ( .ip(n3741), .ck(clk), .q(
        \ANSWER/mem[6][1][1] ) );
  dp_1 \ANSWER/mem_reg[6][2][1]  ( .ip(n3740), .ck(clk), .q(
        \ANSWER/mem[6][2][1] ) );
  dp_1 \ANSWER/mem_reg[6][3][1]  ( .ip(n3739), .ck(clk), .q(
        \ANSWER/mem[6][3][1] ) );
  dp_1 \ANSWER/mem_reg[6][4][1]  ( .ip(n3738), .ck(clk), .q(
        \ANSWER/mem[6][4][1] ) );
  dp_1 \ANSWER/mem_reg[6][5][1]  ( .ip(n3737), .ck(clk), .q(
        \ANSWER/mem[6][5][1] ) );
  dp_1 \ANSWER/mem_reg[6][6][1]  ( .ip(n3736), .ck(clk), .q(
        \ANSWER/mem[6][6][1] ) );
  dp_1 \ANSWER/mem_reg[6][7][1]  ( .ip(n3735), .ck(clk), .q(
        \ANSWER/mem[6][7][1] ) );
  dp_1 \ANSWER/mem_reg[6][8][1]  ( .ip(n3734), .ck(clk), .q(
        \ANSWER/mem[6][8][1] ) );
  dp_1 \ANSWER/mem_reg[6][9][1]  ( .ip(n3733), .ck(clk), .q(
        \ANSWER/mem[6][9][1] ) );
  dp_1 \ANSWER/mem_reg[7][0][1]  ( .ip(n3732), .ck(clk), .q(
        \ANSWER/mem[7][0][1] ) );
  dp_1 \ANSWER/mem_reg[7][1][1]  ( .ip(n3731), .ck(clk), .q(
        \ANSWER/mem[7][1][1] ) );
  dp_1 \ANSWER/mem_reg[7][2][1]  ( .ip(n3730), .ck(clk), .q(
        \ANSWER/mem[7][2][1] ) );
  dp_1 \ANSWER/mem_reg[7][3][1]  ( .ip(n3729), .ck(clk), .q(
        \ANSWER/mem[7][3][1] ) );
  dp_1 \ANSWER/mem_reg[7][4][1]  ( .ip(n3728), .ck(clk), .q(
        \ANSWER/mem[7][4][1] ) );
  dp_1 \ANSWER/mem_reg[7][5][1]  ( .ip(n3727), .ck(clk), .q(
        \ANSWER/mem[7][5][1] ) );
  dp_1 \ANSWER/mem_reg[7][6][1]  ( .ip(n3726), .ck(clk), .q(
        \ANSWER/mem[7][6][1] ) );
  dp_1 \ANSWER/mem_reg[7][7][1]  ( .ip(n3725), .ck(clk), .q(
        \ANSWER/mem[7][7][1] ) );
  dp_1 \ANSWER/mem_reg[7][8][1]  ( .ip(n3724), .ck(clk), .q(
        \ANSWER/mem[7][8][1] ) );
  dp_1 \ANSWER/mem_reg[7][9][1]  ( .ip(n3723), .ck(clk), .q(
        \ANSWER/mem[7][9][1] ) );
  dp_1 \ANSWER/mem_reg[8][0][1]  ( .ip(n3722), .ck(clk), .q(
        \ANSWER/mem[8][0][1] ) );
  dp_1 \ANSWER/mem_reg[8][1][1]  ( .ip(n3721), .ck(clk), .q(
        \ANSWER/mem[8][1][1] ) );
  dp_1 \ANSWER/mem_reg[8][2][1]  ( .ip(n3720), .ck(clk), .q(
        \ANSWER/mem[8][2][1] ) );
  dp_1 \ANSWER/mem_reg[8][3][1]  ( .ip(n3719), .ck(clk), .q(
        \ANSWER/mem[8][3][1] ) );
  dp_1 \ANSWER/mem_reg[8][4][1]  ( .ip(n3718), .ck(clk), .q(
        \ANSWER/mem[8][4][1] ) );
  dp_1 \ANSWER/mem_reg[8][5][1]  ( .ip(n3717), .ck(clk), .q(
        \ANSWER/mem[8][5][1] ) );
  dp_1 \ANSWER/mem_reg[8][6][1]  ( .ip(n3716), .ck(clk), .q(
        \ANSWER/mem[8][6][1] ) );
  dp_1 \ANSWER/mem_reg[8][7][1]  ( .ip(n3715), .ck(clk), .q(
        \ANSWER/mem[8][7][1] ) );
  dp_1 \ANSWER/mem_reg[8][8][1]  ( .ip(n3714), .ck(clk), .q(
        \ANSWER/mem[8][8][1] ) );
  dp_1 \ANSWER/mem_reg[8][9][1]  ( .ip(n3713), .ck(clk), .q(
        \ANSWER/mem[8][9][1] ) );
  dp_1 \ANSWER/mem_reg[9][0][1]  ( .ip(n3712), .ck(clk), .q(
        \ANSWER/mem[9][0][1] ) );
  dp_1 \ANSWER/mem_reg[9][1][1]  ( .ip(n3711), .ck(clk), .q(
        \ANSWER/mem[9][1][1] ) );
  dp_1 \ANSWER/mem_reg[9][2][1]  ( .ip(n3710), .ck(clk), .q(
        \ANSWER/mem[9][2][1] ) );
  dp_1 \ANSWER/mem_reg[9][3][1]  ( .ip(n3709), .ck(clk), .q(
        \ANSWER/mem[9][3][1] ) );
  dp_1 \ANSWER/mem_reg[9][4][1]  ( .ip(n3708), .ck(clk), .q(
        \ANSWER/mem[9][4][1] ) );
  dp_1 \ANSWER/mem_reg[9][5][1]  ( .ip(n3707), .ck(clk), .q(
        \ANSWER/mem[9][5][1] ) );
  dp_1 \ANSWER/mem_reg[9][6][1]  ( .ip(n3706), .ck(clk), .q(
        \ANSWER/mem[9][6][1] ) );
  dp_1 \ANSWER/mem_reg[9][7][1]  ( .ip(n3705), .ck(clk), .q(
        \ANSWER/mem[9][7][1] ) );
  dp_1 \ANSWER/mem_reg[9][8][1]  ( .ip(n3704), .ck(clk), .q(
        \ANSWER/mem[9][8][1] ) );
  dp_1 \ANSWER/mem_reg[9][9][1]  ( .ip(n3703), .ck(clk), .q(
        \ANSWER/mem[9][9][1] ) );
  dp_1 \SIGMOID/lut_out_reg[2]  ( .ip(n3908), .ck(clk), .q(
        \SIGMOID/lut_out [2]) );
  dp_1 \ANSWER/mem_reg[0][0][2]  ( .ip(n3702), .ck(clk), .q(
        \ANSWER/mem[0][0][2] ) );
  dp_1 \ANSWER/mem_reg[0][1][2]  ( .ip(n3701), .ck(clk), .q(
        \ANSWER/mem[0][1][2] ) );
  dp_1 \ANSWER/mem_reg[0][2][2]  ( .ip(n3700), .ck(clk), .q(
        \ANSWER/mem[0][2][2] ) );
  dp_1 \ANSWER/mem_reg[0][3][2]  ( .ip(n3699), .ck(clk), .q(
        \ANSWER/mem[0][3][2] ) );
  dp_1 \ANSWER/mem_reg[0][4][2]  ( .ip(n3698), .ck(clk), .q(
        \ANSWER/mem[0][4][2] ) );
  dp_1 \ANSWER/mem_reg[0][5][2]  ( .ip(n3697), .ck(clk), .q(
        \ANSWER/mem[0][5][2] ) );
  dp_1 \ANSWER/mem_reg[0][6][2]  ( .ip(n3696), .ck(clk), .q(
        \ANSWER/mem[0][6][2] ) );
  dp_1 \ANSWER/mem_reg[0][7][2]  ( .ip(n3695), .ck(clk), .q(
        \ANSWER/mem[0][7][2] ) );
  dp_1 \ANSWER/mem_reg[0][8][2]  ( .ip(n3694), .ck(clk), .q(
        \ANSWER/mem[0][8][2] ) );
  dp_1 \ANSWER/mem_reg[0][9][2]  ( .ip(n3693), .ck(clk), .q(
        \ANSWER/mem[0][9][2] ) );
  dp_1 \ANSWER/mem_reg[1][0][2]  ( .ip(n3692), .ck(clk), .q(
        \ANSWER/mem[1][0][2] ) );
  dp_1 \ANSWER/mem_reg[1][1][2]  ( .ip(n3691), .ck(clk), .q(
        \ANSWER/mem[1][1][2] ) );
  dp_1 \ANSWER/mem_reg[1][2][2]  ( .ip(n3690), .ck(clk), .q(
        \ANSWER/mem[1][2][2] ) );
  dp_1 \ANSWER/mem_reg[1][3][2]  ( .ip(n3689), .ck(clk), .q(
        \ANSWER/mem[1][3][2] ) );
  dp_1 \ANSWER/mem_reg[1][4][2]  ( .ip(n3688), .ck(clk), .q(
        \ANSWER/mem[1][4][2] ) );
  dp_1 \ANSWER/mem_reg[1][5][2]  ( .ip(n3687), .ck(clk), .q(
        \ANSWER/mem[1][5][2] ) );
  dp_1 \ANSWER/mem_reg[1][6][2]  ( .ip(n3686), .ck(clk), .q(
        \ANSWER/mem[1][6][2] ) );
  dp_1 \ANSWER/mem_reg[1][7][2]  ( .ip(n3685), .ck(clk), .q(
        \ANSWER/mem[1][7][2] ) );
  dp_1 \ANSWER/mem_reg[1][8][2]  ( .ip(n3684), .ck(clk), .q(
        \ANSWER/mem[1][8][2] ) );
  dp_1 \ANSWER/mem_reg[1][9][2]  ( .ip(n3683), .ck(clk), .q(
        \ANSWER/mem[1][9][2] ) );
  dp_1 \ANSWER/mem_reg[2][0][2]  ( .ip(n3682), .ck(clk), .q(
        \ANSWER/mem[2][0][2] ) );
  dp_1 \ANSWER/mem_reg[2][1][2]  ( .ip(n3681), .ck(clk), .q(
        \ANSWER/mem[2][1][2] ) );
  dp_1 \ANSWER/mem_reg[2][2][2]  ( .ip(n3680), .ck(clk), .q(
        \ANSWER/mem[2][2][2] ) );
  dp_1 \ANSWER/mem_reg[2][3][2]  ( .ip(n3679), .ck(clk), .q(
        \ANSWER/mem[2][3][2] ) );
  dp_1 \ANSWER/mem_reg[2][4][2]  ( .ip(n3678), .ck(clk), .q(
        \ANSWER/mem[2][4][2] ) );
  dp_1 \ANSWER/mem_reg[2][5][2]  ( .ip(n3677), .ck(clk), .q(
        \ANSWER/mem[2][5][2] ) );
  dp_1 \ANSWER/mem_reg[2][6][2]  ( .ip(n3676), .ck(clk), .q(
        \ANSWER/mem[2][6][2] ) );
  dp_1 \ANSWER/mem_reg[2][7][2]  ( .ip(n3675), .ck(clk), .q(
        \ANSWER/mem[2][7][2] ) );
  dp_1 \ANSWER/mem_reg[2][8][2]  ( .ip(n3674), .ck(clk), .q(
        \ANSWER/mem[2][8][2] ) );
  dp_1 \ANSWER/mem_reg[2][9][2]  ( .ip(n3673), .ck(clk), .q(
        \ANSWER/mem[2][9][2] ) );
  dp_1 \ANSWER/mem_reg[3][0][2]  ( .ip(n3672), .ck(clk), .q(
        \ANSWER/mem[3][0][2] ) );
  dp_1 \ANSWER/mem_reg[3][1][2]  ( .ip(n3671), .ck(clk), .q(
        \ANSWER/mem[3][1][2] ) );
  dp_1 \ANSWER/mem_reg[3][2][2]  ( .ip(n3670), .ck(clk), .q(
        \ANSWER/mem[3][2][2] ) );
  dp_1 \ANSWER/mem_reg[3][3][2]  ( .ip(n3669), .ck(clk), .q(
        \ANSWER/mem[3][3][2] ) );
  dp_1 \ANSWER/mem_reg[3][4][2]  ( .ip(n3668), .ck(clk), .q(
        \ANSWER/mem[3][4][2] ) );
  dp_1 \ANSWER/mem_reg[3][5][2]  ( .ip(n3667), .ck(clk), .q(
        \ANSWER/mem[3][5][2] ) );
  dp_1 \ANSWER/mem_reg[3][6][2]  ( .ip(n3666), .ck(clk), .q(
        \ANSWER/mem[3][6][2] ) );
  dp_1 \ANSWER/mem_reg[3][7][2]  ( .ip(n3665), .ck(clk), .q(
        \ANSWER/mem[3][7][2] ) );
  dp_1 \ANSWER/mem_reg[3][8][2]  ( .ip(n3664), .ck(clk), .q(
        \ANSWER/mem[3][8][2] ) );
  dp_1 \ANSWER/mem_reg[3][9][2]  ( .ip(n3663), .ck(clk), .q(
        \ANSWER/mem[3][9][2] ) );
  dp_1 \ANSWER/mem_reg[4][0][2]  ( .ip(n3662), .ck(clk), .q(
        \ANSWER/mem[4][0][2] ) );
  dp_1 \ANSWER/mem_reg[4][1][2]  ( .ip(n3661), .ck(clk), .q(
        \ANSWER/mem[4][1][2] ) );
  dp_1 \ANSWER/mem_reg[4][2][2]  ( .ip(n3660), .ck(clk), .q(
        \ANSWER/mem[4][2][2] ) );
  dp_1 \ANSWER/mem_reg[4][3][2]  ( .ip(n3659), .ck(clk), .q(
        \ANSWER/mem[4][3][2] ) );
  dp_1 \ANSWER/mem_reg[4][4][2]  ( .ip(n3658), .ck(clk), .q(
        \ANSWER/mem[4][4][2] ) );
  dp_1 \ANSWER/mem_reg[4][5][2]  ( .ip(n3657), .ck(clk), .q(
        \ANSWER/mem[4][5][2] ) );
  dp_1 \ANSWER/mem_reg[4][6][2]  ( .ip(n3656), .ck(clk), .q(
        \ANSWER/mem[4][6][2] ) );
  dp_1 \ANSWER/mem_reg[4][7][2]  ( .ip(n3655), .ck(clk), .q(
        \ANSWER/mem[4][7][2] ) );
  dp_1 \ANSWER/mem_reg[4][8][2]  ( .ip(n3654), .ck(clk), .q(
        \ANSWER/mem[4][8][2] ) );
  dp_1 \ANSWER/mem_reg[4][9][2]  ( .ip(n3653), .ck(clk), .q(
        \ANSWER/mem[4][9][2] ) );
  dp_1 \ANSWER/mem_reg[5][0][2]  ( .ip(n3652), .ck(clk), .q(
        \ANSWER/mem[5][0][2] ) );
  dp_1 \ANSWER/mem_reg[5][1][2]  ( .ip(n3651), .ck(clk), .q(
        \ANSWER/mem[5][1][2] ) );
  dp_1 \ANSWER/mem_reg[5][2][2]  ( .ip(n3650), .ck(clk), .q(
        \ANSWER/mem[5][2][2] ) );
  dp_1 \ANSWER/mem_reg[5][3][2]  ( .ip(n3649), .ck(clk), .q(
        \ANSWER/mem[5][3][2] ) );
  dp_1 \ANSWER/mem_reg[5][4][2]  ( .ip(n3648), .ck(clk), .q(
        \ANSWER/mem[5][4][2] ) );
  dp_1 \ANSWER/mem_reg[5][5][2]  ( .ip(n3647), .ck(clk), .q(
        \ANSWER/mem[5][5][2] ) );
  dp_1 \ANSWER/mem_reg[5][6][2]  ( .ip(n3646), .ck(clk), .q(
        \ANSWER/mem[5][6][2] ) );
  dp_1 \ANSWER/mem_reg[5][7][2]  ( .ip(n3645), .ck(clk), .q(
        \ANSWER/mem[5][7][2] ) );
  dp_1 \ANSWER/mem_reg[5][8][2]  ( .ip(n3644), .ck(clk), .q(
        \ANSWER/mem[5][8][2] ) );
  dp_1 \ANSWER/mem_reg[5][9][2]  ( .ip(n3643), .ck(clk), .q(
        \ANSWER/mem[5][9][2] ) );
  dp_1 \ANSWER/mem_reg[6][0][2]  ( .ip(n3642), .ck(clk), .q(
        \ANSWER/mem[6][0][2] ) );
  dp_1 \ANSWER/mem_reg[6][1][2]  ( .ip(n3641), .ck(clk), .q(
        \ANSWER/mem[6][1][2] ) );
  dp_1 \ANSWER/mem_reg[6][2][2]  ( .ip(n3640), .ck(clk), .q(
        \ANSWER/mem[6][2][2] ) );
  dp_1 \ANSWER/mem_reg[6][3][2]  ( .ip(n3639), .ck(clk), .q(
        \ANSWER/mem[6][3][2] ) );
  dp_1 \ANSWER/mem_reg[6][4][2]  ( .ip(n3638), .ck(clk), .q(
        \ANSWER/mem[6][4][2] ) );
  dp_1 \ANSWER/mem_reg[6][5][2]  ( .ip(n3637), .ck(clk), .q(
        \ANSWER/mem[6][5][2] ) );
  dp_1 \ANSWER/mem_reg[6][6][2]  ( .ip(n3636), .ck(clk), .q(
        \ANSWER/mem[6][6][2] ) );
  dp_1 \ANSWER/mem_reg[6][7][2]  ( .ip(n3635), .ck(clk), .q(
        \ANSWER/mem[6][7][2] ) );
  dp_1 \ANSWER/mem_reg[6][8][2]  ( .ip(n3634), .ck(clk), .q(
        \ANSWER/mem[6][8][2] ) );
  dp_1 \ANSWER/mem_reg[6][9][2]  ( .ip(n3633), .ck(clk), .q(
        \ANSWER/mem[6][9][2] ) );
  dp_1 \ANSWER/mem_reg[7][0][2]  ( .ip(n3632), .ck(clk), .q(
        \ANSWER/mem[7][0][2] ) );
  dp_1 \ANSWER/mem_reg[7][1][2]  ( .ip(n3631), .ck(clk), .q(
        \ANSWER/mem[7][1][2] ) );
  dp_1 \ANSWER/mem_reg[7][2][2]  ( .ip(n3630), .ck(clk), .q(
        \ANSWER/mem[7][2][2] ) );
  dp_1 \ANSWER/mem_reg[7][3][2]  ( .ip(n3629), .ck(clk), .q(
        \ANSWER/mem[7][3][2] ) );
  dp_1 \ANSWER/mem_reg[7][4][2]  ( .ip(n3628), .ck(clk), .q(
        \ANSWER/mem[7][4][2] ) );
  dp_1 \ANSWER/mem_reg[7][5][2]  ( .ip(n3627), .ck(clk), .q(
        \ANSWER/mem[7][5][2] ) );
  dp_1 \ANSWER/mem_reg[7][6][2]  ( .ip(n3626), .ck(clk), .q(
        \ANSWER/mem[7][6][2] ) );
  dp_1 \ANSWER/mem_reg[7][7][2]  ( .ip(n3625), .ck(clk), .q(
        \ANSWER/mem[7][7][2] ) );
  dp_1 \ANSWER/mem_reg[7][8][2]  ( .ip(n3624), .ck(clk), .q(
        \ANSWER/mem[7][8][2] ) );
  dp_1 \ANSWER/mem_reg[7][9][2]  ( .ip(n3623), .ck(clk), .q(
        \ANSWER/mem[7][9][2] ) );
  dp_1 \ANSWER/mem_reg[8][0][2]  ( .ip(n3622), .ck(clk), .q(
        \ANSWER/mem[8][0][2] ) );
  dp_1 \ANSWER/mem_reg[8][1][2]  ( .ip(n3621), .ck(clk), .q(
        \ANSWER/mem[8][1][2] ) );
  dp_1 \ANSWER/mem_reg[8][2][2]  ( .ip(n3620), .ck(clk), .q(
        \ANSWER/mem[8][2][2] ) );
  dp_1 \ANSWER/mem_reg[8][3][2]  ( .ip(n3619), .ck(clk), .q(
        \ANSWER/mem[8][3][2] ) );
  dp_1 \ANSWER/mem_reg[8][4][2]  ( .ip(n3618), .ck(clk), .q(
        \ANSWER/mem[8][4][2] ) );
  dp_1 \ANSWER/mem_reg[8][5][2]  ( .ip(n3617), .ck(clk), .q(
        \ANSWER/mem[8][5][2] ) );
  dp_1 \ANSWER/mem_reg[8][6][2]  ( .ip(n3616), .ck(clk), .q(
        \ANSWER/mem[8][6][2] ) );
  dp_1 \ANSWER/mem_reg[8][7][2]  ( .ip(n3615), .ck(clk), .q(
        \ANSWER/mem[8][7][2] ) );
  dp_1 \ANSWER/mem_reg[8][8][2]  ( .ip(n3614), .ck(clk), .q(
        \ANSWER/mem[8][8][2] ) );
  dp_1 \ANSWER/mem_reg[8][9][2]  ( .ip(n3613), .ck(clk), .q(
        \ANSWER/mem[8][9][2] ) );
  dp_1 \ANSWER/mem_reg[9][0][2]  ( .ip(n3612), .ck(clk), .q(
        \ANSWER/mem[9][0][2] ) );
  dp_1 \ANSWER/mem_reg[9][1][2]  ( .ip(n3611), .ck(clk), .q(
        \ANSWER/mem[9][1][2] ) );
  dp_1 \ANSWER/mem_reg[9][2][2]  ( .ip(n3610), .ck(clk), .q(
        \ANSWER/mem[9][2][2] ) );
  dp_1 \ANSWER/mem_reg[9][3][2]  ( .ip(n3609), .ck(clk), .q(
        \ANSWER/mem[9][3][2] ) );
  dp_1 \ANSWER/mem_reg[9][4][2]  ( .ip(n3608), .ck(clk), .q(
        \ANSWER/mem[9][4][2] ) );
  dp_1 \ANSWER/mem_reg[9][5][2]  ( .ip(n3607), .ck(clk), .q(
        \ANSWER/mem[9][5][2] ) );
  dp_1 \ANSWER/mem_reg[9][6][2]  ( .ip(n3606), .ck(clk), .q(
        \ANSWER/mem[9][6][2] ) );
  dp_1 \ANSWER/mem_reg[9][7][2]  ( .ip(n3605), .ck(clk), .q(
        \ANSWER/mem[9][7][2] ) );
  dp_1 \ANSWER/mem_reg[9][8][2]  ( .ip(n3604), .ck(clk), .q(
        \ANSWER/mem[9][8][2] ) );
  dp_1 \ANSWER/mem_reg[9][9][2]  ( .ip(n3603), .ck(clk), .q(
        \ANSWER/mem[9][9][2] ) );
  dp_1 \SIGMOID/lut_out_reg[3]  ( .ip(n3907), .ck(clk), .q(
        \SIGMOID/lut_out [3]) );
  dp_1 \ANSWER/mem_reg[0][0][3]  ( .ip(n3602), .ck(clk), .q(
        \ANSWER/mem[0][0][3] ) );
  dp_1 \ANSWER/mem_reg[0][1][3]  ( .ip(n3601), .ck(clk), .q(
        \ANSWER/mem[0][1][3] ) );
  dp_1 \ANSWER/mem_reg[0][2][3]  ( .ip(n3600), .ck(clk), .q(
        \ANSWER/mem[0][2][3] ) );
  dp_1 \ANSWER/mem_reg[0][3][3]  ( .ip(n3599), .ck(clk), .q(
        \ANSWER/mem[0][3][3] ) );
  dp_1 \ANSWER/mem_reg[0][4][3]  ( .ip(n3598), .ck(clk), .q(
        \ANSWER/mem[0][4][3] ) );
  dp_1 \ANSWER/mem_reg[0][5][3]  ( .ip(n3597), .ck(clk), .q(
        \ANSWER/mem[0][5][3] ) );
  dp_1 \ANSWER/mem_reg[0][6][3]  ( .ip(n3596), .ck(clk), .q(
        \ANSWER/mem[0][6][3] ) );
  dp_1 \ANSWER/mem_reg[0][7][3]  ( .ip(n3595), .ck(clk), .q(
        \ANSWER/mem[0][7][3] ) );
  dp_1 \ANSWER/mem_reg[0][8][3]  ( .ip(n3594), .ck(clk), .q(
        \ANSWER/mem[0][8][3] ) );
  dp_1 \ANSWER/mem_reg[0][9][3]  ( .ip(n3593), .ck(clk), .q(
        \ANSWER/mem[0][9][3] ) );
  dp_1 \ANSWER/mem_reg[1][0][3]  ( .ip(n3592), .ck(clk), .q(
        \ANSWER/mem[1][0][3] ) );
  dp_1 \ANSWER/mem_reg[1][1][3]  ( .ip(n3591), .ck(clk), .q(
        \ANSWER/mem[1][1][3] ) );
  dp_1 \ANSWER/mem_reg[1][2][3]  ( .ip(n3590), .ck(clk), .q(
        \ANSWER/mem[1][2][3] ) );
  dp_1 \ANSWER/mem_reg[1][3][3]  ( .ip(n3589), .ck(clk), .q(
        \ANSWER/mem[1][3][3] ) );
  dp_1 \ANSWER/mem_reg[1][4][3]  ( .ip(n3588), .ck(clk), .q(
        \ANSWER/mem[1][4][3] ) );
  dp_1 \ANSWER/mem_reg[1][5][3]  ( .ip(n3587), .ck(clk), .q(
        \ANSWER/mem[1][5][3] ) );
  dp_1 \ANSWER/mem_reg[1][6][3]  ( .ip(n3586), .ck(clk), .q(
        \ANSWER/mem[1][6][3] ) );
  dp_1 \ANSWER/mem_reg[1][7][3]  ( .ip(n3585), .ck(clk), .q(
        \ANSWER/mem[1][7][3] ) );
  dp_1 \ANSWER/mem_reg[1][8][3]  ( .ip(n3584), .ck(clk), .q(
        \ANSWER/mem[1][8][3] ) );
  dp_1 \ANSWER/mem_reg[1][9][3]  ( .ip(n3583), .ck(clk), .q(
        \ANSWER/mem[1][9][3] ) );
  dp_1 \ANSWER/mem_reg[2][0][3]  ( .ip(n3582), .ck(clk), .q(
        \ANSWER/mem[2][0][3] ) );
  dp_1 \ANSWER/mem_reg[2][1][3]  ( .ip(n3581), .ck(clk), .q(
        \ANSWER/mem[2][1][3] ) );
  dp_1 \ANSWER/mem_reg[2][2][3]  ( .ip(n3580), .ck(clk), .q(
        \ANSWER/mem[2][2][3] ) );
  dp_1 \ANSWER/mem_reg[2][3][3]  ( .ip(n3579), .ck(clk), .q(
        \ANSWER/mem[2][3][3] ) );
  dp_1 \ANSWER/mem_reg[2][4][3]  ( .ip(n3578), .ck(clk), .q(
        \ANSWER/mem[2][4][3] ) );
  dp_1 \ANSWER/mem_reg[2][5][3]  ( .ip(n3577), .ck(clk), .q(
        \ANSWER/mem[2][5][3] ) );
  dp_1 \ANSWER/mem_reg[2][6][3]  ( .ip(n3576), .ck(clk), .q(
        \ANSWER/mem[2][6][3] ) );
  dp_1 \ANSWER/mem_reg[2][7][3]  ( .ip(n3575), .ck(clk), .q(
        \ANSWER/mem[2][7][3] ) );
  dp_1 \ANSWER/mem_reg[2][8][3]  ( .ip(n3574), .ck(clk), .q(
        \ANSWER/mem[2][8][3] ) );
  dp_1 \ANSWER/mem_reg[2][9][3]  ( .ip(n3573), .ck(clk), .q(
        \ANSWER/mem[2][9][3] ) );
  dp_1 \ANSWER/mem_reg[3][0][3]  ( .ip(n3572), .ck(clk), .q(
        \ANSWER/mem[3][0][3] ) );
  dp_1 \ANSWER/mem_reg[3][1][3]  ( .ip(n3571), .ck(clk), .q(
        \ANSWER/mem[3][1][3] ) );
  dp_1 \ANSWER/mem_reg[3][2][3]  ( .ip(n3570), .ck(clk), .q(
        \ANSWER/mem[3][2][3] ) );
  dp_1 \ANSWER/mem_reg[3][3][3]  ( .ip(n3569), .ck(clk), .q(
        \ANSWER/mem[3][3][3] ) );
  dp_1 \ANSWER/mem_reg[3][4][3]  ( .ip(n3568), .ck(clk), .q(
        \ANSWER/mem[3][4][3] ) );
  dp_1 \ANSWER/mem_reg[3][5][3]  ( .ip(n3567), .ck(clk), .q(
        \ANSWER/mem[3][5][3] ) );
  dp_1 \ANSWER/mem_reg[3][6][3]  ( .ip(n3566), .ck(clk), .q(
        \ANSWER/mem[3][6][3] ) );
  dp_1 \ANSWER/mem_reg[3][7][3]  ( .ip(n3565), .ck(clk), .q(
        \ANSWER/mem[3][7][3] ) );
  dp_1 \ANSWER/mem_reg[3][8][3]  ( .ip(n3564), .ck(clk), .q(
        \ANSWER/mem[3][8][3] ) );
  dp_1 \ANSWER/mem_reg[3][9][3]  ( .ip(n3563), .ck(clk), .q(
        \ANSWER/mem[3][9][3] ) );
  dp_1 \ANSWER/mem_reg[4][0][3]  ( .ip(n3562), .ck(clk), .q(
        \ANSWER/mem[4][0][3] ) );
  dp_1 \ANSWER/mem_reg[4][1][3]  ( .ip(n3561), .ck(clk), .q(
        \ANSWER/mem[4][1][3] ) );
  dp_1 \ANSWER/mem_reg[4][2][3]  ( .ip(n3560), .ck(clk), .q(
        \ANSWER/mem[4][2][3] ) );
  dp_1 \ANSWER/mem_reg[4][3][3]  ( .ip(n3559), .ck(clk), .q(
        \ANSWER/mem[4][3][3] ) );
  dp_1 \ANSWER/mem_reg[4][4][3]  ( .ip(n3558), .ck(clk), .q(
        \ANSWER/mem[4][4][3] ) );
  dp_1 \ANSWER/mem_reg[4][5][3]  ( .ip(n3557), .ck(clk), .q(
        \ANSWER/mem[4][5][3] ) );
  dp_1 \ANSWER/mem_reg[4][6][3]  ( .ip(n3556), .ck(clk), .q(
        \ANSWER/mem[4][6][3] ) );
  dp_1 \ANSWER/mem_reg[4][7][3]  ( .ip(n3555), .ck(clk), .q(
        \ANSWER/mem[4][7][3] ) );
  dp_1 \ANSWER/mem_reg[4][8][3]  ( .ip(n3554), .ck(clk), .q(
        \ANSWER/mem[4][8][3] ) );
  dp_1 \ANSWER/mem_reg[4][9][3]  ( .ip(n3553), .ck(clk), .q(
        \ANSWER/mem[4][9][3] ) );
  dp_1 \ANSWER/mem_reg[5][0][3]  ( .ip(n3552), .ck(clk), .q(
        \ANSWER/mem[5][0][3] ) );
  dp_1 \ANSWER/mem_reg[5][1][3]  ( .ip(n3551), .ck(clk), .q(
        \ANSWER/mem[5][1][3] ) );
  dp_1 \ANSWER/mem_reg[5][2][3]  ( .ip(n3550), .ck(clk), .q(
        \ANSWER/mem[5][2][3] ) );
  dp_1 \ANSWER/mem_reg[5][3][3]  ( .ip(n3549), .ck(clk), .q(
        \ANSWER/mem[5][3][3] ) );
  dp_1 \ANSWER/mem_reg[5][4][3]  ( .ip(n3548), .ck(clk), .q(
        \ANSWER/mem[5][4][3] ) );
  dp_1 \ANSWER/mem_reg[5][5][3]  ( .ip(n3547), .ck(clk), .q(
        \ANSWER/mem[5][5][3] ) );
  dp_1 \ANSWER/mem_reg[5][6][3]  ( .ip(n3546), .ck(clk), .q(
        \ANSWER/mem[5][6][3] ) );
  dp_1 \ANSWER/mem_reg[5][7][3]  ( .ip(n3545), .ck(clk), .q(
        \ANSWER/mem[5][7][3] ) );
  dp_1 \ANSWER/mem_reg[5][8][3]  ( .ip(n3544), .ck(clk), .q(
        \ANSWER/mem[5][8][3] ) );
  dp_1 \ANSWER/mem_reg[5][9][3]  ( .ip(n3543), .ck(clk), .q(
        \ANSWER/mem[5][9][3] ) );
  dp_1 \ANSWER/mem_reg[6][0][3]  ( .ip(n3542), .ck(clk), .q(
        \ANSWER/mem[6][0][3] ) );
  dp_1 \ANSWER/mem_reg[6][1][3]  ( .ip(n3541), .ck(clk), .q(
        \ANSWER/mem[6][1][3] ) );
  dp_1 \ANSWER/mem_reg[6][2][3]  ( .ip(n3540), .ck(clk), .q(
        \ANSWER/mem[6][2][3] ) );
  dp_1 \ANSWER/mem_reg[6][3][3]  ( .ip(n3539), .ck(clk), .q(
        \ANSWER/mem[6][3][3] ) );
  dp_1 \ANSWER/mem_reg[6][4][3]  ( .ip(n3538), .ck(clk), .q(
        \ANSWER/mem[6][4][3] ) );
  dp_1 \ANSWER/mem_reg[6][5][3]  ( .ip(n3537), .ck(clk), .q(
        \ANSWER/mem[6][5][3] ) );
  dp_1 \ANSWER/mem_reg[6][6][3]  ( .ip(n3536), .ck(clk), .q(
        \ANSWER/mem[6][6][3] ) );
  dp_1 \ANSWER/mem_reg[6][7][3]  ( .ip(n3535), .ck(clk), .q(
        \ANSWER/mem[6][7][3] ) );
  dp_1 \ANSWER/mem_reg[6][8][3]  ( .ip(n3534), .ck(clk), .q(
        \ANSWER/mem[6][8][3] ) );
  dp_1 \ANSWER/mem_reg[6][9][3]  ( .ip(n3533), .ck(clk), .q(
        \ANSWER/mem[6][9][3] ) );
  dp_1 \ANSWER/mem_reg[7][0][3]  ( .ip(n3532), .ck(clk), .q(
        \ANSWER/mem[7][0][3] ) );
  dp_1 \ANSWER/mem_reg[7][1][3]  ( .ip(n3531), .ck(clk), .q(
        \ANSWER/mem[7][1][3] ) );
  dp_1 \ANSWER/mem_reg[7][2][3]  ( .ip(n3530), .ck(clk), .q(
        \ANSWER/mem[7][2][3] ) );
  dp_1 \ANSWER/mem_reg[7][3][3]  ( .ip(n3529), .ck(clk), .q(
        \ANSWER/mem[7][3][3] ) );
  dp_1 \ANSWER/mem_reg[7][4][3]  ( .ip(n3528), .ck(clk), .q(
        \ANSWER/mem[7][4][3] ) );
  dp_1 \ANSWER/mem_reg[7][5][3]  ( .ip(n3527), .ck(clk), .q(
        \ANSWER/mem[7][5][3] ) );
  dp_1 \ANSWER/mem_reg[7][6][3]  ( .ip(n3526), .ck(clk), .q(
        \ANSWER/mem[7][6][3] ) );
  dp_1 \ANSWER/mem_reg[7][7][3]  ( .ip(n3525), .ck(clk), .q(
        \ANSWER/mem[7][7][3] ) );
  dp_1 \ANSWER/mem_reg[7][8][3]  ( .ip(n3524), .ck(clk), .q(
        \ANSWER/mem[7][8][3] ) );
  dp_1 \ANSWER/mem_reg[7][9][3]  ( .ip(n3523), .ck(clk), .q(
        \ANSWER/mem[7][9][3] ) );
  dp_1 \ANSWER/mem_reg[8][0][3]  ( .ip(n3522), .ck(clk), .q(
        \ANSWER/mem[8][0][3] ) );
  dp_1 \ANSWER/mem_reg[8][1][3]  ( .ip(n3521), .ck(clk), .q(
        \ANSWER/mem[8][1][3] ) );
  dp_1 \ANSWER/mem_reg[8][2][3]  ( .ip(n3520), .ck(clk), .q(
        \ANSWER/mem[8][2][3] ) );
  dp_1 \ANSWER/mem_reg[8][3][3]  ( .ip(n3519), .ck(clk), .q(
        \ANSWER/mem[8][3][3] ) );
  dp_1 \ANSWER/mem_reg[8][4][3]  ( .ip(n3518), .ck(clk), .q(
        \ANSWER/mem[8][4][3] ) );
  dp_1 \ANSWER/mem_reg[8][5][3]  ( .ip(n3517), .ck(clk), .q(
        \ANSWER/mem[8][5][3] ) );
  dp_1 \ANSWER/mem_reg[8][6][3]  ( .ip(n3516), .ck(clk), .q(
        \ANSWER/mem[8][6][3] ) );
  dp_1 \ANSWER/mem_reg[8][7][3]  ( .ip(n3515), .ck(clk), .q(
        \ANSWER/mem[8][7][3] ) );
  dp_1 \ANSWER/mem_reg[8][8][3]  ( .ip(n3514), .ck(clk), .q(
        \ANSWER/mem[8][8][3] ) );
  dp_1 \ANSWER/mem_reg[8][9][3]  ( .ip(n3513), .ck(clk), .q(
        \ANSWER/mem[8][9][3] ) );
  dp_1 \ANSWER/mem_reg[9][0][3]  ( .ip(n3512), .ck(clk), .q(
        \ANSWER/mem[9][0][3] ) );
  dp_1 \ANSWER/mem_reg[9][1][3]  ( .ip(n3511), .ck(clk), .q(
        \ANSWER/mem[9][1][3] ) );
  dp_1 \ANSWER/mem_reg[9][2][3]  ( .ip(n3510), .ck(clk), .q(
        \ANSWER/mem[9][2][3] ) );
  dp_1 \ANSWER/mem_reg[9][3][3]  ( .ip(n3509), .ck(clk), .q(
        \ANSWER/mem[9][3][3] ) );
  dp_1 \ANSWER/mem_reg[9][4][3]  ( .ip(n3508), .ck(clk), .q(
        \ANSWER/mem[9][4][3] ) );
  dp_1 \ANSWER/mem_reg[9][5][3]  ( .ip(n3507), .ck(clk), .q(
        \ANSWER/mem[9][5][3] ) );
  dp_1 \ANSWER/mem_reg[9][6][3]  ( .ip(n3506), .ck(clk), .q(
        \ANSWER/mem[9][6][3] ) );
  dp_1 \ANSWER/mem_reg[9][7][3]  ( .ip(n3505), .ck(clk), .q(
        \ANSWER/mem[9][7][3] ) );
  dp_1 \ANSWER/mem_reg[9][8][3]  ( .ip(n3504), .ck(clk), .q(
        \ANSWER/mem[9][8][3] ) );
  dp_1 \ANSWER/mem_reg[9][9][3]  ( .ip(n3503), .ck(clk), .q(
        \ANSWER/mem[9][9][3] ) );
  dp_1 \SIGMOID/lut_out_reg[4]  ( .ip(n3906), .ck(clk), .q(
        \SIGMOID/lut_out [4]) );
  dp_1 \ANSWER/mem_reg[0][0][4]  ( .ip(n3502), .ck(clk), .q(
        \ANSWER/mem[0][0][4] ) );
  dp_1 \ANSWER/mem_reg[0][1][4]  ( .ip(n3501), .ck(clk), .q(
        \ANSWER/mem[0][1][4] ) );
  dp_1 \ANSWER/mem_reg[0][2][4]  ( .ip(n3500), .ck(clk), .q(
        \ANSWER/mem[0][2][4] ) );
  dp_1 \ANSWER/mem_reg[0][3][4]  ( .ip(n3499), .ck(clk), .q(
        \ANSWER/mem[0][3][4] ) );
  dp_1 \ANSWER/mem_reg[0][4][4]  ( .ip(n3498), .ck(clk), .q(
        \ANSWER/mem[0][4][4] ) );
  dp_1 \ANSWER/mem_reg[0][5][4]  ( .ip(n3497), .ck(clk), .q(
        \ANSWER/mem[0][5][4] ) );
  dp_1 \ANSWER/mem_reg[0][6][4]  ( .ip(n3496), .ck(clk), .q(
        \ANSWER/mem[0][6][4] ) );
  dp_1 \ANSWER/mem_reg[0][7][4]  ( .ip(n3495), .ck(clk), .q(
        \ANSWER/mem[0][7][4] ) );
  dp_1 \ANSWER/mem_reg[0][8][4]  ( .ip(n3494), .ck(clk), .q(
        \ANSWER/mem[0][8][4] ) );
  dp_1 \ANSWER/mem_reg[0][9][4]  ( .ip(n3493), .ck(clk), .q(
        \ANSWER/mem[0][9][4] ) );
  dp_1 \ANSWER/mem_reg[1][0][4]  ( .ip(n3492), .ck(clk), .q(
        \ANSWER/mem[1][0][4] ) );
  dp_1 \ANSWER/mem_reg[1][1][4]  ( .ip(n3491), .ck(clk), .q(
        \ANSWER/mem[1][1][4] ) );
  dp_1 \ANSWER/mem_reg[1][2][4]  ( .ip(n3490), .ck(clk), .q(
        \ANSWER/mem[1][2][4] ) );
  dp_1 \ANSWER/mem_reg[1][3][4]  ( .ip(n3489), .ck(clk), .q(
        \ANSWER/mem[1][3][4] ) );
  dp_1 \ANSWER/mem_reg[1][4][4]  ( .ip(n3488), .ck(clk), .q(
        \ANSWER/mem[1][4][4] ) );
  dp_1 \ANSWER/mem_reg[1][5][4]  ( .ip(n3487), .ck(clk), .q(
        \ANSWER/mem[1][5][4] ) );
  dp_1 \ANSWER/mem_reg[1][6][4]  ( .ip(n3486), .ck(clk), .q(
        \ANSWER/mem[1][6][4] ) );
  dp_1 \ANSWER/mem_reg[1][7][4]  ( .ip(n3485), .ck(clk), .q(
        \ANSWER/mem[1][7][4] ) );
  dp_1 \ANSWER/mem_reg[1][8][4]  ( .ip(n3484), .ck(clk), .q(
        \ANSWER/mem[1][8][4] ) );
  dp_1 \ANSWER/mem_reg[1][9][4]  ( .ip(n3483), .ck(clk), .q(
        \ANSWER/mem[1][9][4] ) );
  dp_1 \ANSWER/mem_reg[2][0][4]  ( .ip(n3482), .ck(clk), .q(
        \ANSWER/mem[2][0][4] ) );
  dp_1 \ANSWER/mem_reg[2][1][4]  ( .ip(n3481), .ck(clk), .q(
        \ANSWER/mem[2][1][4] ) );
  dp_1 \ANSWER/mem_reg[2][2][4]  ( .ip(n3480), .ck(clk), .q(
        \ANSWER/mem[2][2][4] ) );
  dp_1 \ANSWER/mem_reg[2][3][4]  ( .ip(n3479), .ck(clk), .q(
        \ANSWER/mem[2][3][4] ) );
  dp_1 \ANSWER/mem_reg[2][4][4]  ( .ip(n3478), .ck(clk), .q(
        \ANSWER/mem[2][4][4] ) );
  dp_1 \ANSWER/mem_reg[2][5][4]  ( .ip(n3477), .ck(clk), .q(
        \ANSWER/mem[2][5][4] ) );
  dp_1 \ANSWER/mem_reg[2][6][4]  ( .ip(n3476), .ck(clk), .q(
        \ANSWER/mem[2][6][4] ) );
  dp_1 \ANSWER/mem_reg[2][7][4]  ( .ip(n3475), .ck(clk), .q(
        \ANSWER/mem[2][7][4] ) );
  dp_1 \ANSWER/mem_reg[2][8][4]  ( .ip(n3474), .ck(clk), .q(
        \ANSWER/mem[2][8][4] ) );
  dp_1 \ANSWER/mem_reg[2][9][4]  ( .ip(n3473), .ck(clk), .q(
        \ANSWER/mem[2][9][4] ) );
  dp_1 \ANSWER/mem_reg[3][0][4]  ( .ip(n3472), .ck(clk), .q(
        \ANSWER/mem[3][0][4] ) );
  dp_1 \ANSWER/mem_reg[3][1][4]  ( .ip(n3471), .ck(clk), .q(
        \ANSWER/mem[3][1][4] ) );
  dp_1 \ANSWER/mem_reg[3][2][4]  ( .ip(n3470), .ck(clk), .q(
        \ANSWER/mem[3][2][4] ) );
  dp_1 \ANSWER/mem_reg[3][3][4]  ( .ip(n3469), .ck(clk), .q(
        \ANSWER/mem[3][3][4] ) );
  dp_1 \ANSWER/mem_reg[3][4][4]  ( .ip(n3468), .ck(clk), .q(
        \ANSWER/mem[3][4][4] ) );
  dp_1 \ANSWER/mem_reg[3][5][4]  ( .ip(n3467), .ck(clk), .q(
        \ANSWER/mem[3][5][4] ) );
  dp_1 \ANSWER/mem_reg[3][6][4]  ( .ip(n3466), .ck(clk), .q(
        \ANSWER/mem[3][6][4] ) );
  dp_1 \ANSWER/mem_reg[3][7][4]  ( .ip(n3465), .ck(clk), .q(
        \ANSWER/mem[3][7][4] ) );
  dp_1 \ANSWER/mem_reg[3][8][4]  ( .ip(n3464), .ck(clk), .q(
        \ANSWER/mem[3][8][4] ) );
  dp_1 \ANSWER/mem_reg[3][9][4]  ( .ip(n3463), .ck(clk), .q(
        \ANSWER/mem[3][9][4] ) );
  dp_1 \ANSWER/mem_reg[4][0][4]  ( .ip(n3462), .ck(clk), .q(
        \ANSWER/mem[4][0][4] ) );
  dp_1 \ANSWER/mem_reg[4][1][4]  ( .ip(n3461), .ck(clk), .q(
        \ANSWER/mem[4][1][4] ) );
  dp_1 \ANSWER/mem_reg[4][2][4]  ( .ip(n3460), .ck(clk), .q(
        \ANSWER/mem[4][2][4] ) );
  dp_1 \ANSWER/mem_reg[4][3][4]  ( .ip(n3459), .ck(clk), .q(
        \ANSWER/mem[4][3][4] ) );
  dp_1 \ANSWER/mem_reg[4][4][4]  ( .ip(n3458), .ck(clk), .q(
        \ANSWER/mem[4][4][4] ) );
  dp_1 \ANSWER/mem_reg[4][5][4]  ( .ip(n3457), .ck(clk), .q(
        \ANSWER/mem[4][5][4] ) );
  dp_1 \ANSWER/mem_reg[4][6][4]  ( .ip(n3456), .ck(clk), .q(
        \ANSWER/mem[4][6][4] ) );
  dp_1 \ANSWER/mem_reg[4][7][4]  ( .ip(n3455), .ck(clk), .q(
        \ANSWER/mem[4][7][4] ) );
  dp_1 \ANSWER/mem_reg[4][8][4]  ( .ip(n3454), .ck(clk), .q(
        \ANSWER/mem[4][8][4] ) );
  dp_1 \ANSWER/mem_reg[4][9][4]  ( .ip(n3453), .ck(clk), .q(
        \ANSWER/mem[4][9][4] ) );
  dp_1 \ANSWER/mem_reg[5][0][4]  ( .ip(n3452), .ck(clk), .q(
        \ANSWER/mem[5][0][4] ) );
  dp_1 \ANSWER/mem_reg[5][1][4]  ( .ip(n3451), .ck(clk), .q(
        \ANSWER/mem[5][1][4] ) );
  dp_1 \ANSWER/mem_reg[5][2][4]  ( .ip(n3450), .ck(clk), .q(
        \ANSWER/mem[5][2][4] ) );
  dp_1 \ANSWER/mem_reg[5][3][4]  ( .ip(n3449), .ck(clk), .q(
        \ANSWER/mem[5][3][4] ) );
  dp_1 \ANSWER/mem_reg[5][4][4]  ( .ip(n3448), .ck(clk), .q(
        \ANSWER/mem[5][4][4] ) );
  dp_1 \ANSWER/mem_reg[5][5][4]  ( .ip(n3447), .ck(clk), .q(
        \ANSWER/mem[5][5][4] ) );
  dp_1 \ANSWER/mem_reg[5][6][4]  ( .ip(n3446), .ck(clk), .q(
        \ANSWER/mem[5][6][4] ) );
  dp_1 \ANSWER/mem_reg[5][7][4]  ( .ip(n3445), .ck(clk), .q(
        \ANSWER/mem[5][7][4] ) );
  dp_1 \ANSWER/mem_reg[5][8][4]  ( .ip(n3444), .ck(clk), .q(
        \ANSWER/mem[5][8][4] ) );
  dp_1 \ANSWER/mem_reg[5][9][4]  ( .ip(n3443), .ck(clk), .q(
        \ANSWER/mem[5][9][4] ) );
  dp_1 \ANSWER/mem_reg[6][0][4]  ( .ip(n3442), .ck(clk), .q(
        \ANSWER/mem[6][0][4] ) );
  dp_1 \ANSWER/mem_reg[6][1][4]  ( .ip(n3441), .ck(clk), .q(
        \ANSWER/mem[6][1][4] ) );
  dp_1 \ANSWER/mem_reg[6][2][4]  ( .ip(n3440), .ck(clk), .q(
        \ANSWER/mem[6][2][4] ) );
  dp_1 \ANSWER/mem_reg[6][3][4]  ( .ip(n3439), .ck(clk), .q(
        \ANSWER/mem[6][3][4] ) );
  dp_1 \ANSWER/mem_reg[6][4][4]  ( .ip(n3438), .ck(clk), .q(
        \ANSWER/mem[6][4][4] ) );
  dp_1 \ANSWER/mem_reg[6][5][4]  ( .ip(n3437), .ck(clk), .q(
        \ANSWER/mem[6][5][4] ) );
  dp_1 \ANSWER/mem_reg[6][6][4]  ( .ip(n3436), .ck(clk), .q(
        \ANSWER/mem[6][6][4] ) );
  dp_1 \ANSWER/mem_reg[6][7][4]  ( .ip(n3435), .ck(clk), .q(
        \ANSWER/mem[6][7][4] ) );
  dp_1 \ANSWER/mem_reg[6][8][4]  ( .ip(n3434), .ck(clk), .q(
        \ANSWER/mem[6][8][4] ) );
  dp_1 \ANSWER/mem_reg[6][9][4]  ( .ip(n3433), .ck(clk), .q(
        \ANSWER/mem[6][9][4] ) );
  dp_1 \ANSWER/mem_reg[7][0][4]  ( .ip(n3432), .ck(clk), .q(
        \ANSWER/mem[7][0][4] ) );
  dp_1 \ANSWER/mem_reg[7][1][4]  ( .ip(n3431), .ck(clk), .q(
        \ANSWER/mem[7][1][4] ) );
  dp_1 \ANSWER/mem_reg[7][2][4]  ( .ip(n3430), .ck(clk), .q(
        \ANSWER/mem[7][2][4] ) );
  dp_1 \ANSWER/mem_reg[7][3][4]  ( .ip(n3429), .ck(clk), .q(
        \ANSWER/mem[7][3][4] ) );
  dp_1 \ANSWER/mem_reg[7][4][4]  ( .ip(n3428), .ck(clk), .q(
        \ANSWER/mem[7][4][4] ) );
  dp_1 \ANSWER/mem_reg[7][5][4]  ( .ip(n3427), .ck(clk), .q(
        \ANSWER/mem[7][5][4] ) );
  dp_1 \ANSWER/mem_reg[7][6][4]  ( .ip(n3426), .ck(clk), .q(
        \ANSWER/mem[7][6][4] ) );
  dp_1 \ANSWER/mem_reg[7][7][4]  ( .ip(n3425), .ck(clk), .q(
        \ANSWER/mem[7][7][4] ) );
  dp_1 \ANSWER/mem_reg[7][8][4]  ( .ip(n3424), .ck(clk), .q(
        \ANSWER/mem[7][8][4] ) );
  dp_1 \ANSWER/mem_reg[7][9][4]  ( .ip(n3423), .ck(clk), .q(
        \ANSWER/mem[7][9][4] ) );
  dp_1 \ANSWER/mem_reg[8][0][4]  ( .ip(n3422), .ck(clk), .q(
        \ANSWER/mem[8][0][4] ) );
  dp_1 \ANSWER/mem_reg[8][1][4]  ( .ip(n3421), .ck(clk), .q(
        \ANSWER/mem[8][1][4] ) );
  dp_1 \ANSWER/mem_reg[8][2][4]  ( .ip(n3420), .ck(clk), .q(
        \ANSWER/mem[8][2][4] ) );
  dp_1 \ANSWER/mem_reg[8][3][4]  ( .ip(n3419), .ck(clk), .q(
        \ANSWER/mem[8][3][4] ) );
  dp_1 \ANSWER/mem_reg[8][4][4]  ( .ip(n3418), .ck(clk), .q(
        \ANSWER/mem[8][4][4] ) );
  dp_1 \ANSWER/mem_reg[8][5][4]  ( .ip(n3417), .ck(clk), .q(
        \ANSWER/mem[8][5][4] ) );
  dp_1 \ANSWER/mem_reg[8][6][4]  ( .ip(n3416), .ck(clk), .q(
        \ANSWER/mem[8][6][4] ) );
  dp_1 \ANSWER/mem_reg[8][7][4]  ( .ip(n3415), .ck(clk), .q(
        \ANSWER/mem[8][7][4] ) );
  dp_1 \ANSWER/mem_reg[8][8][4]  ( .ip(n3414), .ck(clk), .q(
        \ANSWER/mem[8][8][4] ) );
  dp_1 \ANSWER/mem_reg[8][9][4]  ( .ip(n3413), .ck(clk), .q(
        \ANSWER/mem[8][9][4] ) );
  dp_1 \ANSWER/mem_reg[9][0][4]  ( .ip(n3412), .ck(clk), .q(
        \ANSWER/mem[9][0][4] ) );
  dp_1 \ANSWER/mem_reg[9][1][4]  ( .ip(n3411), .ck(clk), .q(
        \ANSWER/mem[9][1][4] ) );
  dp_1 \ANSWER/mem_reg[9][2][4]  ( .ip(n3410), .ck(clk), .q(
        \ANSWER/mem[9][2][4] ) );
  dp_1 \ANSWER/mem_reg[9][3][4]  ( .ip(n3409), .ck(clk), .q(
        \ANSWER/mem[9][3][4] ) );
  dp_1 \ANSWER/mem_reg[9][4][4]  ( .ip(n3408), .ck(clk), .q(
        \ANSWER/mem[9][4][4] ) );
  dp_1 \ANSWER/mem_reg[9][5][4]  ( .ip(n3407), .ck(clk), .q(
        \ANSWER/mem[9][5][4] ) );
  dp_1 \ANSWER/mem_reg[9][6][4]  ( .ip(n3406), .ck(clk), .q(
        \ANSWER/mem[9][6][4] ) );
  dp_1 \ANSWER/mem_reg[9][7][4]  ( .ip(n3405), .ck(clk), .q(
        \ANSWER/mem[9][7][4] ) );
  dp_1 \ANSWER/mem_reg[9][8][4]  ( .ip(n3404), .ck(clk), .q(
        \ANSWER/mem[9][8][4] ) );
  dp_1 \ANSWER/mem_reg[9][9][4]  ( .ip(n3403), .ck(clk), .q(
        \ANSWER/mem[9][9][4] ) );
  dp_1 \SIGMOID/lut_out_reg[5]  ( .ip(n3905), .ck(clk), .q(
        \SIGMOID/lut_out [5]) );
  dp_1 \ANSWER/mem_reg[0][0][5]  ( .ip(n3402), .ck(clk), .q(
        \ANSWER/mem[0][0][5] ) );
  dp_1 \ANSWER/mem_reg[0][1][5]  ( .ip(n3401), .ck(clk), .q(
        \ANSWER/mem[0][1][5] ) );
  dp_1 \ANSWER/mem_reg[0][2][5]  ( .ip(n3400), .ck(clk), .q(
        \ANSWER/mem[0][2][5] ) );
  dp_1 \ANSWER/mem_reg[0][3][5]  ( .ip(n3399), .ck(clk), .q(
        \ANSWER/mem[0][3][5] ) );
  dp_1 \ANSWER/mem_reg[0][4][5]  ( .ip(n3398), .ck(clk), .q(
        \ANSWER/mem[0][4][5] ) );
  dp_1 \ANSWER/mem_reg[0][5][5]  ( .ip(n3397), .ck(clk), .q(
        \ANSWER/mem[0][5][5] ) );
  dp_1 \ANSWER/mem_reg[0][6][5]  ( .ip(n3396), .ck(clk), .q(
        \ANSWER/mem[0][6][5] ) );
  dp_1 \ANSWER/mem_reg[0][7][5]  ( .ip(n3395), .ck(clk), .q(
        \ANSWER/mem[0][7][5] ) );
  dp_1 \ANSWER/mem_reg[0][8][5]  ( .ip(n3394), .ck(clk), .q(
        \ANSWER/mem[0][8][5] ) );
  dp_1 \ANSWER/mem_reg[0][9][5]  ( .ip(n3393), .ck(clk), .q(
        \ANSWER/mem[0][9][5] ) );
  dp_1 \ANSWER/mem_reg[1][0][5]  ( .ip(n3392), .ck(clk), .q(
        \ANSWER/mem[1][0][5] ) );
  dp_1 \ANSWER/mem_reg[1][1][5]  ( .ip(n3391), .ck(clk), .q(
        \ANSWER/mem[1][1][5] ) );
  dp_1 \ANSWER/mem_reg[1][2][5]  ( .ip(n3390), .ck(clk), .q(
        \ANSWER/mem[1][2][5] ) );
  dp_1 \ANSWER/mem_reg[1][3][5]  ( .ip(n3389), .ck(clk), .q(
        \ANSWER/mem[1][3][5] ) );
  dp_1 \ANSWER/mem_reg[1][4][5]  ( .ip(n3388), .ck(clk), .q(
        \ANSWER/mem[1][4][5] ) );
  dp_1 \ANSWER/mem_reg[1][5][5]  ( .ip(n3387), .ck(clk), .q(
        \ANSWER/mem[1][5][5] ) );
  dp_1 \ANSWER/mem_reg[1][6][5]  ( .ip(n3386), .ck(clk), .q(
        \ANSWER/mem[1][6][5] ) );
  dp_1 \ANSWER/mem_reg[1][7][5]  ( .ip(n3385), .ck(clk), .q(
        \ANSWER/mem[1][7][5] ) );
  dp_1 \ANSWER/mem_reg[1][8][5]  ( .ip(n3384), .ck(clk), .q(
        \ANSWER/mem[1][8][5] ) );
  dp_1 \ANSWER/mem_reg[1][9][5]  ( .ip(n3383), .ck(clk), .q(
        \ANSWER/mem[1][9][5] ) );
  dp_1 \ANSWER/mem_reg[2][0][5]  ( .ip(n3382), .ck(clk), .q(
        \ANSWER/mem[2][0][5] ) );
  dp_1 \ANSWER/mem_reg[2][1][5]  ( .ip(n3381), .ck(clk), .q(
        \ANSWER/mem[2][1][5] ) );
  dp_1 \ANSWER/mem_reg[2][2][5]  ( .ip(n3380), .ck(clk), .q(
        \ANSWER/mem[2][2][5] ) );
  dp_1 \ANSWER/mem_reg[2][3][5]  ( .ip(n3379), .ck(clk), .q(
        \ANSWER/mem[2][3][5] ) );
  dp_1 \ANSWER/mem_reg[2][4][5]  ( .ip(n3378), .ck(clk), .q(
        \ANSWER/mem[2][4][5] ) );
  dp_1 \ANSWER/mem_reg[2][5][5]  ( .ip(n3377), .ck(clk), .q(
        \ANSWER/mem[2][5][5] ) );
  dp_1 \ANSWER/mem_reg[2][6][5]  ( .ip(n3376), .ck(clk), .q(
        \ANSWER/mem[2][6][5] ) );
  dp_1 \ANSWER/mem_reg[2][7][5]  ( .ip(n3375), .ck(clk), .q(
        \ANSWER/mem[2][7][5] ) );
  dp_1 \ANSWER/mem_reg[2][8][5]  ( .ip(n3374), .ck(clk), .q(
        \ANSWER/mem[2][8][5] ) );
  dp_1 \ANSWER/mem_reg[2][9][5]  ( .ip(n3373), .ck(clk), .q(
        \ANSWER/mem[2][9][5] ) );
  dp_1 \ANSWER/mem_reg[3][0][5]  ( .ip(n3372), .ck(clk), .q(
        \ANSWER/mem[3][0][5] ) );
  dp_1 \ANSWER/mem_reg[3][1][5]  ( .ip(n3371), .ck(clk), .q(
        \ANSWER/mem[3][1][5] ) );
  dp_1 \ANSWER/mem_reg[3][2][5]  ( .ip(n3370), .ck(clk), .q(
        \ANSWER/mem[3][2][5] ) );
  dp_1 \ANSWER/mem_reg[3][3][5]  ( .ip(n3369), .ck(clk), .q(
        \ANSWER/mem[3][3][5] ) );
  dp_1 \ANSWER/mem_reg[3][4][5]  ( .ip(n3368), .ck(clk), .q(
        \ANSWER/mem[3][4][5] ) );
  dp_1 \ANSWER/mem_reg[3][5][5]  ( .ip(n3367), .ck(clk), .q(
        \ANSWER/mem[3][5][5] ) );
  dp_1 \ANSWER/mem_reg[3][6][5]  ( .ip(n3366), .ck(clk), .q(
        \ANSWER/mem[3][6][5] ) );
  dp_1 \ANSWER/mem_reg[3][7][5]  ( .ip(n3365), .ck(clk), .q(
        \ANSWER/mem[3][7][5] ) );
  dp_1 \ANSWER/mem_reg[3][8][5]  ( .ip(n3364), .ck(clk), .q(
        \ANSWER/mem[3][8][5] ) );
  dp_1 \ANSWER/mem_reg[3][9][5]  ( .ip(n3363), .ck(clk), .q(
        \ANSWER/mem[3][9][5] ) );
  dp_1 \ANSWER/mem_reg[4][0][5]  ( .ip(n3362), .ck(clk), .q(
        \ANSWER/mem[4][0][5] ) );
  dp_1 \ANSWER/mem_reg[4][1][5]  ( .ip(n3361), .ck(clk), .q(
        \ANSWER/mem[4][1][5] ) );
  dp_1 \ANSWER/mem_reg[4][2][5]  ( .ip(n3360), .ck(clk), .q(
        \ANSWER/mem[4][2][5] ) );
  dp_1 \ANSWER/mem_reg[4][3][5]  ( .ip(n3359), .ck(clk), .q(
        \ANSWER/mem[4][3][5] ) );
  dp_1 \ANSWER/mem_reg[4][4][5]  ( .ip(n3358), .ck(clk), .q(
        \ANSWER/mem[4][4][5] ) );
  dp_1 \ANSWER/mem_reg[4][5][5]  ( .ip(n3357), .ck(clk), .q(
        \ANSWER/mem[4][5][5] ) );
  dp_1 \ANSWER/mem_reg[4][6][5]  ( .ip(n3356), .ck(clk), .q(
        \ANSWER/mem[4][6][5] ) );
  dp_1 \ANSWER/mem_reg[4][7][5]  ( .ip(n3355), .ck(clk), .q(
        \ANSWER/mem[4][7][5] ) );
  dp_1 \ANSWER/mem_reg[4][8][5]  ( .ip(n3354), .ck(clk), .q(
        \ANSWER/mem[4][8][5] ) );
  dp_1 \ANSWER/mem_reg[4][9][5]  ( .ip(n3353), .ck(clk), .q(
        \ANSWER/mem[4][9][5] ) );
  dp_1 \ANSWER/mem_reg[5][0][5]  ( .ip(n3352), .ck(clk), .q(
        \ANSWER/mem[5][0][5] ) );
  dp_1 \ANSWER/mem_reg[5][1][5]  ( .ip(n3351), .ck(clk), .q(
        \ANSWER/mem[5][1][5] ) );
  dp_1 \ANSWER/mem_reg[5][2][5]  ( .ip(n3350), .ck(clk), .q(
        \ANSWER/mem[5][2][5] ) );
  dp_1 \ANSWER/mem_reg[5][3][5]  ( .ip(n3349), .ck(clk), .q(
        \ANSWER/mem[5][3][5] ) );
  dp_1 \ANSWER/mem_reg[5][4][5]  ( .ip(n3348), .ck(clk), .q(
        \ANSWER/mem[5][4][5] ) );
  dp_1 \ANSWER/mem_reg[5][5][5]  ( .ip(n3347), .ck(clk), .q(
        \ANSWER/mem[5][5][5] ) );
  dp_1 \ANSWER/mem_reg[5][6][5]  ( .ip(n3346), .ck(clk), .q(
        \ANSWER/mem[5][6][5] ) );
  dp_1 \ANSWER/mem_reg[5][7][5]  ( .ip(n3345), .ck(clk), .q(
        \ANSWER/mem[5][7][5] ) );
  dp_1 \ANSWER/mem_reg[5][8][5]  ( .ip(n3344), .ck(clk), .q(
        \ANSWER/mem[5][8][5] ) );
  dp_1 \ANSWER/mem_reg[5][9][5]  ( .ip(n3343), .ck(clk), .q(
        \ANSWER/mem[5][9][5] ) );
  dp_1 \ANSWER/mem_reg[6][0][5]  ( .ip(n3342), .ck(clk), .q(
        \ANSWER/mem[6][0][5] ) );
  dp_1 \ANSWER/mem_reg[6][1][5]  ( .ip(n3341), .ck(clk), .q(
        \ANSWER/mem[6][1][5] ) );
  dp_1 \ANSWER/mem_reg[6][2][5]  ( .ip(n3340), .ck(clk), .q(
        \ANSWER/mem[6][2][5] ) );
  dp_1 \ANSWER/mem_reg[6][3][5]  ( .ip(n3339), .ck(clk), .q(
        \ANSWER/mem[6][3][5] ) );
  dp_1 \ANSWER/mem_reg[6][4][5]  ( .ip(n3338), .ck(clk), .q(
        \ANSWER/mem[6][4][5] ) );
  dp_1 \ANSWER/mem_reg[6][5][5]  ( .ip(n3337), .ck(clk), .q(
        \ANSWER/mem[6][5][5] ) );
  dp_1 \ANSWER/mem_reg[6][6][5]  ( .ip(n3336), .ck(clk), .q(
        \ANSWER/mem[6][6][5] ) );
  dp_1 \ANSWER/mem_reg[6][7][5]  ( .ip(n3335), .ck(clk), .q(
        \ANSWER/mem[6][7][5] ) );
  dp_1 \ANSWER/mem_reg[6][8][5]  ( .ip(n3334), .ck(clk), .q(
        \ANSWER/mem[6][8][5] ) );
  dp_1 \ANSWER/mem_reg[6][9][5]  ( .ip(n3333), .ck(clk), .q(
        \ANSWER/mem[6][9][5] ) );
  dp_1 \ANSWER/mem_reg[7][0][5]  ( .ip(n3332), .ck(clk), .q(
        \ANSWER/mem[7][0][5] ) );
  dp_1 \ANSWER/mem_reg[7][1][5]  ( .ip(n3331), .ck(clk), .q(
        \ANSWER/mem[7][1][5] ) );
  dp_1 \ANSWER/mem_reg[7][2][5]  ( .ip(n3330), .ck(clk), .q(
        \ANSWER/mem[7][2][5] ) );
  dp_1 \ANSWER/mem_reg[7][3][5]  ( .ip(n3329), .ck(clk), .q(
        \ANSWER/mem[7][3][5] ) );
  dp_1 \ANSWER/mem_reg[7][4][5]  ( .ip(n3328), .ck(clk), .q(
        \ANSWER/mem[7][4][5] ) );
  dp_1 \ANSWER/mem_reg[7][5][5]  ( .ip(n3327), .ck(clk), .q(
        \ANSWER/mem[7][5][5] ) );
  dp_1 \ANSWER/mem_reg[7][6][5]  ( .ip(n3326), .ck(clk), .q(
        \ANSWER/mem[7][6][5] ) );
  dp_1 \ANSWER/mem_reg[7][7][5]  ( .ip(n3325), .ck(clk), .q(
        \ANSWER/mem[7][7][5] ) );
  dp_1 \ANSWER/mem_reg[7][8][5]  ( .ip(n3324), .ck(clk), .q(
        \ANSWER/mem[7][8][5] ) );
  dp_1 \ANSWER/mem_reg[7][9][5]  ( .ip(n3323), .ck(clk), .q(
        \ANSWER/mem[7][9][5] ) );
  dp_1 \ANSWER/mem_reg[8][0][5]  ( .ip(n3322), .ck(clk), .q(
        \ANSWER/mem[8][0][5] ) );
  dp_1 \ANSWER/mem_reg[8][1][5]  ( .ip(n3321), .ck(clk), .q(
        \ANSWER/mem[8][1][5] ) );
  dp_1 \ANSWER/mem_reg[8][2][5]  ( .ip(n3320), .ck(clk), .q(
        \ANSWER/mem[8][2][5] ) );
  dp_1 \ANSWER/mem_reg[8][3][5]  ( .ip(n3319), .ck(clk), .q(
        \ANSWER/mem[8][3][5] ) );
  dp_1 \ANSWER/mem_reg[8][4][5]  ( .ip(n3318), .ck(clk), .q(
        \ANSWER/mem[8][4][5] ) );
  dp_1 \ANSWER/mem_reg[8][5][5]  ( .ip(n3317), .ck(clk), .q(
        \ANSWER/mem[8][5][5] ) );
  dp_1 \ANSWER/mem_reg[8][6][5]  ( .ip(n3316), .ck(clk), .q(
        \ANSWER/mem[8][6][5] ) );
  dp_1 \ANSWER/mem_reg[8][7][5]  ( .ip(n3315), .ck(clk), .q(
        \ANSWER/mem[8][7][5] ) );
  dp_1 \ANSWER/mem_reg[8][8][5]  ( .ip(n3314), .ck(clk), .q(
        \ANSWER/mem[8][8][5] ) );
  dp_1 \ANSWER/mem_reg[8][9][5]  ( .ip(n3313), .ck(clk), .q(
        \ANSWER/mem[8][9][5] ) );
  dp_1 \ANSWER/mem_reg[9][0][5]  ( .ip(n3312), .ck(clk), .q(
        \ANSWER/mem[9][0][5] ) );
  dp_1 \ANSWER/mem_reg[9][1][5]  ( .ip(n3311), .ck(clk), .q(
        \ANSWER/mem[9][1][5] ) );
  dp_1 \ANSWER/mem_reg[9][2][5]  ( .ip(n3310), .ck(clk), .q(
        \ANSWER/mem[9][2][5] ) );
  dp_1 \ANSWER/mem_reg[9][3][5]  ( .ip(n3309), .ck(clk), .q(
        \ANSWER/mem[9][3][5] ) );
  dp_1 \ANSWER/mem_reg[9][4][5]  ( .ip(n3308), .ck(clk), .q(
        \ANSWER/mem[9][4][5] ) );
  dp_1 \ANSWER/mem_reg[9][5][5]  ( .ip(n3307), .ck(clk), .q(
        \ANSWER/mem[9][5][5] ) );
  dp_1 \ANSWER/mem_reg[9][6][5]  ( .ip(n3306), .ck(clk), .q(
        \ANSWER/mem[9][6][5] ) );
  dp_1 \ANSWER/mem_reg[9][7][5]  ( .ip(n3305), .ck(clk), .q(
        \ANSWER/mem[9][7][5] ) );
  dp_1 \ANSWER/mem_reg[9][8][5]  ( .ip(n3304), .ck(clk), .q(
        \ANSWER/mem[9][8][5] ) );
  dp_1 \ANSWER/mem_reg[9][9][5]  ( .ip(n3303), .ck(clk), .q(
        \ANSWER/mem[9][9][5] ) );
  dp_1 \SIGMOID/lut_out_reg[6]  ( .ip(n3904), .ck(clk), .q(
        \SIGMOID/lut_out [6]) );
  dp_1 \ANSWER/mem_reg[0][0][6]  ( .ip(n3302), .ck(clk), .q(
        \ANSWER/mem[0][0][6] ) );
  dp_1 \ANSWER/mem_reg[0][1][6]  ( .ip(n3301), .ck(clk), .q(
        \ANSWER/mem[0][1][6] ) );
  dp_1 \ANSWER/mem_reg[0][2][6]  ( .ip(n3300), .ck(clk), .q(
        \ANSWER/mem[0][2][6] ) );
  dp_1 \ANSWER/mem_reg[0][3][6]  ( .ip(n3299), .ck(clk), .q(
        \ANSWER/mem[0][3][6] ) );
  dp_1 \ANSWER/mem_reg[0][4][6]  ( .ip(n3298), .ck(clk), .q(
        \ANSWER/mem[0][4][6] ) );
  dp_1 \ANSWER/mem_reg[0][5][6]  ( .ip(n3297), .ck(clk), .q(
        \ANSWER/mem[0][5][6] ) );
  dp_1 \ANSWER/mem_reg[0][6][6]  ( .ip(n3296), .ck(clk), .q(
        \ANSWER/mem[0][6][6] ) );
  dp_1 \ANSWER/mem_reg[0][7][6]  ( .ip(n3295), .ck(clk), .q(
        \ANSWER/mem[0][7][6] ) );
  dp_1 \ANSWER/mem_reg[0][8][6]  ( .ip(n3294), .ck(clk), .q(
        \ANSWER/mem[0][8][6] ) );
  dp_1 \ANSWER/mem_reg[0][9][6]  ( .ip(n3293), .ck(clk), .q(
        \ANSWER/mem[0][9][6] ) );
  dp_1 \ANSWER/mem_reg[1][0][6]  ( .ip(n3292), .ck(clk), .q(
        \ANSWER/mem[1][0][6] ) );
  dp_1 \ANSWER/mem_reg[1][1][6]  ( .ip(n3291), .ck(clk), .q(
        \ANSWER/mem[1][1][6] ) );
  dp_1 \ANSWER/mem_reg[1][2][6]  ( .ip(n3290), .ck(clk), .q(
        \ANSWER/mem[1][2][6] ) );
  dp_1 \ANSWER/mem_reg[1][3][6]  ( .ip(n3289), .ck(clk), .q(
        \ANSWER/mem[1][3][6] ) );
  dp_1 \ANSWER/mem_reg[1][4][6]  ( .ip(n3288), .ck(clk), .q(
        \ANSWER/mem[1][4][6] ) );
  dp_1 \ANSWER/mem_reg[1][5][6]  ( .ip(n3287), .ck(clk), .q(
        \ANSWER/mem[1][5][6] ) );
  dp_1 \ANSWER/mem_reg[1][6][6]  ( .ip(n3286), .ck(clk), .q(
        \ANSWER/mem[1][6][6] ) );
  dp_1 \ANSWER/mem_reg[1][7][6]  ( .ip(n3285), .ck(clk), .q(
        \ANSWER/mem[1][7][6] ) );
  dp_1 \ANSWER/mem_reg[1][8][6]  ( .ip(n3284), .ck(clk), .q(
        \ANSWER/mem[1][8][6] ) );
  dp_1 \ANSWER/mem_reg[1][9][6]  ( .ip(n3283), .ck(clk), .q(
        \ANSWER/mem[1][9][6] ) );
  dp_1 \ANSWER/mem_reg[2][0][6]  ( .ip(n3282), .ck(clk), .q(
        \ANSWER/mem[2][0][6] ) );
  dp_1 \ANSWER/mem_reg[2][1][6]  ( .ip(n3281), .ck(clk), .q(
        \ANSWER/mem[2][1][6] ) );
  dp_1 \ANSWER/mem_reg[2][2][6]  ( .ip(n3280), .ck(clk), .q(
        \ANSWER/mem[2][2][6] ) );
  dp_1 \ANSWER/mem_reg[2][3][6]  ( .ip(n3279), .ck(clk), .q(
        \ANSWER/mem[2][3][6] ) );
  dp_1 \ANSWER/mem_reg[2][4][6]  ( .ip(n3278), .ck(clk), .q(
        \ANSWER/mem[2][4][6] ) );
  dp_1 \ANSWER/mem_reg[2][5][6]  ( .ip(n3277), .ck(clk), .q(
        \ANSWER/mem[2][5][6] ) );
  dp_1 \ANSWER/mem_reg[2][6][6]  ( .ip(n3276), .ck(clk), .q(
        \ANSWER/mem[2][6][6] ) );
  dp_1 \ANSWER/mem_reg[2][7][6]  ( .ip(n3275), .ck(clk), .q(
        \ANSWER/mem[2][7][6] ) );
  dp_1 \ANSWER/mem_reg[2][8][6]  ( .ip(n3274), .ck(clk), .q(
        \ANSWER/mem[2][8][6] ) );
  dp_1 \ANSWER/mem_reg[2][9][6]  ( .ip(n3273), .ck(clk), .q(
        \ANSWER/mem[2][9][6] ) );
  dp_1 \ANSWER/mem_reg[3][0][6]  ( .ip(n3272), .ck(clk), .q(
        \ANSWER/mem[3][0][6] ) );
  dp_1 \ANSWER/mem_reg[3][1][6]  ( .ip(n3271), .ck(clk), .q(
        \ANSWER/mem[3][1][6] ) );
  dp_1 \ANSWER/mem_reg[3][2][6]  ( .ip(n3270), .ck(clk), .q(
        \ANSWER/mem[3][2][6] ) );
  dp_1 \ANSWER/mem_reg[3][3][6]  ( .ip(n3269), .ck(clk), .q(
        \ANSWER/mem[3][3][6] ) );
  dp_1 \ANSWER/mem_reg[3][4][6]  ( .ip(n3268), .ck(clk), .q(
        \ANSWER/mem[3][4][6] ) );
  dp_1 \ANSWER/mem_reg[3][5][6]  ( .ip(n3267), .ck(clk), .q(
        \ANSWER/mem[3][5][6] ) );
  dp_1 \ANSWER/mem_reg[3][6][6]  ( .ip(n3266), .ck(clk), .q(
        \ANSWER/mem[3][6][6] ) );
  dp_1 \ANSWER/mem_reg[3][7][6]  ( .ip(n3265), .ck(clk), .q(
        \ANSWER/mem[3][7][6] ) );
  dp_1 \ANSWER/mem_reg[3][8][6]  ( .ip(n3264), .ck(clk), .q(
        \ANSWER/mem[3][8][6] ) );
  dp_1 \ANSWER/mem_reg[3][9][6]  ( .ip(n3263), .ck(clk), .q(
        \ANSWER/mem[3][9][6] ) );
  dp_1 \ANSWER/mem_reg[4][0][6]  ( .ip(n3262), .ck(clk), .q(
        \ANSWER/mem[4][0][6] ) );
  dp_1 \ANSWER/mem_reg[4][1][6]  ( .ip(n3261), .ck(clk), .q(
        \ANSWER/mem[4][1][6] ) );
  dp_1 \ANSWER/mem_reg[4][2][6]  ( .ip(n3260), .ck(clk), .q(
        \ANSWER/mem[4][2][6] ) );
  dp_1 \ANSWER/mem_reg[4][3][6]  ( .ip(n3259), .ck(clk), .q(
        \ANSWER/mem[4][3][6] ) );
  dp_1 \ANSWER/mem_reg[4][4][6]  ( .ip(n3258), .ck(clk), .q(
        \ANSWER/mem[4][4][6] ) );
  dp_1 \ANSWER/mem_reg[4][5][6]  ( .ip(n3257), .ck(clk), .q(
        \ANSWER/mem[4][5][6] ) );
  dp_1 \ANSWER/mem_reg[4][6][6]  ( .ip(n3256), .ck(clk), .q(
        \ANSWER/mem[4][6][6] ) );
  dp_1 \ANSWER/mem_reg[4][7][6]  ( .ip(n3255), .ck(clk), .q(
        \ANSWER/mem[4][7][6] ) );
  dp_1 \ANSWER/mem_reg[4][8][6]  ( .ip(n3254), .ck(clk), .q(
        \ANSWER/mem[4][8][6] ) );
  dp_1 \ANSWER/mem_reg[4][9][6]  ( .ip(n3253), .ck(clk), .q(
        \ANSWER/mem[4][9][6] ) );
  dp_1 \ANSWER/mem_reg[5][0][6]  ( .ip(n3252), .ck(clk), .q(
        \ANSWER/mem[5][0][6] ) );
  dp_1 \ANSWER/mem_reg[5][1][6]  ( .ip(n3251), .ck(clk), .q(
        \ANSWER/mem[5][1][6] ) );
  dp_1 \ANSWER/mem_reg[5][2][6]  ( .ip(n3250), .ck(clk), .q(
        \ANSWER/mem[5][2][6] ) );
  dp_1 \ANSWER/mem_reg[5][3][6]  ( .ip(n3249), .ck(clk), .q(
        \ANSWER/mem[5][3][6] ) );
  dp_1 \ANSWER/mem_reg[5][4][6]  ( .ip(n3248), .ck(clk), .q(
        \ANSWER/mem[5][4][6] ) );
  dp_1 \ANSWER/mem_reg[5][5][6]  ( .ip(n3247), .ck(clk), .q(
        \ANSWER/mem[5][5][6] ) );
  dp_1 \ANSWER/mem_reg[5][6][6]  ( .ip(n3246), .ck(clk), .q(
        \ANSWER/mem[5][6][6] ) );
  dp_1 \ANSWER/mem_reg[5][7][6]  ( .ip(n3245), .ck(clk), .q(
        \ANSWER/mem[5][7][6] ) );
  dp_1 \ANSWER/mem_reg[5][8][6]  ( .ip(n3244), .ck(clk), .q(
        \ANSWER/mem[5][8][6] ) );
  dp_1 \ANSWER/mem_reg[5][9][6]  ( .ip(n3243), .ck(clk), .q(
        \ANSWER/mem[5][9][6] ) );
  dp_1 \ANSWER/mem_reg[6][0][6]  ( .ip(n3242), .ck(clk), .q(
        \ANSWER/mem[6][0][6] ) );
  dp_1 \ANSWER/mem_reg[6][1][6]  ( .ip(n3241), .ck(clk), .q(
        \ANSWER/mem[6][1][6] ) );
  dp_1 \ANSWER/mem_reg[6][2][6]  ( .ip(n3240), .ck(clk), .q(
        \ANSWER/mem[6][2][6] ) );
  dp_1 \ANSWER/mem_reg[6][3][6]  ( .ip(n3239), .ck(clk), .q(
        \ANSWER/mem[6][3][6] ) );
  dp_1 \ANSWER/mem_reg[6][4][6]  ( .ip(n3238), .ck(clk), .q(
        \ANSWER/mem[6][4][6] ) );
  dp_1 \ANSWER/mem_reg[6][5][6]  ( .ip(n3237), .ck(clk), .q(
        \ANSWER/mem[6][5][6] ) );
  dp_1 \ANSWER/mem_reg[6][6][6]  ( .ip(n3236), .ck(clk), .q(
        \ANSWER/mem[6][6][6] ) );
  dp_1 \ANSWER/mem_reg[6][7][6]  ( .ip(n3235), .ck(clk), .q(
        \ANSWER/mem[6][7][6] ) );
  dp_1 \ANSWER/mem_reg[6][8][6]  ( .ip(n3234), .ck(clk), .q(
        \ANSWER/mem[6][8][6] ) );
  dp_1 \ANSWER/mem_reg[6][9][6]  ( .ip(n3233), .ck(clk), .q(
        \ANSWER/mem[6][9][6] ) );
  dp_1 \ANSWER/mem_reg[7][0][6]  ( .ip(n3232), .ck(clk), .q(
        \ANSWER/mem[7][0][6] ) );
  dp_1 \ANSWER/mem_reg[7][1][6]  ( .ip(n3231), .ck(clk), .q(
        \ANSWER/mem[7][1][6] ) );
  dp_1 \ANSWER/mem_reg[7][2][6]  ( .ip(n3230), .ck(clk), .q(
        \ANSWER/mem[7][2][6] ) );
  dp_1 \ANSWER/mem_reg[7][3][6]  ( .ip(n3229), .ck(clk), .q(
        \ANSWER/mem[7][3][6] ) );
  dp_1 \ANSWER/mem_reg[7][4][6]  ( .ip(n3228), .ck(clk), .q(
        \ANSWER/mem[7][4][6] ) );
  dp_1 \ANSWER/mem_reg[7][5][6]  ( .ip(n3227), .ck(clk), .q(
        \ANSWER/mem[7][5][6] ) );
  dp_1 \ANSWER/mem_reg[7][6][6]  ( .ip(n3226), .ck(clk), .q(
        \ANSWER/mem[7][6][6] ) );
  dp_1 \ANSWER/mem_reg[7][7][6]  ( .ip(n3225), .ck(clk), .q(
        \ANSWER/mem[7][7][6] ) );
  dp_1 \ANSWER/mem_reg[7][8][6]  ( .ip(n3224), .ck(clk), .q(
        \ANSWER/mem[7][8][6] ) );
  dp_1 \ANSWER/mem_reg[7][9][6]  ( .ip(n3223), .ck(clk), .q(
        \ANSWER/mem[7][9][6] ) );
  dp_1 \ANSWER/mem_reg[8][0][6]  ( .ip(n3222), .ck(clk), .q(
        \ANSWER/mem[8][0][6] ) );
  dp_1 \ANSWER/mem_reg[8][1][6]  ( .ip(n3221), .ck(clk), .q(
        \ANSWER/mem[8][1][6] ) );
  dp_1 \ANSWER/mem_reg[8][2][6]  ( .ip(n3220), .ck(clk), .q(
        \ANSWER/mem[8][2][6] ) );
  dp_1 \ANSWER/mem_reg[8][3][6]  ( .ip(n3219), .ck(clk), .q(
        \ANSWER/mem[8][3][6] ) );
  dp_1 \ANSWER/mem_reg[8][4][6]  ( .ip(n3218), .ck(clk), .q(
        \ANSWER/mem[8][4][6] ) );
  dp_1 \ANSWER/mem_reg[8][5][6]  ( .ip(n3217), .ck(clk), .q(
        \ANSWER/mem[8][5][6] ) );
  dp_1 \ANSWER/mem_reg[8][6][6]  ( .ip(n3216), .ck(clk), .q(
        \ANSWER/mem[8][6][6] ) );
  dp_1 \ANSWER/mem_reg[8][7][6]  ( .ip(n3215), .ck(clk), .q(
        \ANSWER/mem[8][7][6] ) );
  dp_1 \ANSWER/mem_reg[8][8][6]  ( .ip(n3214), .ck(clk), .q(
        \ANSWER/mem[8][8][6] ) );
  dp_1 \ANSWER/mem_reg[8][9][6]  ( .ip(n3213), .ck(clk), .q(
        \ANSWER/mem[8][9][6] ) );
  dp_1 \ANSWER/mem_reg[9][0][6]  ( .ip(n3212), .ck(clk), .q(
        \ANSWER/mem[9][0][6] ) );
  dp_1 \ANSWER/mem_reg[9][1][6]  ( .ip(n3211), .ck(clk), .q(
        \ANSWER/mem[9][1][6] ) );
  dp_1 \ANSWER/mem_reg[9][2][6]  ( .ip(n3210), .ck(clk), .q(
        \ANSWER/mem[9][2][6] ) );
  dp_1 \ANSWER/mem_reg[9][3][6]  ( .ip(n3209), .ck(clk), .q(
        \ANSWER/mem[9][3][6] ) );
  dp_1 \ANSWER/mem_reg[9][4][6]  ( .ip(n3208), .ck(clk), .q(
        \ANSWER/mem[9][4][6] ) );
  dp_1 \ANSWER/mem_reg[9][5][6]  ( .ip(n3207), .ck(clk), .q(
        \ANSWER/mem[9][5][6] ) );
  dp_1 \ANSWER/mem_reg[9][6][6]  ( .ip(n3206), .ck(clk), .q(
        \ANSWER/mem[9][6][6] ) );
  dp_1 \ANSWER/mem_reg[9][7][6]  ( .ip(n3205), .ck(clk), .q(
        \ANSWER/mem[9][7][6] ) );
  dp_1 \ANSWER/mem_reg[9][8][6]  ( .ip(n3204), .ck(clk), .q(
        \ANSWER/mem[9][8][6] ) );
  dp_1 \ANSWER/mem_reg[9][9][6]  ( .ip(n3203), .ck(clk), .q(
        \ANSWER/mem[9][9][6] ) );
  dp_1 \SIGMOID/lut_out_reg[7]  ( .ip(n3903), .ck(clk), .q(
        \SIGMOID/lut_out [7]) );
  dp_1 \ANSWER/mem_reg[0][0][7]  ( .ip(n3202), .ck(clk), .q(
        \ANSWER/mem[0][0][7] ) );
  dp_1 \ANSWER/mem_reg[0][1][7]  ( .ip(n3201), .ck(clk), .q(
        \ANSWER/mem[0][1][7] ) );
  dp_1 \ANSWER/mem_reg[0][2][7]  ( .ip(n3200), .ck(clk), .q(
        \ANSWER/mem[0][2][7] ) );
  dp_1 \ANSWER/mem_reg[0][3][7]  ( .ip(n3199), .ck(clk), .q(
        \ANSWER/mem[0][3][7] ) );
  dp_1 \ANSWER/mem_reg[0][4][7]  ( .ip(n3198), .ck(clk), .q(
        \ANSWER/mem[0][4][7] ) );
  dp_1 \ANSWER/mem_reg[0][5][7]  ( .ip(n3197), .ck(clk), .q(
        \ANSWER/mem[0][5][7] ) );
  dp_1 \ANSWER/mem_reg[0][6][7]  ( .ip(n3196), .ck(clk), .q(
        \ANSWER/mem[0][6][7] ) );
  dp_1 \ANSWER/mem_reg[0][7][7]  ( .ip(n3195), .ck(clk), .q(
        \ANSWER/mem[0][7][7] ) );
  dp_1 \ANSWER/mem_reg[0][8][7]  ( .ip(n3194), .ck(clk), .q(
        \ANSWER/mem[0][8][7] ) );
  dp_1 \ANSWER/mem_reg[0][9][7]  ( .ip(n3193), .ck(clk), .q(
        \ANSWER/mem[0][9][7] ) );
  dp_1 \ANSWER/mem_reg[1][0][7]  ( .ip(n3192), .ck(clk), .q(
        \ANSWER/mem[1][0][7] ) );
  dp_1 \ANSWER/mem_reg[1][1][7]  ( .ip(n3191), .ck(clk), .q(
        \ANSWER/mem[1][1][7] ) );
  dp_1 \ANSWER/mem_reg[1][2][7]  ( .ip(n3190), .ck(clk), .q(
        \ANSWER/mem[1][2][7] ) );
  dp_1 \ANSWER/mem_reg[1][3][7]  ( .ip(n3189), .ck(clk), .q(
        \ANSWER/mem[1][3][7] ) );
  dp_1 \ANSWER/mem_reg[1][4][7]  ( .ip(n3188), .ck(clk), .q(
        \ANSWER/mem[1][4][7] ) );
  dp_1 \ANSWER/mem_reg[1][5][7]  ( .ip(n3187), .ck(clk), .q(
        \ANSWER/mem[1][5][7] ) );
  dp_1 \ANSWER/mem_reg[1][6][7]  ( .ip(n3186), .ck(clk), .q(
        \ANSWER/mem[1][6][7] ) );
  dp_1 \ANSWER/mem_reg[1][7][7]  ( .ip(n3185), .ck(clk), .q(
        \ANSWER/mem[1][7][7] ) );
  dp_1 \ANSWER/mem_reg[1][8][7]  ( .ip(n3184), .ck(clk), .q(
        \ANSWER/mem[1][8][7] ) );
  dp_1 \ANSWER/mem_reg[1][9][7]  ( .ip(n3183), .ck(clk), .q(
        \ANSWER/mem[1][9][7] ) );
  dp_1 \ANSWER/mem_reg[2][0][7]  ( .ip(n3182), .ck(clk), .q(
        \ANSWER/mem[2][0][7] ) );
  dp_1 \ANSWER/mem_reg[2][1][7]  ( .ip(n3181), .ck(clk), .q(
        \ANSWER/mem[2][1][7] ) );
  dp_1 \ANSWER/mem_reg[2][2][7]  ( .ip(n3180), .ck(clk), .q(
        \ANSWER/mem[2][2][7] ) );
  dp_1 \ANSWER/mem_reg[2][3][7]  ( .ip(n3179), .ck(clk), .q(
        \ANSWER/mem[2][3][7] ) );
  dp_1 \ANSWER/mem_reg[2][4][7]  ( .ip(n3178), .ck(clk), .q(
        \ANSWER/mem[2][4][7] ) );
  dp_1 \ANSWER/mem_reg[2][5][7]  ( .ip(n3177), .ck(clk), .q(
        \ANSWER/mem[2][5][7] ) );
  dp_1 \ANSWER/mem_reg[2][6][7]  ( .ip(n3176), .ck(clk), .q(
        \ANSWER/mem[2][6][7] ) );
  dp_1 \ANSWER/mem_reg[2][7][7]  ( .ip(n3175), .ck(clk), .q(
        \ANSWER/mem[2][7][7] ) );
  dp_1 \ANSWER/mem_reg[2][8][7]  ( .ip(n3174), .ck(clk), .q(
        \ANSWER/mem[2][8][7] ) );
  dp_1 \ANSWER/mem_reg[2][9][7]  ( .ip(n3173), .ck(clk), .q(
        \ANSWER/mem[2][9][7] ) );
  dp_1 \ANSWER/mem_reg[3][0][7]  ( .ip(n3172), .ck(clk), .q(
        \ANSWER/mem[3][0][7] ) );
  dp_1 \ANSWER/mem_reg[3][1][7]  ( .ip(n3171), .ck(clk), .q(
        \ANSWER/mem[3][1][7] ) );
  dp_1 \ANSWER/mem_reg[3][2][7]  ( .ip(n3170), .ck(clk), .q(
        \ANSWER/mem[3][2][7] ) );
  dp_1 \ANSWER/mem_reg[3][3][7]  ( .ip(n3169), .ck(clk), .q(
        \ANSWER/mem[3][3][7] ) );
  dp_1 \ANSWER/mem_reg[3][4][7]  ( .ip(n3168), .ck(clk), .q(
        \ANSWER/mem[3][4][7] ) );
  dp_1 \ANSWER/mem_reg[3][5][7]  ( .ip(n3167), .ck(clk), .q(
        \ANSWER/mem[3][5][7] ) );
  dp_1 \ANSWER/mem_reg[3][6][7]  ( .ip(n3166), .ck(clk), .q(
        \ANSWER/mem[3][6][7] ) );
  dp_1 \ANSWER/mem_reg[3][7][7]  ( .ip(n3165), .ck(clk), .q(
        \ANSWER/mem[3][7][7] ) );
  dp_1 \ANSWER/mem_reg[3][8][7]  ( .ip(n3164), .ck(clk), .q(
        \ANSWER/mem[3][8][7] ) );
  dp_1 \ANSWER/mem_reg[3][9][7]  ( .ip(n3163), .ck(clk), .q(
        \ANSWER/mem[3][9][7] ) );
  dp_1 \ANSWER/mem_reg[4][0][7]  ( .ip(n3162), .ck(clk), .q(
        \ANSWER/mem[4][0][7] ) );
  dp_1 \ANSWER/mem_reg[4][1][7]  ( .ip(n3161), .ck(clk), .q(
        \ANSWER/mem[4][1][7] ) );
  dp_1 \ANSWER/mem_reg[4][2][7]  ( .ip(n3160), .ck(clk), .q(
        \ANSWER/mem[4][2][7] ) );
  dp_1 \ANSWER/mem_reg[4][3][7]  ( .ip(n3159), .ck(clk), .q(
        \ANSWER/mem[4][3][7] ) );
  dp_1 \ANSWER/mem_reg[4][4][7]  ( .ip(n3158), .ck(clk), .q(
        \ANSWER/mem[4][4][7] ) );
  dp_1 \ANSWER/mem_reg[4][5][7]  ( .ip(n3157), .ck(clk), .q(
        \ANSWER/mem[4][5][7] ) );
  dp_1 \ANSWER/mem_reg[4][6][7]  ( .ip(n3156), .ck(clk), .q(
        \ANSWER/mem[4][6][7] ) );
  dp_1 \ANSWER/mem_reg[4][7][7]  ( .ip(n3155), .ck(clk), .q(
        \ANSWER/mem[4][7][7] ) );
  dp_1 \ANSWER/mem_reg[4][8][7]  ( .ip(n3154), .ck(clk), .q(
        \ANSWER/mem[4][8][7] ) );
  dp_1 \ANSWER/mem_reg[4][9][7]  ( .ip(n3153), .ck(clk), .q(
        \ANSWER/mem[4][9][7] ) );
  dp_1 \ANSWER/mem_reg[5][0][7]  ( .ip(n3152), .ck(clk), .q(
        \ANSWER/mem[5][0][7] ) );
  dp_1 \ANSWER/mem_reg[5][1][7]  ( .ip(n3151), .ck(clk), .q(
        \ANSWER/mem[5][1][7] ) );
  dp_1 \ANSWER/mem_reg[5][2][7]  ( .ip(n3150), .ck(clk), .q(
        \ANSWER/mem[5][2][7] ) );
  dp_1 \ANSWER/mem_reg[5][3][7]  ( .ip(n3149), .ck(clk), .q(
        \ANSWER/mem[5][3][7] ) );
  dp_1 \ANSWER/mem_reg[5][4][7]  ( .ip(n3148), .ck(clk), .q(
        \ANSWER/mem[5][4][7] ) );
  dp_1 \ANSWER/mem_reg[5][5][7]  ( .ip(n3147), .ck(clk), .q(
        \ANSWER/mem[5][5][7] ) );
  dp_1 \ANSWER/mem_reg[5][6][7]  ( .ip(n3146), .ck(clk), .q(
        \ANSWER/mem[5][6][7] ) );
  dp_1 \ANSWER/mem_reg[5][7][7]  ( .ip(n3145), .ck(clk), .q(
        \ANSWER/mem[5][7][7] ) );
  dp_1 \ANSWER/mem_reg[5][8][7]  ( .ip(n3144), .ck(clk), .q(
        \ANSWER/mem[5][8][7] ) );
  dp_1 \ANSWER/mem_reg[5][9][7]  ( .ip(n3143), .ck(clk), .q(
        \ANSWER/mem[5][9][7] ) );
  dp_1 \ANSWER/mem_reg[6][0][7]  ( .ip(n3142), .ck(clk), .q(
        \ANSWER/mem[6][0][7] ) );
  dp_1 \ANSWER/mem_reg[6][1][7]  ( .ip(n3141), .ck(clk), .q(
        \ANSWER/mem[6][1][7] ) );
  dp_1 \ANSWER/mem_reg[6][2][7]  ( .ip(n3140), .ck(clk), .q(
        \ANSWER/mem[6][2][7] ) );
  dp_1 \ANSWER/mem_reg[6][3][7]  ( .ip(n3139), .ck(clk), .q(
        \ANSWER/mem[6][3][7] ) );
  dp_1 \ANSWER/mem_reg[6][4][7]  ( .ip(n3138), .ck(clk), .q(
        \ANSWER/mem[6][4][7] ) );
  dp_1 \ANSWER/mem_reg[6][5][7]  ( .ip(n3137), .ck(clk), .q(
        \ANSWER/mem[6][5][7] ) );
  dp_1 \ANSWER/mem_reg[6][6][7]  ( .ip(n3136), .ck(clk), .q(
        \ANSWER/mem[6][6][7] ) );
  dp_1 \ANSWER/mem_reg[6][7][7]  ( .ip(n3135), .ck(clk), .q(
        \ANSWER/mem[6][7][7] ) );
  dp_1 \ANSWER/mem_reg[6][8][7]  ( .ip(n3134), .ck(clk), .q(
        \ANSWER/mem[6][8][7] ) );
  dp_1 \ANSWER/mem_reg[6][9][7]  ( .ip(n3133), .ck(clk), .q(
        \ANSWER/mem[6][9][7] ) );
  dp_1 \ANSWER/mem_reg[7][0][7]  ( .ip(n3132), .ck(clk), .q(
        \ANSWER/mem[7][0][7] ) );
  dp_1 \ANSWER/mem_reg[7][1][7]  ( .ip(n3131), .ck(clk), .q(
        \ANSWER/mem[7][1][7] ) );
  dp_1 \ANSWER/mem_reg[7][2][7]  ( .ip(n3130), .ck(clk), .q(
        \ANSWER/mem[7][2][7] ) );
  dp_1 \ANSWER/mem_reg[7][3][7]  ( .ip(n3129), .ck(clk), .q(
        \ANSWER/mem[7][3][7] ) );
  dp_1 \ANSWER/mem_reg[7][4][7]  ( .ip(n3128), .ck(clk), .q(
        \ANSWER/mem[7][4][7] ) );
  dp_1 \ANSWER/mem_reg[7][5][7]  ( .ip(n3127), .ck(clk), .q(
        \ANSWER/mem[7][5][7] ) );
  dp_1 \ANSWER/mem_reg[7][6][7]  ( .ip(n3126), .ck(clk), .q(
        \ANSWER/mem[7][6][7] ) );
  dp_1 \ANSWER/mem_reg[7][7][7]  ( .ip(n3125), .ck(clk), .q(
        \ANSWER/mem[7][7][7] ) );
  dp_1 \ANSWER/mem_reg[7][8][7]  ( .ip(n3124), .ck(clk), .q(
        \ANSWER/mem[7][8][7] ) );
  dp_1 \ANSWER/mem_reg[7][9][7]  ( .ip(n3123), .ck(clk), .q(
        \ANSWER/mem[7][9][7] ) );
  dp_1 \ANSWER/mem_reg[8][0][7]  ( .ip(n3122), .ck(clk), .q(
        \ANSWER/mem[8][0][7] ) );
  dp_1 \ANSWER/mem_reg[8][1][7]  ( .ip(n3121), .ck(clk), .q(
        \ANSWER/mem[8][1][7] ) );
  dp_1 \ANSWER/mem_reg[8][2][7]  ( .ip(n3120), .ck(clk), .q(
        \ANSWER/mem[8][2][7] ) );
  dp_1 \ANSWER/mem_reg[8][3][7]  ( .ip(n3119), .ck(clk), .q(
        \ANSWER/mem[8][3][7] ) );
  dp_1 \ANSWER/mem_reg[8][4][7]  ( .ip(n3118), .ck(clk), .q(
        \ANSWER/mem[8][4][7] ) );
  dp_1 \ANSWER/mem_reg[8][5][7]  ( .ip(n3117), .ck(clk), .q(
        \ANSWER/mem[8][5][7] ) );
  dp_1 \ANSWER/mem_reg[8][6][7]  ( .ip(n3116), .ck(clk), .q(
        \ANSWER/mem[8][6][7] ) );
  dp_1 \ANSWER/mem_reg[8][7][7]  ( .ip(n3115), .ck(clk), .q(
        \ANSWER/mem[8][7][7] ) );
  dp_1 \ANSWER/mem_reg[8][8][7]  ( .ip(n3114), .ck(clk), .q(
        \ANSWER/mem[8][8][7] ) );
  dp_1 \ANSWER/mem_reg[8][9][7]  ( .ip(n3113), .ck(clk), .q(
        \ANSWER/mem[8][9][7] ) );
  dp_1 \ANSWER/mem_reg[9][0][7]  ( .ip(n3112), .ck(clk), .q(
        \ANSWER/mem[9][0][7] ) );
  dp_1 \ANSWER/mem_reg[9][1][7]  ( .ip(n3111), .ck(clk), .q(
        \ANSWER/mem[9][1][7] ) );
  dp_1 \ANSWER/mem_reg[9][2][7]  ( .ip(n3110), .ck(clk), .q(
        \ANSWER/mem[9][2][7] ) );
  dp_1 \ANSWER/mem_reg[9][3][7]  ( .ip(n3109), .ck(clk), .q(
        \ANSWER/mem[9][3][7] ) );
  dp_1 \ANSWER/mem_reg[9][4][7]  ( .ip(n3108), .ck(clk), .q(
        \ANSWER/mem[9][4][7] ) );
  dp_1 \ANSWER/mem_reg[9][5][7]  ( .ip(n3107), .ck(clk), .q(
        \ANSWER/mem[9][5][7] ) );
  dp_1 \ANSWER/mem_reg[9][6][7]  ( .ip(n3106), .ck(clk), .q(
        \ANSWER/mem[9][6][7] ) );
  dp_1 \ANSWER/mem_reg[9][7][7]  ( .ip(n3105), .ck(clk), .q(
        \ANSWER/mem[9][7][7] ) );
  dp_1 \ANSWER/mem_reg[9][8][7]  ( .ip(n3104), .ck(clk), .q(
        \ANSWER/mem[9][8][7] ) );
  dp_1 \ANSWER/mem_reg[9][9][7]  ( .ip(n3103), .ck(clk), .q(
        \ANSWER/mem[9][9][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][0]  ( .ip(n2302), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][0] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][1]  ( .ip(n2301), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][1] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][2]  ( .ip(n2300), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][2] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][3]  ( .ip(n2299), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][3] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][4]  ( .ip(n2298), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][4] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][5]  ( .ip(n2297), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][5] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][6]  ( .ip(n2296), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][6] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][7]  ( .ip(n2295), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][8]  ( .ip(n2294), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][8] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][9]  ( .ip(n2293), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][9] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][10]  ( .ip(n2292), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][10] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][11]  ( .ip(n2291), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][11] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][12]  ( .ip(n2290), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][12] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][13]  ( .ip(n2289), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][13] ) );
  dp_1 \INPUTSRAM/mem_i_reg[0][14]  ( .ip(n2288), .ck(clk), .q(
        \INPUTSRAM/mem_i[0][14] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][0]  ( .ip(n2287), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][0] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][1]  ( .ip(n2286), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][1] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][2]  ( .ip(n2285), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][2] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][3]  ( .ip(n2284), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][3] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][4]  ( .ip(n2283), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][4] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][5]  ( .ip(n2282), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][5] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][6]  ( .ip(n2281), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][6] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][7]  ( .ip(n2280), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][8]  ( .ip(n2279), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][8] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][9]  ( .ip(n2278), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][9] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][10]  ( .ip(n2277), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][10] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][11]  ( .ip(n2276), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][11] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][12]  ( .ip(n2275), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][12] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][13]  ( .ip(n2274), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][13] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][14]  ( .ip(n2273), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][14] ) );
  dp_1 \INPUTSRAM/mem_i_reg[1][15]  ( .ip(n2272), .ck(clk), .q(
        \INPUTSRAM/mem_i[1][15] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][0]  ( .ip(n2271), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][0] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][1]  ( .ip(n2270), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][1] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][2]  ( .ip(n2269), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][2] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][3]  ( .ip(n2268), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][3] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][4]  ( .ip(n2267), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][4] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][5]  ( .ip(n2266), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][5] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][6]  ( .ip(n2265), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][6] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][7]  ( .ip(n2264), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][8]  ( .ip(n2263), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][8] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][9]  ( .ip(n2262), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][9] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][10]  ( .ip(n2261), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][10] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][11]  ( .ip(n2260), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][11] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][12]  ( .ip(n2259), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][12] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][13]  ( .ip(n2258), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][13] ) );
  dp_1 \INPUTSRAM/mem_i_reg[2][14]  ( .ip(n2257), .ck(clk), .q(
        \INPUTSRAM/mem_i[2][14] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][0]  ( .ip(n2256), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][0] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][1]  ( .ip(n2255), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][1] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][2]  ( .ip(n2254), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][2] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][3]  ( .ip(n2253), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][3] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][4]  ( .ip(n2252), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][4] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][5]  ( .ip(n2251), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][5] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][6]  ( .ip(n2250), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][6] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][7]  ( .ip(n2249), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][8]  ( .ip(n2248), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][8] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][9]  ( .ip(n2247), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][9] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][10]  ( .ip(n2246), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][10] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][11]  ( .ip(n2245), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][11] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][12]  ( .ip(n2244), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][12] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][13]  ( .ip(n2243), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][13] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][14]  ( .ip(n2242), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][14] ) );
  dp_1 \INPUTSRAM/mem_i_reg[3][15]  ( .ip(n2241), .ck(clk), .q(
        \INPUTSRAM/mem_i[3][15] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][0]  ( .ip(n2240), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][0] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][1]  ( .ip(n2239), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][1] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][2]  ( .ip(n2238), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][2] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][3]  ( .ip(n2237), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][3] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][4]  ( .ip(n2236), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][4] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][5]  ( .ip(n2235), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][5] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][6]  ( .ip(n2234), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][6] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][7]  ( .ip(n2233), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][8]  ( .ip(n2232), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][8] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][9]  ( .ip(n2231), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][9] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][10]  ( .ip(n2230), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][10] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][11]  ( .ip(n2229), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][11] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][12]  ( .ip(n2228), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][12] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][13]  ( .ip(n2227), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][13] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][14]  ( .ip(n2226), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][14] ) );
  dp_1 \INPUTSRAM/mem_i_reg[4][15]  ( .ip(n2225), .ck(clk), .q(
        \INPUTSRAM/mem_i[4][15] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][0]  ( .ip(n2224), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][0] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][1]  ( .ip(n2223), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][1] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][2]  ( .ip(n2222), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][2] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][3]  ( .ip(n2221), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][3] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][4]  ( .ip(n2220), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][4] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][5]  ( .ip(n2219), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][5] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][6]  ( .ip(n2218), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][6] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][7]  ( .ip(n2217), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][8]  ( .ip(n2216), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][8] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][9]  ( .ip(n2215), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][9] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][10]  ( .ip(n2214), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][10] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][11]  ( .ip(n2213), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][11] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][12]  ( .ip(n2212), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][12] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][13]  ( .ip(n2211), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][13] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][14]  ( .ip(n2210), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][14] ) );
  dp_1 \INPUTSRAM/mem_i_reg[5][15]  ( .ip(n2209), .ck(clk), .q(
        \INPUTSRAM/mem_i[5][15] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][0]  ( .ip(n2208), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][0] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][1]  ( .ip(n2207), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][1] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][2]  ( .ip(n2206), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][2] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][3]  ( .ip(n2205), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][3] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][4]  ( .ip(n2204), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][4] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][5]  ( .ip(n2203), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][5] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][6]  ( .ip(n2202), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][6] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][7]  ( .ip(n2201), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][8]  ( .ip(n2200), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][8] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][9]  ( .ip(n2199), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][9] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][10]  ( .ip(n2198), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][10] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][11]  ( .ip(n2197), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][11] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][12]  ( .ip(n2196), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][12] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][13]  ( .ip(n2195), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][13] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][14]  ( .ip(n2194), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][14] ) );
  dp_1 \INPUTSRAM/mem_i_reg[6][15]  ( .ip(n2193), .ck(clk), .q(
        \INPUTSRAM/mem_i[6][15] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][0]  ( .ip(n2192), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][0] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][1]  ( .ip(n2191), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][1] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][2]  ( .ip(n2190), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][2] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][3]  ( .ip(n2189), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][3] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][4]  ( .ip(n2188), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][4] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][5]  ( .ip(n2187), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][5] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][6]  ( .ip(n2186), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][6] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][7]  ( .ip(n2185), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][8]  ( .ip(n2184), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][8] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][9]  ( .ip(n2183), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][9] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][10]  ( .ip(n2182), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][10] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][11]  ( .ip(n2181), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][11] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][12]  ( .ip(n2180), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][12] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][13]  ( .ip(n2179), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][13] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][14]  ( .ip(n2178), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][14] ) );
  dp_1 \INPUTSRAM/mem_i_reg[7][15]  ( .ip(n2177), .ck(clk), .q(
        \INPUTSRAM/mem_i[7][15] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][0]  ( .ip(n2176), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][0] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][1]  ( .ip(n2175), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][1] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][2]  ( .ip(n2174), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][2] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][3]  ( .ip(n2173), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][3] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][4]  ( .ip(n2172), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][4] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][5]  ( .ip(n2171), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][5] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][6]  ( .ip(n2170), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][6] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][7]  ( .ip(n2169), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][8]  ( .ip(n2168), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][8] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][9]  ( .ip(n2167), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][9] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][10]  ( .ip(n2166), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][10] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][11]  ( .ip(n2165), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][11] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][12]  ( .ip(n2164), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][12] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][13]  ( .ip(n2163), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][13] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][14]  ( .ip(n2162), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][14] ) );
  dp_1 \INPUTSRAM/mem_i_reg[8][15]  ( .ip(n2161), .ck(clk), .q(
        \INPUTSRAM/mem_i[8][15] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][0]  ( .ip(n2160), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][0] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][1]  ( .ip(n2159), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][1] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][2]  ( .ip(n2158), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][2] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][3]  ( .ip(n2157), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][3] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][4]  ( .ip(n2156), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][4] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][5]  ( .ip(n2155), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][5] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][6]  ( .ip(n2154), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][6] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][7]  ( .ip(n2153), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][7] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][8]  ( .ip(n2152), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][8] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][9]  ( .ip(n2151), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][9] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][10]  ( .ip(n2150), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][10] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][11]  ( .ip(n2149), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][11] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][12]  ( .ip(n2148), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][12] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][13]  ( .ip(n2147), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][13] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][14]  ( .ip(n2146), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][14] ) );
  dp_1 \INPUTSRAM/mem_i_reg[9][15]  ( .ip(n2145), .ck(clk), .q(
        \INPUTSRAM/mem_i[9][15] ) );
  dp_1 \WEIGHT_2/q_reg[14]  ( .ip(n2130), .ck(clk), .q(q_w2[14]) );
  dp_1 \WEIGHT_2/q_reg[15]  ( .ip(n2129), .ck(clk), .q(q_w2[15]) );
  dp_1 \ROUTEDATA/regData_reg[8]  ( .ip(n2128), .ck(clk), .q(
        \ROUTEDATA/regData [8]) );
  dp_1 \ROUTEDATA/regData_reg[24]  ( .ip(n2127), .ck(clk), .q(
        \ROUTEDATA/regData [24]) );
  dp_1 \ROUTEDATA/regData_reg[40]  ( .ip(n2126), .ck(clk), .q(
        \ROUTEDATA/regData [40]) );
  dp_1 \ROUTEDATA/regData_reg[56]  ( .ip(n2125), .ck(clk), .q(
        \ROUTEDATA/regData [56]) );
  dp_1 \ROUTEDATA/regData_reg[72]  ( .ip(n2124), .ck(clk), .q(
        \ROUTEDATA/regData [72]) );
  dp_1 \ROUTEDATA/regData_reg[88]  ( .ip(n2123), .ck(clk), .q(
        \ROUTEDATA/regData [88]) );
  dp_1 \ROUTEDATA/regData_reg[104]  ( .ip(n2122), .ck(clk), .q(
        \ROUTEDATA/regData [104]) );
  dp_1 \ROUTEDATA/regData_reg[120]  ( .ip(n2121), .ck(clk), .q(
        \ROUTEDATA/regData [120]) );
  dp_1 \ROUTEDATA/regData_reg[136]  ( .ip(n2120), .ck(clk), .q(
        \ROUTEDATA/regData [136]) );
  dp_1 \ROUTEDATA/regData_reg[152]  ( .ip(n2119), .ck(clk), .q(
        \ROUTEDATA/regData [152]) );
  dp_1 \ROUTEDATA/regData_reg[9]  ( .ip(n2118), .ck(clk), .q(
        \ROUTEDATA/regData [9]) );
  dp_1 \ROUTEDATA/regData_reg[25]  ( .ip(n2117), .ck(clk), .q(
        \ROUTEDATA/regData [25]) );
  dp_1 \ROUTEDATA/regData_reg[41]  ( .ip(n2116), .ck(clk), .q(
        \ROUTEDATA/regData [41]) );
  dp_1 \ROUTEDATA/regData_reg[57]  ( .ip(n2115), .ck(clk), .q(
        \ROUTEDATA/regData [57]) );
  dp_1 \ROUTEDATA/regData_reg[73]  ( .ip(n2114), .ck(clk), .q(
        \ROUTEDATA/regData [73]) );
  dp_1 \ROUTEDATA/regData_reg[89]  ( .ip(n2113), .ck(clk), .q(
        \ROUTEDATA/regData [89]) );
  dp_1 \ROUTEDATA/regData_reg[105]  ( .ip(n2112), .ck(clk), .q(
        \ROUTEDATA/regData [105]) );
  dp_1 \ROUTEDATA/regData_reg[121]  ( .ip(n2111), .ck(clk), .q(
        \ROUTEDATA/regData [121]) );
  dp_1 \ROUTEDATA/regData_reg[137]  ( .ip(n2110), .ck(clk), .q(
        \ROUTEDATA/regData [137]) );
  dp_1 \ROUTEDATA/regData_reg[153]  ( .ip(n2109), .ck(clk), .q(
        \ROUTEDATA/regData [153]) );
  dp_1 \ROUTEDATA/regData_reg[10]  ( .ip(n2108), .ck(clk), .q(
        \ROUTEDATA/regData [10]) );
  dp_1 \ROUTEDATA/regData_reg[26]  ( .ip(n2107), .ck(clk), .q(
        \ROUTEDATA/regData [26]) );
  dp_1 \ROUTEDATA/regData_reg[42]  ( .ip(n2106), .ck(clk), .q(
        \ROUTEDATA/regData [42]) );
  dp_1 \ROUTEDATA/regData_reg[58]  ( .ip(n2105), .ck(clk), .q(
        \ROUTEDATA/regData [58]) );
  dp_1 \ROUTEDATA/regData_reg[74]  ( .ip(n2104), .ck(clk), .q(
        \ROUTEDATA/regData [74]) );
  dp_1 \ROUTEDATA/regData_reg[90]  ( .ip(n2103), .ck(clk), .q(
        \ROUTEDATA/regData [90]) );
  dp_1 \ROUTEDATA/regData_reg[106]  ( .ip(n2102), .ck(clk), .q(
        \ROUTEDATA/regData [106]) );
  dp_1 \ROUTEDATA/regData_reg[122]  ( .ip(n2101), .ck(clk), .q(
        \ROUTEDATA/regData [122]) );
  dp_1 \ROUTEDATA/regData_reg[138]  ( .ip(n2100), .ck(clk), .q(
        \ROUTEDATA/regData [138]) );
  dp_1 \ROUTEDATA/regData_reg[154]  ( .ip(n2099), .ck(clk), .q(
        \ROUTEDATA/regData [154]) );
  dp_1 \ROUTEDATA/regData_reg[11]  ( .ip(n2098), .ck(clk), .q(
        \ROUTEDATA/regData [11]) );
  dp_1 \ROUTEDATA/regData_reg[27]  ( .ip(n2097), .ck(clk), .q(
        \ROUTEDATA/regData [27]) );
  dp_1 \ROUTEDATA/regData_reg[43]  ( .ip(n2096), .ck(clk), .q(
        \ROUTEDATA/regData [43]) );
  dp_1 \ROUTEDATA/regData_reg[59]  ( .ip(n2095), .ck(clk), .q(
        \ROUTEDATA/regData [59]) );
  dp_1 \ROUTEDATA/regData_reg[75]  ( .ip(n2094), .ck(clk), .q(
        \ROUTEDATA/regData [75]) );
  dp_1 \ROUTEDATA/regData_reg[91]  ( .ip(n2093), .ck(clk), .q(
        \ROUTEDATA/regData [91]) );
  dp_1 \ROUTEDATA/regData_reg[107]  ( .ip(n2092), .ck(clk), .q(
        \ROUTEDATA/regData [107]) );
  dp_1 \ROUTEDATA/regData_reg[123]  ( .ip(n2091), .ck(clk), .q(
        \ROUTEDATA/regData [123]) );
  dp_1 \ROUTEDATA/regData_reg[139]  ( .ip(n2090), .ck(clk), .q(
        \ROUTEDATA/regData [139]) );
  dp_1 \ROUTEDATA/regData_reg[155]  ( .ip(n2089), .ck(clk), .q(
        \ROUTEDATA/regData [155]) );
  dp_1 \ROUTEDATA/regData_reg[12]  ( .ip(n2088), .ck(clk), .q(
        \ROUTEDATA/regData [12]) );
  dp_1 \ROUTEDATA/regData_reg[28]  ( .ip(n2087), .ck(clk), .q(
        \ROUTEDATA/regData [28]) );
  dp_1 \ROUTEDATA/regData_reg[44]  ( .ip(n2086), .ck(clk), .q(
        \ROUTEDATA/regData [44]) );
  dp_1 \ROUTEDATA/regData_reg[60]  ( .ip(n2085), .ck(clk), .q(
        \ROUTEDATA/regData [60]) );
  dp_1 \ROUTEDATA/regData_reg[76]  ( .ip(n2084), .ck(clk), .q(
        \ROUTEDATA/regData [76]) );
  dp_1 \ROUTEDATA/regData_reg[92]  ( .ip(n2083), .ck(clk), .q(
        \ROUTEDATA/regData [92]) );
  dp_1 \ROUTEDATA/regData_reg[108]  ( .ip(n2082), .ck(clk), .q(
        \ROUTEDATA/regData [108]) );
  dp_1 \ROUTEDATA/regData_reg[124]  ( .ip(n2081), .ck(clk), .q(
        \ROUTEDATA/regData [124]) );
  dp_1 \ROUTEDATA/regData_reg[140]  ( .ip(n2080), .ck(clk), .q(
        \ROUTEDATA/regData [140]) );
  dp_1 \ROUTEDATA/regData_reg[156]  ( .ip(n2079), .ck(clk), .q(
        \ROUTEDATA/regData [156]) );
  dp_1 \ROUTEDATA/regData_reg[13]  ( .ip(n2078), .ck(clk), .q(
        \ROUTEDATA/regData [13]) );
  dp_1 \ROUTEDATA/regData_reg[29]  ( .ip(n2077), .ck(clk), .q(
        \ROUTEDATA/regData [29]) );
  dp_1 \ROUTEDATA/regData_reg[45]  ( .ip(n2076), .ck(clk), .q(
        \ROUTEDATA/regData [45]) );
  dp_1 \ROUTEDATA/regData_reg[61]  ( .ip(n2075), .ck(clk), .q(
        \ROUTEDATA/regData [61]) );
  dp_1 \ROUTEDATA/regData_reg[77]  ( .ip(n2074), .ck(clk), .q(
        \ROUTEDATA/regData [77]) );
  dp_1 \ROUTEDATA/regData_reg[93]  ( .ip(n2073), .ck(clk), .q(
        \ROUTEDATA/regData [93]) );
  dp_1 \ROUTEDATA/regData_reg[109]  ( .ip(n2072), .ck(clk), .q(
        \ROUTEDATA/regData [109]) );
  dp_1 \ROUTEDATA/regData_reg[125]  ( .ip(n2071), .ck(clk), .q(
        \ROUTEDATA/regData [125]) );
  dp_1 \ROUTEDATA/regData_reg[141]  ( .ip(n2070), .ck(clk), .q(
        \ROUTEDATA/regData [141]) );
  dp_1 \ROUTEDATA/regData_reg[157]  ( .ip(n2069), .ck(clk), .q(
        \ROUTEDATA/regData [157]) );
  dp_1 \ROUTEDATA/regData_reg[14]  ( .ip(n2068), .ck(clk), .q(
        \ROUTEDATA/regData [14]) );
  dp_1 \ROUTEDATA/regData_reg[30]  ( .ip(n2067), .ck(clk), .q(
        \ROUTEDATA/regData [30]) );
  dp_1 \ROUTEDATA/regData_reg[46]  ( .ip(n2066), .ck(clk), .q(
        \ROUTEDATA/regData [46]) );
  dp_1 \ROUTEDATA/regData_reg[62]  ( .ip(n2065), .ck(clk), .q(
        \ROUTEDATA/regData [62]) );
  dp_1 \ROUTEDATA/regData_reg[78]  ( .ip(n2064), .ck(clk), .q(
        \ROUTEDATA/regData [78]) );
  dp_1 \ROUTEDATA/regData_reg[94]  ( .ip(n2063), .ck(clk), .q(
        \ROUTEDATA/regData [94]) );
  dp_1 \ROUTEDATA/regData_reg[110]  ( .ip(n2062), .ck(clk), .q(
        \ROUTEDATA/regData [110]) );
  dp_1 \ROUTEDATA/regData_reg[126]  ( .ip(n2061), .ck(clk), .q(
        \ROUTEDATA/regData [126]) );
  dp_1 \ROUTEDATA/regData_reg[142]  ( .ip(n2060), .ck(clk), .q(
        \ROUTEDATA/regData [142]) );
  dp_1 \ROUTEDATA/regData_reg[158]  ( .ip(n2059), .ck(clk), .q(
        \ROUTEDATA/regData [158]) );
  dp_1 \ROUTEDATA/regData_reg[15]  ( .ip(n2058), .ck(clk), .q(
        \ROUTEDATA/regData [15]) );
  dp_1 \ROUTEDATA/regData_reg[31]  ( .ip(n2057), .ck(clk), .q(
        \ROUTEDATA/regData [31]) );
  dp_1 \ROUTEDATA/regData_reg[47]  ( .ip(n2056), .ck(clk), .q(
        \ROUTEDATA/regData [47]) );
  dp_1 \ROUTEDATA/regData_reg[63]  ( .ip(n2055), .ck(clk), .q(
        \ROUTEDATA/regData [63]) );
  dp_1 \ROUTEDATA/regData_reg[79]  ( .ip(n2054), .ck(clk), .q(
        \ROUTEDATA/regData [79]) );
  dp_1 \ROUTEDATA/regData_reg[95]  ( .ip(n2053), .ck(clk), .q(
        \ROUTEDATA/regData [95]) );
  dp_1 \ROUTEDATA/regData_reg[111]  ( .ip(n2052), .ck(clk), .q(
        \ROUTEDATA/regData [111]) );
  dp_1 \ROUTEDATA/regData_reg[127]  ( .ip(n2051), .ck(clk), .q(
        \ROUTEDATA/regData [127]) );
  dp_1 \ROUTEDATA/regData_reg[143]  ( .ip(n2050), .ck(clk), .q(
        \ROUTEDATA/regData [143]) );
  dp_1 \ROUTEDATA/regData_reg[159]  ( .ip(n2049), .ck(clk), .q(
        \ROUTEDATA/regData [159]) );
  dp_1 \ROUTEDATA/regData_reg[0]  ( .ip(n2048), .ck(clk), .q(
        \ROUTEDATA/regData [0]) );
  dp_1 \ROUTEDATA/regData_reg[16]  ( .ip(n2047), .ck(clk), .q(
        \ROUTEDATA/regData [16]) );
  dp_1 \ROUTEDATA/regData_reg[32]  ( .ip(n2046), .ck(clk), .q(
        \ROUTEDATA/regData [32]) );
  dp_1 \ROUTEDATA/regData_reg[48]  ( .ip(n2045), .ck(clk), .q(
        \ROUTEDATA/regData [48]) );
  dp_1 \ROUTEDATA/regData_reg[64]  ( .ip(n2044), .ck(clk), .q(
        \ROUTEDATA/regData [64]) );
  dp_1 \ROUTEDATA/regData_reg[80]  ( .ip(n2043), .ck(clk), .q(
        \ROUTEDATA/regData [80]) );
  dp_1 \ROUTEDATA/regData_reg[96]  ( .ip(n2042), .ck(clk), .q(
        \ROUTEDATA/regData [96]) );
  dp_1 \ROUTEDATA/regData_reg[112]  ( .ip(n2041), .ck(clk), .q(
        \ROUTEDATA/regData [112]) );
  dp_1 \ROUTEDATA/regData_reg[128]  ( .ip(n2040), .ck(clk), .q(
        \ROUTEDATA/regData [128]) );
  dp_1 \ROUTEDATA/regData_reg[144]  ( .ip(n2039), .ck(clk), .q(
        \ROUTEDATA/regData [144]) );
  dp_1 \ROUTEDATA/regData_reg[1]  ( .ip(n2038), .ck(clk), .q(
        \ROUTEDATA/regData [1]) );
  dp_1 \ROUTEDATA/regData_reg[17]  ( .ip(n2037), .ck(clk), .q(
        \ROUTEDATA/regData [17]) );
  dp_1 \ROUTEDATA/regData_reg[33]  ( .ip(n2036), .ck(clk), .q(
        \ROUTEDATA/regData [33]) );
  dp_1 \ROUTEDATA/regData_reg[49]  ( .ip(n2035), .ck(clk), .q(
        \ROUTEDATA/regData [49]) );
  dp_1 \ROUTEDATA/regData_reg[65]  ( .ip(n2034), .ck(clk), .q(
        \ROUTEDATA/regData [65]) );
  dp_1 \ROUTEDATA/regData_reg[81]  ( .ip(n2033), .ck(clk), .q(
        \ROUTEDATA/regData [81]) );
  dp_1 \ROUTEDATA/regData_reg[97]  ( .ip(n2032), .ck(clk), .q(
        \ROUTEDATA/regData [97]) );
  dp_1 \ROUTEDATA/regData_reg[113]  ( .ip(n2031), .ck(clk), .q(
        \ROUTEDATA/regData [113]) );
  dp_1 \ROUTEDATA/regData_reg[129]  ( .ip(n2030), .ck(clk), .q(
        \ROUTEDATA/regData [129]) );
  dp_1 \ROUTEDATA/regData_reg[145]  ( .ip(n2029), .ck(clk), .q(
        \ROUTEDATA/regData [145]) );
  dp_1 \ROUTEDATA/regData_reg[2]  ( .ip(n2028), .ck(clk), .q(
        \ROUTEDATA/regData [2]) );
  dp_1 \ROUTEDATA/regData_reg[18]  ( .ip(n2027), .ck(clk), .q(
        \ROUTEDATA/regData [18]) );
  dp_1 \ROUTEDATA/regData_reg[34]  ( .ip(n2026), .ck(clk), .q(
        \ROUTEDATA/regData [34]) );
  dp_1 \ROUTEDATA/regData_reg[50]  ( .ip(n2025), .ck(clk), .q(
        \ROUTEDATA/regData [50]) );
  dp_1 \ROUTEDATA/regData_reg[66]  ( .ip(n2024), .ck(clk), .q(
        \ROUTEDATA/regData [66]) );
  dp_1 \ROUTEDATA/regData_reg[82]  ( .ip(n2023), .ck(clk), .q(
        \ROUTEDATA/regData [82]) );
  dp_1 \ROUTEDATA/regData_reg[98]  ( .ip(n2022), .ck(clk), .q(
        \ROUTEDATA/regData [98]) );
  dp_1 \ROUTEDATA/regData_reg[114]  ( .ip(n2021), .ck(clk), .q(
        \ROUTEDATA/regData [114]) );
  dp_1 \ROUTEDATA/regData_reg[130]  ( .ip(n2020), .ck(clk), .q(
        \ROUTEDATA/regData [130]) );
  dp_1 \ROUTEDATA/regData_reg[146]  ( .ip(n2019), .ck(clk), .q(
        \ROUTEDATA/regData [146]) );
  dp_1 \ROUTEDATA/regData_reg[3]  ( .ip(n2018), .ck(clk), .q(
        \ROUTEDATA/regData [3]) );
  dp_1 \ROUTEDATA/regData_reg[19]  ( .ip(n2017), .ck(clk), .q(
        \ROUTEDATA/regData [19]) );
  dp_1 \ROUTEDATA/regData_reg[35]  ( .ip(n2016), .ck(clk), .q(
        \ROUTEDATA/regData [35]) );
  dp_1 \ROUTEDATA/regData_reg[51]  ( .ip(n2015), .ck(clk), .q(
        \ROUTEDATA/regData [51]) );
  dp_1 \ROUTEDATA/regData_reg[67]  ( .ip(n2014), .ck(clk), .q(
        \ROUTEDATA/regData [67]) );
  dp_1 \ROUTEDATA/regData_reg[83]  ( .ip(n2013), .ck(clk), .q(
        \ROUTEDATA/regData [83]) );
  dp_1 \ROUTEDATA/regData_reg[99]  ( .ip(n2012), .ck(clk), .q(
        \ROUTEDATA/regData [99]) );
  dp_1 \ROUTEDATA/regData_reg[115]  ( .ip(n2011), .ck(clk), .q(
        \ROUTEDATA/regData [115]) );
  dp_1 \ROUTEDATA/regData_reg[131]  ( .ip(n2010), .ck(clk), .q(
        \ROUTEDATA/regData [131]) );
  dp_1 \ROUTEDATA/regData_reg[147]  ( .ip(n2009), .ck(clk), .q(
        \ROUTEDATA/regData [147]) );
  dp_1 \ROUTEDATA/regData_reg[4]  ( .ip(n2008), .ck(clk), .q(
        \ROUTEDATA/regData [4]) );
  dp_1 \ROUTEDATA/regData_reg[20]  ( .ip(n2007), .ck(clk), .q(
        \ROUTEDATA/regData [20]) );
  dp_1 \ROUTEDATA/regData_reg[36]  ( .ip(n2006), .ck(clk), .q(
        \ROUTEDATA/regData [36]) );
  dp_1 \ROUTEDATA/regData_reg[52]  ( .ip(n2005), .ck(clk), .q(
        \ROUTEDATA/regData [52]) );
  dp_1 \ROUTEDATA/regData_reg[68]  ( .ip(n2004), .ck(clk), .q(
        \ROUTEDATA/regData [68]) );
  dp_1 \ROUTEDATA/regData_reg[84]  ( .ip(n2003), .ck(clk), .q(
        \ROUTEDATA/regData [84]) );
  dp_1 \ROUTEDATA/regData_reg[100]  ( .ip(n2002), .ck(clk), .q(
        \ROUTEDATA/regData [100]) );
  dp_1 \ROUTEDATA/regData_reg[116]  ( .ip(n2001), .ck(clk), .q(
        \ROUTEDATA/regData [116]) );
  dp_1 \ROUTEDATA/regData_reg[132]  ( .ip(n2000), .ck(clk), .q(
        \ROUTEDATA/regData [132]) );
  dp_1 \ROUTEDATA/regData_reg[148]  ( .ip(n1999), .ck(clk), .q(
        \ROUTEDATA/regData [148]) );
  dp_1 \ROUTEDATA/regData_reg[5]  ( .ip(n1998), .ck(clk), .q(
        \ROUTEDATA/regData [5]) );
  dp_1 \ROUTEDATA/regData_reg[21]  ( .ip(n1997), .ck(clk), .q(
        \ROUTEDATA/regData [21]) );
  dp_1 \ROUTEDATA/regData_reg[37]  ( .ip(n1996), .ck(clk), .q(
        \ROUTEDATA/regData [37]) );
  dp_1 \ROUTEDATA/regData_reg[53]  ( .ip(n1995), .ck(clk), .q(
        \ROUTEDATA/regData [53]) );
  dp_1 \ROUTEDATA/regData_reg[69]  ( .ip(n1994), .ck(clk), .q(
        \ROUTEDATA/regData [69]) );
  dp_1 \ROUTEDATA/regData_reg[85]  ( .ip(n1993), .ck(clk), .q(
        \ROUTEDATA/regData [85]) );
  dp_1 \ROUTEDATA/regData_reg[101]  ( .ip(n1992), .ck(clk), .q(
        \ROUTEDATA/regData [101]) );
  dp_1 \ROUTEDATA/regData_reg[117]  ( .ip(n1991), .ck(clk), .q(
        \ROUTEDATA/regData [117]) );
  dp_1 \ROUTEDATA/regData_reg[133]  ( .ip(n1990), .ck(clk), .q(
        \ROUTEDATA/regData [133]) );
  dp_1 \ROUTEDATA/regData_reg[149]  ( .ip(n1989), .ck(clk), .q(
        \ROUTEDATA/regData [149]) );
  dp_1 \ROUTEDATA/regData_reg[6]  ( .ip(n1988), .ck(clk), .q(
        \ROUTEDATA/regData [6]) );
  dp_1 \ROUTEDATA/regData_reg[22]  ( .ip(n1987), .ck(clk), .q(
        \ROUTEDATA/regData [22]) );
  dp_1 \ROUTEDATA/regData_reg[38]  ( .ip(n1986), .ck(clk), .q(
        \ROUTEDATA/regData [38]) );
  dp_1 \ROUTEDATA/regData_reg[54]  ( .ip(n1985), .ck(clk), .q(
        \ROUTEDATA/regData [54]) );
  dp_1 \ROUTEDATA/regData_reg[70]  ( .ip(n1984), .ck(clk), .q(
        \ROUTEDATA/regData [70]) );
  dp_1 \ROUTEDATA/regData_reg[86]  ( .ip(n1983), .ck(clk), .q(
        \ROUTEDATA/regData [86]) );
  dp_1 \ROUTEDATA/regData_reg[102]  ( .ip(n1982), .ck(clk), .q(
        \ROUTEDATA/regData [102]) );
  dp_1 \ROUTEDATA/regData_reg[118]  ( .ip(n1981), .ck(clk), .q(
        \ROUTEDATA/regData [118]) );
  dp_1 \ROUTEDATA/regData_reg[134]  ( .ip(n1980), .ck(clk), .q(
        \ROUTEDATA/regData [134]) );
  dp_1 \ROUTEDATA/regData_reg[150]  ( .ip(n1979), .ck(clk), .q(
        \ROUTEDATA/regData [150]) );
  dp_1 \ROUTEDATA/regData_reg[7]  ( .ip(n1978), .ck(clk), .q(
        \ROUTEDATA/regData [7]) );
  dp_1 \ROUTEDATA/regData_reg[23]  ( .ip(n1977), .ck(clk), .q(
        \ROUTEDATA/regData [23]) );
  dp_1 \ROUTEDATA/regData_reg[39]  ( .ip(n1976), .ck(clk), .q(
        \ROUTEDATA/regData [39]) );
  dp_1 \ROUTEDATA/regData_reg[55]  ( .ip(n1975), .ck(clk), .q(
        \ROUTEDATA/regData [55]) );
  dp_1 \ROUTEDATA/regData_reg[71]  ( .ip(n1974), .ck(clk), .q(
        \ROUTEDATA/regData [71]) );
  dp_1 \ROUTEDATA/regData_reg[87]  ( .ip(n1973), .ck(clk), .q(
        \ROUTEDATA/regData [87]) );
  dp_1 \ROUTEDATA/regData_reg[103]  ( .ip(n1972), .ck(clk), .q(
        \ROUTEDATA/regData [103]) );
  dp_1 \ROUTEDATA/regData_reg[119]  ( .ip(n1971), .ck(clk), .q(
        \ROUTEDATA/regData [119]) );
  dp_1 \ROUTEDATA/regData_reg[135]  ( .ip(n1970), .ck(clk), .q(
        \ROUTEDATA/regData [135]) );
  dp_1 \ROUTEDATA/regData_reg[151]  ( .ip(n1969), .ck(clk), .q(
        \ROUTEDATA/regData [151]) );
  dp_1 \STAGE_1/weightReg_reg[15]  ( .ip(weight1[15]), .ck(clk), .q(
        \STAGE_1/weightReg [15]) );
  dp_1 \INPUTSRAM/q_reg[23]  ( .ip(\INPUTSRAM/mem_i[1][7] ), .ck(clk), .q(
        m1Inputs[23]) );
  dp_1 \INPUTSRAM/q_reg[24]  ( .ip(\INPUTSRAM/mem_i[1][8] ), .ck(clk), .q(
        m1Inputs[24]) );
  dp_1 \INPUTSRAM/q_reg[133]  ( .ip(\INPUTSRAM/mem_i[8][5] ), .ck(clk), .q(
        m1Inputs[133]) );
  dp_1 \INPUTSRAM/q_reg[37]  ( .ip(\INPUTSRAM/mem_i[2][5] ), .ck(clk), .q(
        m1Inputs[37]) );
  dp_1 \INPUTSRAM/q_reg[96]  ( .ip(\INPUTSRAM/mem_i[6][0] ), .ck(clk), .q(
        m1Inputs[96]) );
  dp_1 \INPUTSRAM/q_reg[101]  ( .ip(\INPUTSRAM/mem_i[6][5] ), .ck(clk), .q(
        m1Inputs[101]) );
  dp_1 \STAGE_1/weightReg_reg[6]  ( .ip(weight1[6]), .ck(clk), .q(
        \STAGE_1/weightReg [6]) );
  dp_1 \STAGE_1/weightReg_reg[3]  ( .ip(weight1[3]), .ck(clk), .q(
        \STAGE_1/weightReg [3]) );
  dp_1 \STAGE_1/weightReg_reg[7]  ( .ip(weight1[7]), .ck(clk), .q(
        \STAGE_1/weightReg [7]) );
  dp_1 \INPUTSRAM/q_reg[19]  ( .ip(\INPUTSRAM/mem_i[1][3] ), .ck(clk), .q(
        m1Inputs[19]) );
  dp_1 \WEIGHT_2/q_reg[13]  ( .ip(n2131), .ck(clk), .q(q_w2[13]) );
  dp_1 \WEIGHT_2/q_reg[12]  ( .ip(n2132), .ck(clk), .q(q_w2[12]) );
  dp_1 \INPUTSRAM/q_reg[22]  ( .ip(\INPUTSRAM/mem_i[1][6] ), .ck(clk), .q(
        m1Inputs[22]) );
  dp_1 \WEIGHT_2/q_reg[10]  ( .ip(n2134), .ck(clk), .q(q_w2[10]) );
  dp_1 \INPUTSRAM/q_reg[157]  ( .ip(\INPUTSRAM/mem_i[9][13] ), .ck(clk), .q(
        m1Inputs[157]) );
  dp_1 \INPUTSRAM/q_reg[156]  ( .ip(\INPUTSRAM/mem_i[9][12] ), .ck(clk), .q(
        m1Inputs[156]) );
  dp_1 \WEIGHT_2/q_reg[11]  ( .ip(n2133), .ck(clk), .q(q_w2[11]) );
  dp_1 \INPUTSRAM/q_reg[140]  ( .ip(\INPUTSRAM/mem_i[8][12] ), .ck(clk), .q(
        m1Inputs[140]) );
  dp_1 \INPUTSRAM/q_reg[150]  ( .ip(\INPUTSRAM/mem_i[9][6] ), .ck(clk), .q(
        m1Inputs[150]) );
  dp_1 \INPUTSRAM/q_reg[141]  ( .ip(\INPUTSRAM/mem_i[8][13] ), .ck(clk), .q(
        m1Inputs[141]) );
  dp_1 \INPUTSRAM/q_reg[134]  ( .ip(\INPUTSRAM/mem_i[8][6] ), .ck(clk), .q(
        m1Inputs[134]) );
  dp_1 \INPUTSRAM/q_reg[26]  ( .ip(\INPUTSRAM/mem_i[1][10] ), .ck(clk), .q(
        m1Inputs[26]) );
  dp_1 \INPUTSRAM/q_reg[155]  ( .ip(\INPUTSRAM/mem_i[9][11] ), .ck(clk), .q(
        m1Inputs[155]) );
  dp_1 \INPUTSRAM/q_reg[27]  ( .ip(\INPUTSRAM/mem_i[1][11] ), .ck(clk), .q(
        m1Inputs[27]) );
  dp_1 \INPUTSRAM/q_reg[25]  ( .ip(\INPUTSRAM/mem_i[1][9] ), .ck(clk), .q(
        m1Inputs[25]) );
  dp_1 \WEIGHT_2/q_reg[9]  ( .ip(n2135), .ck(clk), .q(q_w2[9]) );
  dp_1 \INPUTSRAM/q_reg[139]  ( .ip(\INPUTSRAM/mem_i[8][11] ), .ck(clk), .q(
        m1Inputs[139]) );
  dp_1 \WEIGHT_2/q_reg[8]  ( .ip(n2136), .ck(clk), .q(q_w2[8]) );
  dp_1 \INPUTSRAM/q_reg[28]  ( .ip(\INPUTSRAM/mem_i[1][12] ), .ck(clk), .q(
        m1Inputs[28]) );
  dp_1 \INPUTSRAM/q_reg[154]  ( .ip(\INPUTSRAM/mem_i[9][10] ), .ck(clk), .q(
        m1Inputs[154]) );
  dp_1 \INPUTSRAM/q_reg[153]  ( .ip(\INPUTSRAM/mem_i[9][9] ), .ck(clk), .q(
        m1Inputs[153]) );
  dp_1 \INPUTSRAM/q_reg[51]  ( .ip(\INPUTSRAM/mem_i[3][3] ), .ck(clk), .q(
        m1Inputs[51]) );
  dp_1 \WEIGHT_2/q_reg[7]  ( .ip(n2137), .ck(clk), .q(q_w2[7]) );
  dp_1 \INPUTSRAM/q_reg[138]  ( .ip(\INPUTSRAM/mem_i[8][10] ), .ck(clk), .q(
        m1Inputs[138]) );
  dp_1 \INPUTSRAM/q_reg[137]  ( .ip(\INPUTSRAM/mem_i[8][9] ), .ck(clk), .q(
        m1Inputs[137]) );
  dp_1 \INPUTSRAM/q_reg[124]  ( .ip(\INPUTSRAM/mem_i[7][12] ), .ck(clk), .q(
        m1Inputs[124]) );
  dp_1 \INPUTSRAM/q_reg[3]  ( .ip(\INPUTSRAM/mem_i[0][3] ), .ck(clk), .q(
        m1Inputs[3]) );
  dp_1 \INPUTSRAM/q_reg[6]  ( .ip(\INPUTSRAM/mem_i[0][6] ), .ck(clk), .q(
        m1Inputs[6]) );
  dp_1 \INPUTSRAM/q_reg[131]  ( .ip(\INPUTSRAM/mem_i[8][3] ), .ck(clk), .q(
        m1Inputs[131]) );
  dp_1 \WEIGHT_2/q_reg[6]  ( .ip(n2138), .ck(clk), .q(q_w2[6]) );
  dp_1 \INPUTSRAM/q_reg[54]  ( .ip(\INPUTSRAM/mem_i[3][6] ), .ck(clk), .q(
        m1Inputs[54]) );
  dp_1 \INPUTSRAM/q_reg[118]  ( .ip(\INPUTSRAM/mem_i[7][6] ), .ck(clk), .q(
        m1Inputs[118]) );
  dp_1 \INPUTSRAM/q_reg[146]  ( .ip(\INPUTSRAM/mem_i[9][2] ), .ck(clk), .q(
        m1Inputs[146]) );
  dp_1 \WEIGHT_2/q_reg[5]  ( .ip(n2139), .ck(clk), .q(q_w2[5]) );
  dp_1 \INPUTSRAM/q_reg[115]  ( .ip(\INPUTSRAM/mem_i[7][3] ), .ck(clk), .q(
        m1Inputs[115]) );
  dp_1 \INPUTSRAM/q_reg[70]  ( .ip(\INPUTSRAM/mem_i[4][6] ), .ck(clk), .q(
        m1Inputs[70]) );
  dp_1 \INPUTSRAM/q_reg[130]  ( .ip(\INPUTSRAM/mem_i[8][2] ), .ck(clk), .q(
        m1Inputs[130]) );
  dp_1 \INPUTSRAM/q_reg[83]  ( .ip(\INPUTSRAM/mem_i[5][3] ), .ck(clk), .q(
        m1Inputs[83]) );
  dp_1 \INPUTSRAM/q_reg[64]  ( .ip(\INPUTSRAM/mem_i[4][0] ), .ck(clk), .q(
        m1Inputs[64]) );
  dp_1 \INPUTSRAM/q_reg[99]  ( .ip(\INPUTSRAM/mem_i[6][3] ), .ck(clk), .q(
        m1Inputs[99]) );
  dp_1 \INPUTSRAM/q_reg[86]  ( .ip(\INPUTSRAM/mem_i[5][6] ), .ck(clk), .q(
        m1Inputs[86]) );
  dp_1 \INPUTSRAM/q_reg[18]  ( .ip(\INPUTSRAM/mem_i[1][2] ), .ck(clk), .q(
        m1Inputs[18]) );
  dp_1 \INPUTSRAM/q_reg[102]  ( .ip(\INPUTSRAM/mem_i[6][6] ), .ck(clk), .q(
        m1Inputs[102]) );
  dp_1 \INPUTSRAM/q_reg[80]  ( .ip(\INPUTSRAM/mem_i[5][0] ), .ck(clk), .q(
        m1Inputs[80]) );
  dp_1 \INPUTSRAM/q_reg[123]  ( .ip(\INPUTSRAM/mem_i[7][11] ), .ck(clk), .q(
        m1Inputs[123]) );
  dp_1 \INPUTSRAM/q_reg[147]  ( .ip(\INPUTSRAM/mem_i[9][3] ), .ck(clk), .q(
        m1Inputs[147]) );
  dp_1 \INPUTSRAM/q_reg[62]  ( .ip(\INPUTSRAM/mem_i[3][14] ), .ck(clk), .q(
        m1Inputs[62]) );
  dp_1 \WEIGHT_2/q_reg[2]  ( .ip(n2142), .ck(clk), .q(q_w2[2]) );
  dp_1 \INPUTSRAM/q_reg[112]  ( .ip(\INPUTSRAM/mem_i[7][0] ), .ck(clk), .q(
        m1Inputs[112]) );
  dp_1 \INPUTSRAM/q_reg[67]  ( .ip(\INPUTSRAM/mem_i[4][3] ), .ck(clk), .q(
        m1Inputs[67]) );
  dp_1 \INPUTSRAM/q_reg[13]  ( .ip(\INPUTSRAM/mem_i[0][13] ), .ck(clk), .q(
        m1Inputs[13]) );
  dp_1 \INPUTSRAM/q_reg[12]  ( .ip(\INPUTSRAM/mem_i[0][12] ), .ck(clk), .q(
        m1Inputs[12]) );
  dp_1 \INPUTSRAM/q_reg[108]  ( .ip(\INPUTSRAM/mem_i[6][12] ), .ck(clk), .q(
        m1Inputs[108]) );
  dp_1 \INPUTSRAM/q_reg[151]  ( .ip(\INPUTSRAM/mem_i[9][7] ), .ck(clk), .q(
        m1Inputs[151]) );
  dp_1 \INPUTSRAM/q_reg[148]  ( .ip(\INPUTSRAM/mem_i[9][4] ), .ck(clk), .q(
        m1Inputs[148]) );
  dp_1 \WEIGHT_2/q_reg[4]  ( .ip(n2140), .ck(clk), .q(q_w2[4]) );
  dp_1 \INPUTSRAM/q_reg[121]  ( .ip(\INPUTSRAM/mem_i[7][9] ), .ck(clk), .q(
        m1Inputs[121]) );
  dp_1 \INPUTSRAM/q_reg[122]  ( .ip(\INPUTSRAM/mem_i[7][10] ), .ck(clk), .q(
        m1Inputs[122]) );
  dp_1 \INPUTSRAM/q_reg[152]  ( .ip(\INPUTSRAM/mem_i[9][8] ), .ck(clk), .q(
        m1Inputs[152]) );
  dp_1 \INPUTSRAM/q_reg[58]  ( .ip(\INPUTSRAM/mem_i[3][10] ), .ck(clk), .q(
        m1Inputs[58]) );
  dp_1 \INPUTSRAM/q_reg[135]  ( .ip(\INPUTSRAM/mem_i[8][7] ), .ck(clk), .q(
        m1Inputs[135]) );
  dp_1 \INPUTSRAM/q_reg[149]  ( .ip(\INPUTSRAM/mem_i[9][5] ), .ck(clk), .q(
        m1Inputs[149]) );
  dp_1 \INPUTSRAM/q_reg[76]  ( .ip(\INPUTSRAM/mem_i[4][12] ), .ck(clk), .q(
        m1Inputs[76]) );
  dp_1 \INPUTSRAM/q_reg[107]  ( .ip(\INPUTSRAM/mem_i[6][11] ), .ck(clk), .q(
        m1Inputs[107]) );
  dp_1 \INPUTSRAM/q_reg[77]  ( .ip(\INPUTSRAM/mem_i[4][13] ), .ck(clk), .q(
        m1Inputs[77]) );
  dp_1 \INPUTSRAM/q_reg[132]  ( .ip(\INPUTSRAM/mem_i[8][4] ), .ck(clk), .q(
        m1Inputs[132]) );
  dp_1 \INPUTSRAM/q_reg[59]  ( .ip(\INPUTSRAM/mem_i[3][11] ), .ck(clk), .q(
        m1Inputs[59]) );
  dp_1 \INPUTSRAM/q_reg[20]  ( .ip(\INPUTSRAM/mem_i[1][4] ), .ck(clk), .q(
        m1Inputs[20]) );
  dp_1 \INPUTSRAM/q_reg[57]  ( .ip(\INPUTSRAM/mem_i[3][9] ), .ck(clk), .q(
        m1Inputs[57]) );
  dp_1 \INPUTSRAM/q_reg[9]  ( .ip(\INPUTSRAM/mem_i[0][9] ), .ck(clk), .q(
        m1Inputs[9]) );
  dp_1 \INPUTSRAM/q_reg[136]  ( .ip(\INPUTSRAM/mem_i[8][8] ), .ck(clk), .q(
        m1Inputs[136]) );
  dp_1 \INPUTSRAM/q_reg[92]  ( .ip(\INPUTSRAM/mem_i[5][12] ), .ck(clk), .q(
        m1Inputs[92]) );
  dp_1 \INPUTSRAM/q_reg[93]  ( .ip(\INPUTSRAM/mem_i[5][13] ), .ck(clk), .q(
        m1Inputs[93]) );
  dp_1 \INPUTSRAM/q_reg[21]  ( .ip(\INPUTSRAM/mem_i[1][5] ), .ck(clk), .q(
        m1Inputs[21]) );
  dp_1 \INPUTSRAM/q_reg[105]  ( .ip(\INPUTSRAM/mem_i[6][9] ), .ck(clk), .q(
        m1Inputs[105]) );
  dp_1 \INPUTSRAM/q_reg[60]  ( .ip(\INPUTSRAM/mem_i[3][12] ), .ck(clk), .q(
        m1Inputs[60]) );
  dp_1 \INPUTSRAM/q_reg[61]  ( .ip(\INPUTSRAM/mem_i[3][13] ), .ck(clk), .q(
        m1Inputs[61]) );
  dp_1 \INPUTSRAM/q_reg[106]  ( .ip(\INPUTSRAM/mem_i[6][10] ), .ck(clk), .q(
        m1Inputs[106]) );
  dp_1 \INPUTSRAM/q_reg[103]  ( .ip(\INPUTSRAM/mem_i[6][7] ), .ck(clk), .q(
        m1Inputs[103]) );
  dp_1 \INPUTSRAM/q_reg[89]  ( .ip(\INPUTSRAM/mem_i[5][9] ), .ck(clk), .q(
        m1Inputs[89]) );
  dp_1 \INPUTSRAM/q_reg[104]  ( .ip(\INPUTSRAM/mem_i[6][8] ), .ck(clk), .q(
        m1Inputs[104]) );
  dp_1 \INPUTSRAM/q_reg[114]  ( .ip(\INPUTSRAM/mem_i[7][2] ), .ck(clk), .q(
        m1Inputs[114]) );
  dp_1 \INPUTSRAM/q_reg[73]  ( .ip(\INPUTSRAM/mem_i[4][9] ), .ck(clk), .q(
        m1Inputs[73]) );
  dp_1 \INPUTSRAM/q_reg[10]  ( .ip(\INPUTSRAM/mem_i[0][10] ), .ck(clk), .q(
        m1Inputs[10]) );
  dp_1 \INPUTSRAM/q_reg[11]  ( .ip(\INPUTSRAM/mem_i[0][11] ), .ck(clk), .q(
        m1Inputs[11]) );
  dp_1 \INPUTSRAM/q_reg[35]  ( .ip(\INPUTSRAM/mem_i[2][3] ), .ck(clk), .q(
        m1Inputs[35]) );
  dp_1 \INPUTSRAM/q_reg[38]  ( .ip(\INPUTSRAM/mem_i[2][6] ), .ck(clk), .q(
        m1Inputs[38]) );
  dp_1 \INPUTSRAM/q_reg[71]  ( .ip(\INPUTSRAM/mem_i[4][7] ), .ck(clk), .q(
        m1Inputs[71]) );
  dp_1 \WEIGHT_2/q_reg[1]  ( .ip(n2143), .ck(clk), .q(q_w2[1]) );
  dp_1 \WEIGHT_2/q_reg[3]  ( .ip(n2141), .ck(clk), .q(q_w2[3]) );
  dp_1 \WEIGHT_2/q_reg[0]  ( .ip(n2144), .ck(clk), .q(q_w2[0]) );
  dp_1 \INPUTSRAM/q_reg[46]  ( .ip(\INPUTSRAM/mem_i[2][14] ), .ck(clk), .q(
        m1Inputs[46]) );
  dp_1 \INPUTSRAM/q_reg[72]  ( .ip(\INPUTSRAM/mem_i[4][8] ), .ck(clk), .q(
        m1Inputs[72]) );
  dp_1 \INPUTSRAM/q_reg[90]  ( .ip(\INPUTSRAM/mem_i[5][10] ), .ck(clk), .q(
        m1Inputs[90]) );
  dp_1 \INPUTSRAM/q_reg[116]  ( .ip(\INPUTSRAM/mem_i[7][4] ), .ck(clk), .q(
        m1Inputs[116]) );
  dp_1 \INPUTSRAM/q_reg[66]  ( .ip(\INPUTSRAM/mem_i[4][2] ), .ck(clk), .q(
        m1Inputs[66]) );
  dp_1 \INPUTSRAM/q_reg[91]  ( .ip(\INPUTSRAM/mem_i[5][11] ), .ck(clk), .q(
        m1Inputs[91]) );
  dp_1 \INPUTSRAM/q_reg[119]  ( .ip(\INPUTSRAM/mem_i[7][7] ), .ck(clk), .q(
        m1Inputs[119]) );
  dp_1 \INPUTSRAM/q_reg[74]  ( .ip(\INPUTSRAM/mem_i[4][10] ), .ck(clk), .q(
        m1Inputs[74]) );
  dp_1 \INPUTSRAM/q_reg[117]  ( .ip(\INPUTSRAM/mem_i[7][5] ), .ck(clk), .q(
        m1Inputs[117]) );
  dp_1 \INPUTSRAM/q_reg[120]  ( .ip(\INPUTSRAM/mem_i[7][8] ), .ck(clk), .q(
        m1Inputs[120]) );
  dp_1 \INPUTSRAM/q_reg[75]  ( .ip(\INPUTSRAM/mem_i[4][11] ), .ck(clk), .q(
        m1Inputs[75]) );
  dp_1 \INPUTSRAM/q_reg[2]  ( .ip(\INPUTSRAM/mem_i[0][2] ), .ck(clk), .q(
        m1Inputs[2]) );
  dp_1 \INPUTSRAM/q_reg[98]  ( .ip(\INPUTSRAM/mem_i[6][2] ), .ck(clk), .q(
        m1Inputs[98]) );
  dp_1 \INPUTSRAM/q_reg[50]  ( .ip(\INPUTSRAM/mem_i[3][2] ), .ck(clk), .q(
        m1Inputs[50]) );
  dp_1 \INPUTSRAM/q_reg[45]  ( .ip(\INPUTSRAM/mem_i[2][13] ), .ck(clk), .q(
        m1Inputs[45]) );
  dp_1 \INPUTSRAM/q_reg[44]  ( .ip(\INPUTSRAM/mem_i[2][12] ), .ck(clk), .q(
        m1Inputs[44]) );
  dp_1 \INPUTSRAM/q_reg[68]  ( .ip(\INPUTSRAM/mem_i[4][4] ), .ck(clk), .q(
        m1Inputs[68]) );
  dp_1 \INPUTSRAM/q_reg[41]  ( .ip(\INPUTSRAM/mem_i[2][9] ), .ck(clk), .q(
        m1Inputs[41]) );
  dp_1 \INPUTSRAM/q_reg[69]  ( .ip(\INPUTSRAM/mem_i[4][5] ), .ck(clk), .q(
        m1Inputs[69]) );
  dp_1 \INPUTSRAM/q_reg[82]  ( .ip(\INPUTSRAM/mem_i[5][2] ), .ck(clk), .q(
        m1Inputs[82]) );
  dp_1 \INPUTSRAM/q_reg[4]  ( .ip(\INPUTSRAM/mem_i[0][4] ), .ck(clk), .q(
        m1Inputs[4]) );
  dp_1 \INPUTSRAM/q_reg[7]  ( .ip(\INPUTSRAM/mem_i[0][7] ), .ck(clk), .q(
        m1Inputs[7]) );
  dp_1 \INPUTSRAM/q_reg[8]  ( .ip(\INPUTSRAM/mem_i[0][8] ), .ck(clk), .q(
        m1Inputs[8]) );
  dp_1 \INPUTSRAM/q_reg[5]  ( .ip(\INPUTSRAM/mem_i[0][5] ), .ck(clk), .q(
        m1Inputs[5]) );
  dp_1 \INPUTSRAM/q_reg[52]  ( .ip(\INPUTSRAM/mem_i[3][4] ), .ck(clk), .q(
        m1Inputs[52]) );
  dp_1 \INPUTSRAM/q_reg[53]  ( .ip(\INPUTSRAM/mem_i[3][5] ), .ck(clk), .q(
        m1Inputs[53]) );
  dp_1 \INPUTSRAM/q_reg[55]  ( .ip(\INPUTSRAM/mem_i[3][7] ), .ck(clk), .q(
        m1Inputs[55]) );
  dp_1 \INPUTSRAM/q_reg[100]  ( .ip(\INPUTSRAM/mem_i[6][4] ), .ck(clk), .q(
        m1Inputs[100]) );
  dp_1 \INPUTSRAM/q_reg[56]  ( .ip(\INPUTSRAM/mem_i[3][8] ), .ck(clk), .q(
        m1Inputs[56]) );
  dp_1 \INPUTSRAM/q_reg[42]  ( .ip(\INPUTSRAM/mem_i[2][10] ), .ck(clk), .q(
        m1Inputs[42]) );
  dp_1 \INPUTSRAM/q_reg[84]  ( .ip(\INPUTSRAM/mem_i[5][4] ), .ck(clk), .q(
        m1Inputs[84]) );
  dp_1 \INPUTSRAM/q_reg[43]  ( .ip(\INPUTSRAM/mem_i[2][11] ), .ck(clk), .q(
        m1Inputs[43]) );
  dp_1 \INPUTSRAM/q_reg[87]  ( .ip(\INPUTSRAM/mem_i[5][7] ), .ck(clk), .q(
        m1Inputs[87]) );
  dp_1 \INPUTSRAM/q_reg[85]  ( .ip(\INPUTSRAM/mem_i[5][5] ), .ck(clk), .q(
        m1Inputs[85]) );
  dp_1 \INPUTSRAM/q_reg[88]  ( .ip(\INPUTSRAM/mem_i[5][8] ), .ck(clk), .q(
        m1Inputs[88]) );
  dp_1 \INPUTSRAM/q_reg[34]  ( .ip(\INPUTSRAM/mem_i[2][2] ), .ck(clk), .q(
        m1Inputs[34]) );
  dp_1 \INPUTSRAM/q_reg[36]  ( .ip(\INPUTSRAM/mem_i[2][4] ), .ck(clk), .q(
        m1Inputs[36]) );
  dp_1 \INPUTSRAM/q_reg[39]  ( .ip(\INPUTSRAM/mem_i[2][7] ), .ck(clk), .q(
        m1Inputs[39]) );
  dp_1 \INPUTSRAM/q_reg[40]  ( .ip(\INPUTSRAM/mem_i[2][8] ), .ck(clk), .q(
        m1Inputs[40]) );
  nand2_1 U4336 ( .ip1(w2SramWeOffChip), .ip2(q_w2[10]), .op(n4140) );
  nor2_1 U4337 ( .ip1(\CNTRL/currentState [0]), .ip2(\CNTRL/currentState [1]), 
        .op(n15092) );
  nand2_1 U4338 ( .ip1(n15092), .ip2(\CNTRL/currentState [2]), .op(n15087) );
  inv_1 U4339 ( .ip(n15087), .op(n15624) );
  nand2_1 U4340 ( .ip1(n15624), .ip2(\CNTRL/count_10Q [3]), .op(n4358) );
  nor3_1 U4341 ( .ip1(\CNTRL/count_10Q [0]), .ip2(w2SramWeOffChip), .ip3(n4358), .op(n4337) );
  nand2_1 U4342 ( .ip1(n4337), .ip2(\WEIGHT_2/mem_w2[8][10] ), .op(n4139) );
  inv_1 U4343 ( .ip(\CNTRL/count_10Q [0]), .op(n15132) );
  nor2_1 U4344 ( .ip1(n15087), .ip2(n15132), .op(n4354) );
  inv_1 U4345 ( .ip(w2SramWeOffChip), .op(n4113) );
  and3_1 U4346 ( .ip1(\CNTRL/count_10Q [3]), .ip2(n4354), .ip3(n4113), .op(
        n4338) );
  nand2_1 U4347 ( .ip1(n4338), .ip2(\WEIGHT_2/mem_w2[9][10] ), .op(n4138) );
  and2_1 U4348 ( .ip1(n4358), .ip2(n4113), .op(n4349) );
  mux2_1 U4349 ( .ip1(n4354), .ip2(weight2AddrOffChip[0]), .s(w2SramWeOffChip), 
        .op(n4132) );
  inv_1 U4350 ( .ip(n4132), .op(n4124) );
  nand2_1 U4351 ( .ip1(n15624), .ip2(\CNTRL/count_10Q [1]), .op(n4390) );
  nor2_1 U4352 ( .ip1(w2SramWeOffChip), .ip2(n4390), .op(n4114) );
  or2_1 U4353 ( .ip1(weight2AddrOffChip[1]), .ip2(n4114), .op(n4116) );
  or2_1 U4354 ( .ip1(w2SramWeOffChip), .ip2(n4114), .op(n4115) );
  nand2_1 U4355 ( .ip1(n4116), .ip2(n4115), .op(n4117) );
  inv_1 U4356 ( .ip(\CNTRL/count_10Q [2]), .op(n15136) );
  nor2_1 U4357 ( .ip1(n15087), .ip2(n15136), .op(n4391) );
  mux2_1 U4358 ( .ip1(n4391), .ip2(weight2AddrOffChip[2]), .s(w2SramWeOffChip), 
        .op(n4121) );
  nand2_1 U4359 ( .ip1(n4117), .ip2(n4121), .op(n4119) );
  nor2_1 U4360 ( .ip1(n4124), .ip2(n4119), .op(n15402) );
  nand2_1 U4361 ( .ip1(\WEIGHT_2/mem_w2[5][10] ), .ip2(n15402), .op(n4135) );
  inv_1 U4362 ( .ip(n4121), .op(n4118) );
  inv_1 U4363 ( .ip(n4117), .op(n4120) );
  nand2_1 U4364 ( .ip1(n4118), .ip2(n4120), .op(n4123) );
  nor2_1 U4365 ( .ip1(n4132), .ip2(n4123), .op(n15396) );
  nand2_1 U4366 ( .ip1(n4118), .ip2(n4117), .op(n4131) );
  nor2_1 U4367 ( .ip1(n4131), .ip2(n4124), .op(n15411) );
  and2_1 U4368 ( .ip1(n15411), .ip2(\WEIGHT_2/mem_w2[1][10] ), .op(n4130) );
  nor2_1 U4369 ( .ip1(n4132), .ip2(n4119), .op(n15400) );
  nand2_1 U4370 ( .ip1(n15400), .ip2(\WEIGHT_2/mem_w2[4][10] ), .op(n4128) );
  nand2_1 U4371 ( .ip1(n4121), .ip2(n4120), .op(n4122) );
  nor2_1 U4372 ( .ip1(n4124), .ip2(n4122), .op(n15407) );
  nand2_1 U4373 ( .ip1(n15407), .ip2(\WEIGHT_2/mem_w2[7][10] ), .op(n4127) );
  nor2_1 U4374 ( .ip1(n4132), .ip2(n4122), .op(n15404) );
  nand2_1 U4375 ( .ip1(n15404), .ip2(\WEIGHT_2/mem_w2[6][10] ), .op(n4126) );
  nor2_1 U4376 ( .ip1(n4124), .ip2(n4123), .op(n15398) );
  nand2_1 U4377 ( .ip1(n15398), .ip2(\WEIGHT_2/mem_w2[3][10] ), .op(n4125) );
  nand4_1 U4378 ( .ip1(n4128), .ip2(n4127), .ip3(n4126), .ip4(n4125), .op(
        n4129) );
  not_ab_or_c_or_d U4379 ( .ip1(\WEIGHT_2/mem_w2[2][10] ), .ip2(n15396), .ip3(
        n4130), .ip4(n4129), .op(n4134) );
  nor2_1 U4380 ( .ip1(n4132), .ip2(n4131), .op(n15409) );
  nand2_1 U4381 ( .ip1(n15409), .ip2(\WEIGHT_2/mem_w2[0][10] ), .op(n4133) );
  nand3_1 U4382 ( .ip1(n4135), .ip2(n4134), .ip3(n4133), .op(n4136) );
  nand2_1 U4383 ( .ip1(n4349), .ip2(n4136), .op(n4137) );
  nand4_1 U4384 ( .ip1(n4140), .ip2(n4139), .ip3(n4138), .ip4(n4137), .op(
        n2134) );
  nand2_1 U4385 ( .ip1(n4337), .ip2(\WEIGHT_2/mem_w2[8][14] ), .op(n4154) );
  nand2_1 U4386 ( .ip1(w2SramWeOffChip), .ip2(q_w2[14]), .op(n4153) );
  nand2_1 U4387 ( .ip1(n4338), .ip2(\WEIGHT_2/mem_w2[9][14] ), .op(n4152) );
  nand2_1 U4388 ( .ip1(\WEIGHT_2/mem_w2[0][14] ), .ip2(n15409), .op(n4149) );
  and2_1 U4389 ( .ip1(n15411), .ip2(\WEIGHT_2/mem_w2[1][14] ), .op(n4146) );
  nand2_1 U4390 ( .ip1(n15400), .ip2(\WEIGHT_2/mem_w2[4][14] ), .op(n4144) );
  nand2_1 U4391 ( .ip1(n15407), .ip2(\WEIGHT_2/mem_w2[7][14] ), .op(n4143) );
  nand2_1 U4392 ( .ip1(n15396), .ip2(\WEIGHT_2/mem_w2[2][14] ), .op(n4142) );
  nand2_1 U4393 ( .ip1(n15404), .ip2(\WEIGHT_2/mem_w2[6][14] ), .op(n4141) );
  nand4_1 U4394 ( .ip1(n4144), .ip2(n4143), .ip3(n4142), .ip4(n4141), .op(
        n4145) );
  not_ab_or_c_or_d U4395 ( .ip1(\WEIGHT_2/mem_w2[5][14] ), .ip2(n15402), .ip3(
        n4146), .ip4(n4145), .op(n4148) );
  nand2_1 U4396 ( .ip1(n15398), .ip2(\WEIGHT_2/mem_w2[3][14] ), .op(n4147) );
  nand3_1 U4397 ( .ip1(n4149), .ip2(n4148), .ip3(n4147), .op(n4150) );
  nand2_1 U4398 ( .ip1(n4349), .ip2(n4150), .op(n4151) );
  nand4_1 U4399 ( .ip1(n4154), .ip2(n4153), .ip3(n4152), .ip4(n4151), .op(
        n2130) );
  nand2_1 U4400 ( .ip1(w2SramWeOffChip), .ip2(q_w2[15]), .op(n4168) );
  nand2_1 U4401 ( .ip1(n4337), .ip2(\WEIGHT_2/mem_w2[8][15] ), .op(n4167) );
  nand2_1 U4402 ( .ip1(n4338), .ip2(\WEIGHT_2/mem_w2[9][15] ), .op(n4166) );
  nand2_1 U4403 ( .ip1(\WEIGHT_2/mem_w2[0][15] ), .ip2(n15409), .op(n4163) );
  and2_1 U4404 ( .ip1(n15411), .ip2(\WEIGHT_2/mem_w2[1][15] ), .op(n4160) );
  nand2_1 U4405 ( .ip1(n15400), .ip2(\WEIGHT_2/mem_w2[4][15] ), .op(n4158) );
  nand2_1 U4406 ( .ip1(n15407), .ip2(\WEIGHT_2/mem_w2[7][15] ), .op(n4157) );
  nand2_1 U4407 ( .ip1(n15396), .ip2(\WEIGHT_2/mem_w2[2][15] ), .op(n4156) );
  nand2_1 U4408 ( .ip1(n15402), .ip2(\WEIGHT_2/mem_w2[5][15] ), .op(n4155) );
  nand4_1 U4409 ( .ip1(n4158), .ip2(n4157), .ip3(n4156), .ip4(n4155), .op(
        n4159) );
  not_ab_or_c_or_d U4410 ( .ip1(\WEIGHT_2/mem_w2[3][15] ), .ip2(n15398), .ip3(
        n4160), .ip4(n4159), .op(n4162) );
  nand2_1 U4411 ( .ip1(n15404), .ip2(\WEIGHT_2/mem_w2[6][15] ), .op(n4161) );
  nand3_1 U4412 ( .ip1(n4163), .ip2(n4162), .ip3(n4161), .op(n4164) );
  nand2_1 U4413 ( .ip1(n4349), .ip2(n4164), .op(n4165) );
  nand4_1 U4414 ( .ip1(n4168), .ip2(n4167), .ip3(n4166), .ip4(n4165), .op(
        n2129) );
  nand2_1 U4415 ( .ip1(w2SramWeOffChip), .ip2(q_w2[12]), .op(n4182) );
  nand2_1 U4416 ( .ip1(n4337), .ip2(\WEIGHT_2/mem_w2[8][12] ), .op(n4181) );
  nand2_1 U4417 ( .ip1(n4338), .ip2(\WEIGHT_2/mem_w2[9][12] ), .op(n4180) );
  nand2_1 U4418 ( .ip1(\WEIGHT_2/mem_w2[0][12] ), .ip2(n15409), .op(n4177) );
  and2_1 U4419 ( .ip1(n15411), .ip2(\WEIGHT_2/mem_w2[1][12] ), .op(n4174) );
  nand2_1 U4420 ( .ip1(n15402), .ip2(\WEIGHT_2/mem_w2[5][12] ), .op(n4172) );
  nand2_1 U4421 ( .ip1(n15396), .ip2(\WEIGHT_2/mem_w2[2][12] ), .op(n4171) );
  nand2_1 U4422 ( .ip1(n15400), .ip2(\WEIGHT_2/mem_w2[4][12] ), .op(n4170) );
  nand2_1 U4423 ( .ip1(n15407), .ip2(\WEIGHT_2/mem_w2[7][12] ), .op(n4169) );
  nand4_1 U4424 ( .ip1(n4172), .ip2(n4171), .ip3(n4170), .ip4(n4169), .op(
        n4173) );
  not_ab_or_c_or_d U4425 ( .ip1(n15404), .ip2(\WEIGHT_2/mem_w2[6][12] ), .ip3(
        n4174), .ip4(n4173), .op(n4176) );
  nand2_1 U4426 ( .ip1(n15398), .ip2(\WEIGHT_2/mem_w2[3][12] ), .op(n4175) );
  nand3_1 U4427 ( .ip1(n4177), .ip2(n4176), .ip3(n4175), .op(n4178) );
  nand2_1 U4428 ( .ip1(n4349), .ip2(n4178), .op(n4179) );
  nand4_1 U4429 ( .ip1(n4182), .ip2(n4181), .ip3(n4180), .ip4(n4179), .op(
        n2132) );
  nand2_1 U4430 ( .ip1(n4337), .ip2(\WEIGHT_2/mem_w2[8][6] ), .op(n4196) );
  nand2_1 U4431 ( .ip1(w2SramWeOffChip), .ip2(q_w2[6]), .op(n4195) );
  nand2_1 U4432 ( .ip1(n4338), .ip2(\WEIGHT_2/mem_w2[9][6] ), .op(n4194) );
  nand2_1 U4433 ( .ip1(\WEIGHT_2/mem_w2[5][6] ), .ip2(n15402), .op(n4191) );
  and2_1 U4434 ( .ip1(n15411), .ip2(\WEIGHT_2/mem_w2[1][6] ), .op(n4188) );
  nand2_1 U4435 ( .ip1(n15398), .ip2(\WEIGHT_2/mem_w2[3][6] ), .op(n4186) );
  nand2_1 U4436 ( .ip1(n15400), .ip2(\WEIGHT_2/mem_w2[4][6] ), .op(n4185) );
  nand2_1 U4437 ( .ip1(n15396), .ip2(\WEIGHT_2/mem_w2[2][6] ), .op(n4184) );
  nand2_1 U4438 ( .ip1(n15404), .ip2(\WEIGHT_2/mem_w2[6][6] ), .op(n4183) );
  nand4_1 U4439 ( .ip1(n4186), .ip2(n4185), .ip3(n4184), .ip4(n4183), .op(
        n4187) );
  not_ab_or_c_or_d U4440 ( .ip1(n15407), .ip2(\WEIGHT_2/mem_w2[7][6] ), .ip3(
        n4188), .ip4(n4187), .op(n4190) );
  nand2_1 U4441 ( .ip1(n15409), .ip2(\WEIGHT_2/mem_w2[0][6] ), .op(n4189) );
  nand3_1 U4442 ( .ip1(n4191), .ip2(n4190), .ip3(n4189), .op(n4192) );
  nand2_1 U4443 ( .ip1(n4349), .ip2(n4192), .op(n4193) );
  nand4_1 U4444 ( .ip1(n4196), .ip2(n4195), .ip3(n4194), .ip4(n4193), .op(
        n2138) );
  nand2_1 U4445 ( .ip1(w2SramWeOffChip), .ip2(q_w2[11]), .op(n4210) );
  nand2_1 U4446 ( .ip1(n4337), .ip2(\WEIGHT_2/mem_w2[8][11] ), .op(n4209) );
  nand2_1 U4447 ( .ip1(n4338), .ip2(\WEIGHT_2/mem_w2[9][11] ), .op(n4208) );
  nand2_1 U4448 ( .ip1(\WEIGHT_2/mem_w2[0][11] ), .ip2(n15409), .op(n4205) );
  and2_1 U4449 ( .ip1(n15411), .ip2(\WEIGHT_2/mem_w2[1][11] ), .op(n4202) );
  nand2_1 U4450 ( .ip1(n15400), .ip2(\WEIGHT_2/mem_w2[4][11] ), .op(n4200) );
  nand2_1 U4451 ( .ip1(n15402), .ip2(\WEIGHT_2/mem_w2[5][11] ), .op(n4199) );
  nand2_1 U4452 ( .ip1(n15396), .ip2(\WEIGHT_2/mem_w2[2][11] ), .op(n4198) );
  nand2_1 U4453 ( .ip1(n15404), .ip2(\WEIGHT_2/mem_w2[6][11] ), .op(n4197) );
  nand4_1 U4454 ( .ip1(n4200), .ip2(n4199), .ip3(n4198), .ip4(n4197), .op(
        n4201) );
  not_ab_or_c_or_d U4455 ( .ip1(n15407), .ip2(\WEIGHT_2/mem_w2[7][11] ), .ip3(
        n4202), .ip4(n4201), .op(n4204) );
  nand2_1 U4456 ( .ip1(n15398), .ip2(\WEIGHT_2/mem_w2[3][11] ), .op(n4203) );
  nand3_1 U4457 ( .ip1(n4205), .ip2(n4204), .ip3(n4203), .op(n4206) );
  nand2_1 U4458 ( .ip1(n4349), .ip2(n4206), .op(n4207) );
  nand4_1 U4459 ( .ip1(n4210), .ip2(n4209), .ip3(n4208), .ip4(n4207), .op(
        n2133) );
  nand2_1 U4460 ( .ip1(q_w2[2]), .ip2(w2SramWeOffChip), .op(n4224) );
  nand2_1 U4461 ( .ip1(n4337), .ip2(\WEIGHT_2/mem_w2[8][2] ), .op(n4223) );
  nand2_1 U4462 ( .ip1(n4338), .ip2(\WEIGHT_2/mem_w2[9][2] ), .op(n4222) );
  nand2_1 U4463 ( .ip1(n15396), .ip2(\WEIGHT_2/mem_w2[2][2] ), .op(n4219) );
  and2_1 U4464 ( .ip1(n15411), .ip2(\WEIGHT_2/mem_w2[1][2] ), .op(n4216) );
  nand2_1 U4465 ( .ip1(n15398), .ip2(\WEIGHT_2/mem_w2[3][2] ), .op(n4214) );
  nand2_1 U4466 ( .ip1(n15400), .ip2(\WEIGHT_2/mem_w2[4][2] ), .op(n4213) );
  nand2_1 U4467 ( .ip1(n15402), .ip2(\WEIGHT_2/mem_w2[5][2] ), .op(n4212) );
  nand2_1 U4468 ( .ip1(n15407), .ip2(\WEIGHT_2/mem_w2[7][2] ), .op(n4211) );
  nand4_1 U4469 ( .ip1(n4214), .ip2(n4213), .ip3(n4212), .ip4(n4211), .op(
        n4215) );
  not_ab_or_c_or_d U4470 ( .ip1(n15409), .ip2(\WEIGHT_2/mem_w2[0][2] ), .ip3(
        n4216), .ip4(n4215), .op(n4218) );
  nand2_1 U4471 ( .ip1(n15404), .ip2(\WEIGHT_2/mem_w2[6][2] ), .op(n4217) );
  nand3_1 U4472 ( .ip1(n4219), .ip2(n4218), .ip3(n4217), .op(n4220) );
  nand2_1 U4473 ( .ip1(n4349), .ip2(n4220), .op(n4221) );
  nand4_1 U4474 ( .ip1(n4224), .ip2(n4223), .ip3(n4222), .ip4(n4221), .op(
        n2142) );
  nand2_1 U4475 ( .ip1(q_w2[1]), .ip2(w2SramWeOffChip), .op(n4238) );
  nand2_1 U4476 ( .ip1(n4337), .ip2(\WEIGHT_2/mem_w2[8][1] ), .op(n4237) );
  nand2_1 U4477 ( .ip1(n4338), .ip2(\WEIGHT_2/mem_w2[9][1] ), .op(n4236) );
  nand2_1 U4478 ( .ip1(\WEIGHT_2/mem_w2[4][1] ), .ip2(n15400), .op(n4233) );
  and2_1 U4479 ( .ip1(n15411), .ip2(\WEIGHT_2/mem_w2[1][1] ), .op(n4230) );
  nand2_1 U4480 ( .ip1(n15402), .ip2(\WEIGHT_2/mem_w2[5][1] ), .op(n4228) );
  nand2_1 U4481 ( .ip1(n15404), .ip2(\WEIGHT_2/mem_w2[6][1] ), .op(n4227) );
  nand2_1 U4482 ( .ip1(n15409), .ip2(\WEIGHT_2/mem_w2[0][1] ), .op(n4226) );
  nand2_1 U4483 ( .ip1(n15407), .ip2(\WEIGHT_2/mem_w2[7][1] ), .op(n4225) );
  nand4_1 U4484 ( .ip1(n4228), .ip2(n4227), .ip3(n4226), .ip4(n4225), .op(
        n4229) );
  not_ab_or_c_or_d U4485 ( .ip1(\WEIGHT_2/mem_w2[2][1] ), .ip2(n15396), .ip3(
        n4230), .ip4(n4229), .op(n4232) );
  nand2_1 U4486 ( .ip1(n15398), .ip2(\WEIGHT_2/mem_w2[3][1] ), .op(n4231) );
  nand3_1 U4487 ( .ip1(n4233), .ip2(n4232), .ip3(n4231), .op(n4234) );
  nand2_1 U4488 ( .ip1(n4349), .ip2(n4234), .op(n4235) );
  nand4_1 U4489 ( .ip1(n4238), .ip2(n4237), .ip3(n4236), .ip4(n4235), .op(
        n2143) );
  nand2_1 U4490 ( .ip1(w2SramWeOffChip), .ip2(q_w2[5]), .op(n4252) );
  nand2_1 U4491 ( .ip1(n4337), .ip2(\WEIGHT_2/mem_w2[8][5] ), .op(n4251) );
  nand2_1 U4492 ( .ip1(n4338), .ip2(\WEIGHT_2/mem_w2[9][5] ), .op(n4250) );
  nand2_1 U4493 ( .ip1(n15396), .ip2(\WEIGHT_2/mem_w2[2][5] ), .op(n4247) );
  and2_1 U4494 ( .ip1(n15411), .ip2(\WEIGHT_2/mem_w2[1][5] ), .op(n4244) );
  nand2_1 U4495 ( .ip1(n15400), .ip2(\WEIGHT_2/mem_w2[4][5] ), .op(n4242) );
  nand2_1 U4496 ( .ip1(n15409), .ip2(\WEIGHT_2/mem_w2[0][5] ), .op(n4241) );
  nand2_1 U4497 ( .ip1(n15402), .ip2(\WEIGHT_2/mem_w2[5][5] ), .op(n4240) );
  nand2_1 U4498 ( .ip1(n15398), .ip2(\WEIGHT_2/mem_w2[3][5] ), .op(n4239) );
  nand4_1 U4499 ( .ip1(n4242), .ip2(n4241), .ip3(n4240), .ip4(n4239), .op(
        n4243) );
  not_ab_or_c_or_d U4500 ( .ip1(\WEIGHT_2/mem_w2[7][5] ), .ip2(n15407), .ip3(
        n4244), .ip4(n4243), .op(n4246) );
  nand2_1 U4501 ( .ip1(n15404), .ip2(\WEIGHT_2/mem_w2[6][5] ), .op(n4245) );
  nand3_1 U4502 ( .ip1(n4247), .ip2(n4246), .ip3(n4245), .op(n4248) );
  nand2_1 U4503 ( .ip1(n4349), .ip2(n4248), .op(n4249) );
  nand4_1 U4504 ( .ip1(n4252), .ip2(n4251), .ip3(n4250), .ip4(n4249), .op(
        n2139) );
  nand2_1 U4505 ( .ip1(n4337), .ip2(\WEIGHT_2/mem_w2[8][0] ), .op(n4266) );
  nand2_1 U4506 ( .ip1(q_w2[0]), .ip2(w2SramWeOffChip), .op(n4265) );
  nand2_1 U4507 ( .ip1(n4338), .ip2(\WEIGHT_2/mem_w2[9][0] ), .op(n4264) );
  nand2_1 U4508 ( .ip1(n15402), .ip2(\WEIGHT_2/mem_w2[5][0] ), .op(n4261) );
  and2_1 U4509 ( .ip1(n15411), .ip2(\WEIGHT_2/mem_w2[1][0] ), .op(n4258) );
  nand2_1 U4510 ( .ip1(n15409), .ip2(\WEIGHT_2/mem_w2[0][0] ), .op(n4256) );
  nand2_1 U4511 ( .ip1(n15404), .ip2(\WEIGHT_2/mem_w2[6][0] ), .op(n4255) );
  nand2_1 U4512 ( .ip1(n15407), .ip2(\WEIGHT_2/mem_w2[7][0] ), .op(n4254) );
  nand2_1 U4513 ( .ip1(n15398), .ip2(\WEIGHT_2/mem_w2[3][0] ), .op(n4253) );
  nand4_1 U4514 ( .ip1(n4256), .ip2(n4255), .ip3(n4254), .ip4(n4253), .op(
        n4257) );
  not_ab_or_c_or_d U4515 ( .ip1(n15400), .ip2(\WEIGHT_2/mem_w2[4][0] ), .ip3(
        n4258), .ip4(n4257), .op(n4260) );
  nand2_1 U4516 ( .ip1(n15396), .ip2(\WEIGHT_2/mem_w2[2][0] ), .op(n4259) );
  nand3_1 U4517 ( .ip1(n4261), .ip2(n4260), .ip3(n4259), .op(n4262) );
  nand2_1 U4518 ( .ip1(n4349), .ip2(n4262), .op(n4263) );
  nand4_1 U4519 ( .ip1(n4266), .ip2(n4265), .ip3(n4264), .ip4(n4263), .op(
        n2144) );
  nand2_1 U4520 ( .ip1(w2SramWeOffChip), .ip2(q_w2[9]), .op(n4280) );
  nand2_1 U4521 ( .ip1(n4337), .ip2(\WEIGHT_2/mem_w2[8][9] ), .op(n4279) );
  nand2_1 U4522 ( .ip1(n4338), .ip2(\WEIGHT_2/mem_w2[9][9] ), .op(n4278) );
  nand2_1 U4523 ( .ip1(n15402), .ip2(\WEIGHT_2/mem_w2[5][9] ), .op(n4275) );
  and2_1 U4524 ( .ip1(n15411), .ip2(\WEIGHT_2/mem_w2[1][9] ), .op(n4272) );
  nand2_1 U4525 ( .ip1(n15404), .ip2(\WEIGHT_2/mem_w2[6][9] ), .op(n4270) );
  nand2_1 U4526 ( .ip1(n15396), .ip2(\WEIGHT_2/mem_w2[2][9] ), .op(n4269) );
  nand2_1 U4527 ( .ip1(n15398), .ip2(\WEIGHT_2/mem_w2[3][9] ), .op(n4268) );
  nand2_1 U4528 ( .ip1(n15409), .ip2(\WEIGHT_2/mem_w2[0][9] ), .op(n4267) );
  nand4_1 U4529 ( .ip1(n4270), .ip2(n4269), .ip3(n4268), .ip4(n4267), .op(
        n4271) );
  not_ab_or_c_or_d U4530 ( .ip1(\WEIGHT_2/mem_w2[7][9] ), .ip2(n15407), .ip3(
        n4272), .ip4(n4271), .op(n4274) );
  nand2_1 U4531 ( .ip1(n15400), .ip2(\WEIGHT_2/mem_w2[4][9] ), .op(n4273) );
  nand3_1 U4532 ( .ip1(n4275), .ip2(n4274), .ip3(n4273), .op(n4276) );
  nand2_1 U4533 ( .ip1(n4349), .ip2(n4276), .op(n4277) );
  nand4_1 U4534 ( .ip1(n4280), .ip2(n4279), .ip3(n4278), .ip4(n4277), .op(
        n2135) );
  nand2_1 U4535 ( .ip1(w2SramWeOffChip), .ip2(q_w2[7]), .op(n4294) );
  nand2_1 U4536 ( .ip1(n4337), .ip2(\WEIGHT_2/mem_w2[8][7] ), .op(n4293) );
  nand2_1 U4537 ( .ip1(n4338), .ip2(\WEIGHT_2/mem_w2[9][7] ), .op(n4292) );
  nand2_1 U4538 ( .ip1(n15402), .ip2(\WEIGHT_2/mem_w2[5][7] ), .op(n4289) );
  and2_1 U4539 ( .ip1(n15411), .ip2(\WEIGHT_2/mem_w2[1][7] ), .op(n4286) );
  nand2_1 U4540 ( .ip1(n15409), .ip2(\WEIGHT_2/mem_w2[0][7] ), .op(n4284) );
  nand2_1 U4541 ( .ip1(n15398), .ip2(\WEIGHT_2/mem_w2[3][7] ), .op(n4283) );
  nand2_1 U4542 ( .ip1(n15400), .ip2(\WEIGHT_2/mem_w2[4][7] ), .op(n4282) );
  nand2_1 U4543 ( .ip1(n15396), .ip2(\WEIGHT_2/mem_w2[2][7] ), .op(n4281) );
  nand4_1 U4544 ( .ip1(n4284), .ip2(n4283), .ip3(n4282), .ip4(n4281), .op(
        n4285) );
  not_ab_or_c_or_d U4545 ( .ip1(n15404), .ip2(\WEIGHT_2/mem_w2[6][7] ), .ip3(
        n4286), .ip4(n4285), .op(n4288) );
  nand2_1 U4546 ( .ip1(n15407), .ip2(\WEIGHT_2/mem_w2[7][7] ), .op(n4287) );
  nand3_1 U4547 ( .ip1(n4289), .ip2(n4288), .ip3(n4287), .op(n4290) );
  nand2_1 U4548 ( .ip1(n4349), .ip2(n4290), .op(n4291) );
  nand4_1 U4549 ( .ip1(n4294), .ip2(n4293), .ip3(n4292), .ip4(n4291), .op(
        n2137) );
  nand2_1 U4550 ( .ip1(n4337), .ip2(\WEIGHT_2/mem_w2[8][8] ), .op(n4308) );
  nand2_1 U4551 ( .ip1(w2SramWeOffChip), .ip2(q_w2[8]), .op(n4307) );
  nand2_1 U4552 ( .ip1(n4338), .ip2(\WEIGHT_2/mem_w2[9][8] ), .op(n4306) );
  nand2_1 U4553 ( .ip1(n15404), .ip2(\WEIGHT_2/mem_w2[6][8] ), .op(n4303) );
  and2_1 U4554 ( .ip1(n15411), .ip2(\WEIGHT_2/mem_w2[1][8] ), .op(n4300) );
  nand2_1 U4555 ( .ip1(n15407), .ip2(\WEIGHT_2/mem_w2[7][8] ), .op(n4298) );
  nand2_1 U4556 ( .ip1(n15400), .ip2(\WEIGHT_2/mem_w2[4][8] ), .op(n4297) );
  nand2_1 U4557 ( .ip1(n15409), .ip2(\WEIGHT_2/mem_w2[0][8] ), .op(n4296) );
  nand2_1 U4558 ( .ip1(n15396), .ip2(\WEIGHT_2/mem_w2[2][8] ), .op(n4295) );
  nand4_1 U4559 ( .ip1(n4298), .ip2(n4297), .ip3(n4296), .ip4(n4295), .op(
        n4299) );
  not_ab_or_c_or_d U4560 ( .ip1(n15402), .ip2(\WEIGHT_2/mem_w2[5][8] ), .ip3(
        n4300), .ip4(n4299), .op(n4302) );
  nand2_1 U4561 ( .ip1(n15398), .ip2(\WEIGHT_2/mem_w2[3][8] ), .op(n4301) );
  nand3_1 U4562 ( .ip1(n4303), .ip2(n4302), .ip3(n4301), .op(n4304) );
  nand2_1 U4563 ( .ip1(n4349), .ip2(n4304), .op(n4305) );
  nand4_1 U4564 ( .ip1(n4308), .ip2(n4307), .ip3(n4306), .ip4(n4305), .op(
        n2136) );
  nand2_1 U4565 ( .ip1(w2SramWeOffChip), .ip2(q_w2[4]), .op(n4322) );
  nand2_1 U4566 ( .ip1(n4337), .ip2(\WEIGHT_2/mem_w2[8][4] ), .op(n4321) );
  nand2_1 U4567 ( .ip1(n4338), .ip2(\WEIGHT_2/mem_w2[9][4] ), .op(n4320) );
  nand2_1 U4568 ( .ip1(\WEIGHT_2/mem_w2[6][4] ), .ip2(n15404), .op(n4317) );
  and2_1 U4569 ( .ip1(n15411), .ip2(\WEIGHT_2/mem_w2[1][4] ), .op(n4314) );
  nand2_1 U4570 ( .ip1(n15396), .ip2(\WEIGHT_2/mem_w2[2][4] ), .op(n4312) );
  nand2_1 U4571 ( .ip1(n15398), .ip2(\WEIGHT_2/mem_w2[3][4] ), .op(n4311) );
  nand2_1 U4572 ( .ip1(n15409), .ip2(\WEIGHT_2/mem_w2[0][4] ), .op(n4310) );
  nand2_1 U4573 ( .ip1(n15400), .ip2(\WEIGHT_2/mem_w2[4][4] ), .op(n4309) );
  nand4_1 U4574 ( .ip1(n4312), .ip2(n4311), .ip3(n4310), .ip4(n4309), .op(
        n4313) );
  not_ab_or_c_or_d U4575 ( .ip1(n15402), .ip2(\WEIGHT_2/mem_w2[5][4] ), .ip3(
        n4314), .ip4(n4313), .op(n4316) );
  nand2_1 U4576 ( .ip1(n15407), .ip2(\WEIGHT_2/mem_w2[7][4] ), .op(n4315) );
  nand3_1 U4577 ( .ip1(n4317), .ip2(n4316), .ip3(n4315), .op(n4318) );
  nand2_1 U4578 ( .ip1(n4349), .ip2(n4318), .op(n4319) );
  nand4_1 U4579 ( .ip1(n4322), .ip2(n4321), .ip3(n4320), .ip4(n4319), .op(
        n2140) );
  nand2_1 U4580 ( .ip1(n4337), .ip2(\WEIGHT_2/mem_w2[8][13] ), .op(n4336) );
  nand2_1 U4581 ( .ip1(w2SramWeOffChip), .ip2(q_w2[13]), .op(n4335) );
  nand2_1 U4582 ( .ip1(n4338), .ip2(\WEIGHT_2/mem_w2[9][13] ), .op(n4334) );
  nand2_1 U4583 ( .ip1(\WEIGHT_2/mem_w2[6][13] ), .ip2(n15404), .op(n4331) );
  and2_1 U4584 ( .ip1(n15411), .ip2(\WEIGHT_2/mem_w2[1][13] ), .op(n4328) );
  nand2_1 U4585 ( .ip1(n15402), .ip2(\WEIGHT_2/mem_w2[5][13] ), .op(n4326) );
  nand2_1 U4586 ( .ip1(n15409), .ip2(\WEIGHT_2/mem_w2[0][13] ), .op(n4325) );
  nand2_1 U4587 ( .ip1(n15396), .ip2(\WEIGHT_2/mem_w2[2][13] ), .op(n4324) );
  nand2_1 U4588 ( .ip1(n15400), .ip2(\WEIGHT_2/mem_w2[4][13] ), .op(n4323) );
  nand4_1 U4589 ( .ip1(n4326), .ip2(n4325), .ip3(n4324), .ip4(n4323), .op(
        n4327) );
  not_ab_or_c_or_d U4590 ( .ip1(n15407), .ip2(\WEIGHT_2/mem_w2[7][13] ), .ip3(
        n4328), .ip4(n4327), .op(n4330) );
  nand2_1 U4591 ( .ip1(n15398), .ip2(\WEIGHT_2/mem_w2[3][13] ), .op(n4329) );
  nand3_1 U4592 ( .ip1(n4331), .ip2(n4330), .ip3(n4329), .op(n4332) );
  nand2_1 U4593 ( .ip1(n4349), .ip2(n4332), .op(n4333) );
  nand4_1 U4594 ( .ip1(n4336), .ip2(n4335), .ip3(n4334), .ip4(n4333), .op(
        n2131) );
  nand2_1 U4595 ( .ip1(q_w2[3]), .ip2(w2SramWeOffChip), .op(n4353) );
  nand2_1 U4596 ( .ip1(n4337), .ip2(\WEIGHT_2/mem_w2[8][3] ), .op(n4352) );
  nand2_1 U4597 ( .ip1(n4338), .ip2(\WEIGHT_2/mem_w2[9][3] ), .op(n4351) );
  nand2_1 U4598 ( .ip1(n15404), .ip2(\WEIGHT_2/mem_w2[6][3] ), .op(n4347) );
  and2_1 U4599 ( .ip1(n15411), .ip2(\WEIGHT_2/mem_w2[1][3] ), .op(n4344) );
  nand2_1 U4600 ( .ip1(n15402), .ip2(\WEIGHT_2/mem_w2[5][3] ), .op(n4342) );
  nand2_1 U4601 ( .ip1(n15398), .ip2(\WEIGHT_2/mem_w2[3][3] ), .op(n4341) );
  nand2_1 U4602 ( .ip1(n15396), .ip2(\WEIGHT_2/mem_w2[2][3] ), .op(n4340) );
  nand2_1 U4603 ( .ip1(n15409), .ip2(\WEIGHT_2/mem_w2[0][3] ), .op(n4339) );
  nand4_1 U4604 ( .ip1(n4342), .ip2(n4341), .ip3(n4340), .ip4(n4339), .op(
        n4343) );
  not_ab_or_c_or_d U4605 ( .ip1(n15400), .ip2(\WEIGHT_2/mem_w2[4][3] ), .ip3(
        n4344), .ip4(n4343), .op(n4346) );
  nand2_1 U4606 ( .ip1(n15407), .ip2(\WEIGHT_2/mem_w2[7][3] ), .op(n4345) );
  nand3_1 U4607 ( .ip1(n4347), .ip2(n4346), .ip3(n4345), .op(n4348) );
  nand2_1 U4608 ( .ip1(n4349), .ip2(n4348), .op(n4350) );
  nand4_1 U4609 ( .ip1(n4353), .ip2(n4352), .ip3(n4351), .ip4(n4350), .op(
        n2141) );
  or2_1 U4610 ( .ip1(\CNTRL/count_10_2Q [0]), .ip2(n4354), .op(n4356) );
  inv_1 U4611 ( .ip(\CNTRL/currentState [2]), .op(n15083) );
  nor2_1 U4612 ( .ip1(n15092), .ip2(n15083), .op(n15085) );
  or2_1 U4613 ( .ip1(n15085), .ip2(n4354), .op(n4355) );
  nand2_1 U4614 ( .ip1(n4356), .ip2(n4355), .op(n4466) );
  nand2_1 U4615 ( .ip1(n15085), .ip2(\CNTRL/count_10_2Q [3]), .op(n4357) );
  and2_1 U4616 ( .ip1(n4358), .ip2(n4357), .op(n18888) );
  nor2_1 U4617 ( .ip1(n4466), .ip2(n18888), .op(n18899) );
  inv_1 U4618 ( .ip(\CNTRL/count_20Q [1]), .op(n15186) );
  nor2_1 U4619 ( .ip1(n15087), .ip2(n15186), .op(n4359) );
  or2_1 U4620 ( .ip1(\CNTRL/count_10Q [0]), .ip2(n4359), .op(n4361) );
  or2_1 U4621 ( .ip1(n15085), .ip2(n4359), .op(n4360) );
  nand2_1 U4622 ( .ip1(n4361), .ip2(n4360), .op(n4362) );
  inv_1 U4623 ( .ip(n4362), .op(n17610) );
  inv_1 U4624 ( .ip(n4362), .op(n17401) );
  buf_1 U4625 ( .ip(n17401), .op(n15643) );
  mux2_1 U4626 ( .ip1(\ANSWER/mem[0][9][1] ), .ip2(\ANSWER/mem[1][9][1] ), .s(
        n15643), .op(n4368) );
  mux2_1 U4627 ( .ip1(\ANSWER/mem[2][9][1] ), .ip2(\ANSWER/mem[3][9][1] ), .s(
        n15643), .op(n4367) );
  inv_1 U4628 ( .ip(\CNTRL/count_20Q [2]), .op(n15110) );
  nor2_1 U4629 ( .ip1(n15087), .ip2(n15110), .op(n4363) );
  or2_1 U4630 ( .ip1(\CNTRL/count_10Q [1]), .ip2(n4363), .op(n4365) );
  or2_1 U4631 ( .ip1(n15085), .ip2(n4363), .op(n4364) );
  nand2_1 U4632 ( .ip1(n4365), .ip2(n4364), .op(n4366) );
  inv_1 U4633 ( .ip(n4366), .op(n18901) );
  inv_1 U4634 ( .ip(n4366), .op(n15636) );
  mux2_1 U4635 ( .ip1(n4368), .ip2(n4367), .s(n15636), .op(n4375) );
  mux2_1 U4636 ( .ip1(\ANSWER/mem[4][9][1] ), .ip2(\ANSWER/mem[5][9][1] ), .s(
        n15643), .op(n4370) );
  mux2_1 U4637 ( .ip1(\ANSWER/mem[6][9][1] ), .ip2(\ANSWER/mem[7][9][1] ), .s(
        n15643), .op(n4369) );
  mux2_1 U4638 ( .ip1(n4370), .ip2(n4369), .s(n15636), .op(n4374) );
  inv_1 U4639 ( .ip(\CNTRL/count_20Q [3]), .op(n15174) );
  nor2_1 U4640 ( .ip1(n15087), .ip2(n15174), .op(n4371) );
  or2_1 U4641 ( .ip1(\CNTRL/count_10Q [2]), .ip2(n4371), .op(n4373) );
  or2_1 U4642 ( .ip1(n15085), .ip2(n4371), .op(n4372) );
  nand2_1 U4643 ( .ip1(n4373), .ip2(n4372), .op(n17488) );
  inv_1 U4644 ( .ip(n17488), .op(n18878) );
  buf_1 U4645 ( .ip(n18878), .op(n18859) );
  mux2_1 U4646 ( .ip1(n4375), .ip2(n4374), .s(n18859), .op(n4378) );
  mux2_1 U4647 ( .ip1(\ANSWER/mem[8][9][1] ), .ip2(\ANSWER/mem[9][9][1] ), .s(
        n15643), .op(n4377) );
  inv_1 U4648 ( .ip(\CNTRL/count_20Q [4]), .op(n15184) );
  nor2_1 U4649 ( .ip1(\CNTRL/count_10Q [3]), .ip2(n15092), .op(n4376) );
  not_ab_or_c_or_d U4650 ( .ip1(n15092), .ip2(n15184), .ip3(n4376), .ip4(
        n15083), .op(n18252) );
  inv_1 U4651 ( .ip(n18252), .op(n18165) );
  inv_1 U4652 ( .ip(n18165), .op(n18227) );
  mux2_1 U4653 ( .ip1(n4378), .ip2(n4377), .s(n18227), .op(n4379) );
  nand2_1 U4654 ( .ip1(n18899), .ip2(n4379), .op(n4484) );
  inv_1 U4655 ( .ip(n4466), .op(n4453) );
  nor2_1 U4656 ( .ip1(n4453), .ip2(n18888), .op(n18914) );
  mux2_1 U4657 ( .ip1(\ANSWER/mem[0][8][1] ), .ip2(\ANSWER/mem[1][8][1] ), .s(
        n15643), .op(n4381) );
  mux2_1 U4658 ( .ip1(\ANSWER/mem[2][8][1] ), .ip2(\ANSWER/mem[3][8][1] ), .s(
        n15643), .op(n4380) );
  mux2_1 U4659 ( .ip1(n4381), .ip2(n4380), .s(n15636), .op(n4385) );
  mux2_1 U4660 ( .ip1(\ANSWER/mem[4][8][1] ), .ip2(\ANSWER/mem[5][8][1] ), .s(
        n15643), .op(n4383) );
  mux2_1 U4661 ( .ip1(\ANSWER/mem[6][8][1] ), .ip2(\ANSWER/mem[7][8][1] ), .s(
        n15643), .op(n4382) );
  mux2_1 U4662 ( .ip1(n4383), .ip2(n4382), .s(n15636), .op(n4384) );
  mux2_1 U4663 ( .ip1(n4385), .ip2(n4384), .s(n18859), .op(n4387) );
  mux2_1 U4664 ( .ip1(\ANSWER/mem[8][8][1] ), .ip2(\ANSWER/mem[9][8][1] ), .s(
        n15643), .op(n4386) );
  mux2_1 U4665 ( .ip1(n4387), .ip2(n4386), .s(n18227), .op(n4388) );
  nand2_1 U4666 ( .ip1(n18914), .ip2(n4388), .op(n4483) );
  nand2_1 U4667 ( .ip1(n15085), .ip2(\CNTRL/count_10_2Q [1]), .op(n4389) );
  nand2_1 U4668 ( .ip1(n4390), .ip2(n4389), .op(n4411) );
  inv_1 U4669 ( .ip(n4411), .op(n4465) );
  and2_1 U4670 ( .ip1(n15085), .ip2(\CNTRL/count_10_2Q [2]), .op(n4392) );
  nor2_1 U4671 ( .ip1(n4392), .ip2(n4391), .op(n4464) );
  nand2_1 U4672 ( .ip1(n4465), .ip2(n4464), .op(n15630) );
  nor2_1 U4673 ( .ip1(n15630), .ip2(n4466), .op(n18872) );
  and2_1 U4674 ( .ip1(n18888), .ip2(n18872), .op(n15648) );
  inv_1 U4675 ( .ip(n4362), .op(n17506) );
  buf_1 U4676 ( .ip(n17506), .op(n17536) );
  mux2_1 U4677 ( .ip1(\ANSWER/mem[0][1][1] ), .ip2(\ANSWER/mem[1][1][1] ), .s(
        n17536), .op(n4394) );
  mux2_1 U4678 ( .ip1(\ANSWER/mem[2][1][1] ), .ip2(\ANSWER/mem[3][1][1] ), .s(
        n17536), .op(n4393) );
  inv_1 U4679 ( .ip(n4366), .op(n4456) );
  mux2_1 U4680 ( .ip1(n4394), .ip2(n4393), .s(n4456), .op(n4398) );
  mux2_1 U4681 ( .ip1(\ANSWER/mem[4][1][1] ), .ip2(\ANSWER/mem[5][1][1] ), .s(
        n17536), .op(n4396) );
  mux2_1 U4682 ( .ip1(\ANSWER/mem[6][1][1] ), .ip2(\ANSWER/mem[7][1][1] ), .s(
        n17536), .op(n4395) );
  mux2_1 U4683 ( .ip1(n4396), .ip2(n4395), .s(n4456), .op(n4397) );
  mux2_1 U4684 ( .ip1(n4398), .ip2(n4397), .s(n18859), .op(n4400) );
  mux2_1 U4685 ( .ip1(\ANSWER/mem[8][1][1] ), .ip2(\ANSWER/mem[9][1][1] ), .s(
        n17536), .op(n4399) );
  mux2_1 U4686 ( .ip1(n4400), .ip2(n4399), .s(n18227), .op(n4401) );
  nand2_1 U4687 ( .ip1(n15648), .ip2(n4401), .op(n4482) );
  nor3_1 U4688 ( .ip1(n4411), .ip2(n4466), .ip3(n4464), .op(n18832) );
  mux2_1 U4689 ( .ip1(\ANSWER/mem[0][5][1] ), .ip2(\ANSWER/mem[1][5][1] ), .s(
        n17401), .op(n4403) );
  mux2_1 U4690 ( .ip1(\ANSWER/mem[2][5][1] ), .ip2(\ANSWER/mem[3][5][1] ), .s(
        n17401), .op(n4402) );
  mux2_1 U4691 ( .ip1(n4403), .ip2(n4402), .s(n4456), .op(n4407) );
  mux2_1 U4692 ( .ip1(\ANSWER/mem[4][5][1] ), .ip2(\ANSWER/mem[5][5][1] ), .s(
        n17401), .op(n4405) );
  mux2_1 U4693 ( .ip1(\ANSWER/mem[6][5][1] ), .ip2(\ANSWER/mem[7][5][1] ), .s(
        n17401), .op(n4404) );
  mux2_1 U4694 ( .ip1(n4405), .ip2(n4404), .s(n4456), .op(n4406) );
  mux2_1 U4695 ( .ip1(n4407), .ip2(n4406), .s(n18859), .op(n4409) );
  mux2_1 U4696 ( .ip1(\ANSWER/mem[8][5][1] ), .ip2(\ANSWER/mem[9][5][1] ), .s(
        n17401), .op(n4408) );
  mux2_1 U4697 ( .ip1(n4409), .ip2(n4408), .s(n18227), .op(n4410) );
  nand2_1 U4698 ( .ip1(n18832), .ip2(n4410), .op(n4442) );
  nor3_1 U4699 ( .ip1(n4411), .ip2(n4453), .ip3(n4464), .op(n18843) );
  mux2_1 U4700 ( .ip1(\ANSWER/mem[0][4][1] ), .ip2(\ANSWER/mem[1][4][1] ), .s(
        n15643), .op(n4413) );
  mux2_1 U4701 ( .ip1(\ANSWER/mem[2][4][1] ), .ip2(\ANSWER/mem[3][4][1] ), .s(
        n17401), .op(n4412) );
  mux2_1 U4702 ( .ip1(n4413), .ip2(n4412), .s(n4456), .op(n4417) );
  mux2_1 U4703 ( .ip1(\ANSWER/mem[4][4][1] ), .ip2(\ANSWER/mem[5][4][1] ), .s(
        n17401), .op(n4415) );
  mux2_1 U4704 ( .ip1(\ANSWER/mem[6][4][1] ), .ip2(\ANSWER/mem[7][4][1] ), .s(
        n17401), .op(n4414) );
  mux2_1 U4705 ( .ip1(n4415), .ip2(n4414), .s(n4456), .op(n4416) );
  mux2_1 U4706 ( .ip1(n4417), .ip2(n4416), .s(n18859), .op(n4419) );
  mux2_1 U4707 ( .ip1(\ANSWER/mem[8][4][1] ), .ip2(\ANSWER/mem[9][4][1] ), .s(
        n15643), .op(n4418) );
  mux2_1 U4708 ( .ip1(n4419), .ip2(n4418), .s(n18227), .op(n4420) );
  nand2_1 U4709 ( .ip1(n18843), .ip2(n4420), .op(n4441) );
  nor2_1 U4710 ( .ip1(n4453), .ip2(n15630), .op(n18800) );
  mux2_1 U4711 ( .ip1(\ANSWER/mem[0][0][1] ), .ip2(\ANSWER/mem[1][0][1] ), .s(
        n17536), .op(n4422) );
  mux2_1 U4712 ( .ip1(\ANSWER/mem[2][0][1] ), .ip2(\ANSWER/mem[3][0][1] ), .s(
        n17536), .op(n4421) );
  mux2_1 U4713 ( .ip1(n4422), .ip2(n4421), .s(n4456), .op(n4426) );
  mux2_1 U4714 ( .ip1(\ANSWER/mem[4][0][1] ), .ip2(\ANSWER/mem[5][0][1] ), .s(
        n17536), .op(n4424) );
  mux2_1 U4715 ( .ip1(\ANSWER/mem[6][0][1] ), .ip2(\ANSWER/mem[7][0][1] ), .s(
        n17536), .op(n4423) );
  mux2_1 U4716 ( .ip1(n4424), .ip2(n4423), .s(n4456), .op(n4425) );
  mux2_1 U4717 ( .ip1(n4426), .ip2(n4425), .s(n18859), .op(n4428) );
  mux2_1 U4718 ( .ip1(\ANSWER/mem[8][0][1] ), .ip2(\ANSWER/mem[9][0][1] ), .s(
        n17536), .op(n4427) );
  mux2_1 U4719 ( .ip1(n4428), .ip2(n4427), .s(n18227), .op(n4429) );
  nand2_1 U4720 ( .ip1(n18800), .ip2(n4429), .op(n4440) );
  inv_1 U4721 ( .ip(n4464), .op(n4452) );
  nor3_1 U4722 ( .ip1(n4452), .ip2(n4466), .ip3(n4465), .op(n18854) );
  mux2_1 U4723 ( .ip1(\ANSWER/mem[0][3][1] ), .ip2(\ANSWER/mem[1][3][1] ), .s(
        n17401), .op(n4431) );
  mux2_1 U4724 ( .ip1(\ANSWER/mem[2][3][1] ), .ip2(\ANSWER/mem[3][3][1] ), .s(
        n17401), .op(n4430) );
  mux2_1 U4725 ( .ip1(n4431), .ip2(n4430), .s(n4456), .op(n4435) );
  mux2_1 U4726 ( .ip1(\ANSWER/mem[4][3][1] ), .ip2(\ANSWER/mem[5][3][1] ), .s(
        n17401), .op(n4433) );
  mux2_1 U4727 ( .ip1(\ANSWER/mem[6][3][1] ), .ip2(\ANSWER/mem[7][3][1] ), .s(
        n17401), .op(n4432) );
  mux2_1 U4728 ( .ip1(n4433), .ip2(n4432), .s(n4456), .op(n4434) );
  mux2_1 U4729 ( .ip1(n4435), .ip2(n4434), .s(n18859), .op(n4437) );
  mux2_1 U4730 ( .ip1(\ANSWER/mem[8][3][1] ), .ip2(\ANSWER/mem[9][3][1] ), .s(
        n15643), .op(n4436) );
  mux2_1 U4731 ( .ip1(n4437), .ip2(n4436), .s(n18227), .op(n4438) );
  nand2_1 U4732 ( .ip1(n18854), .ip2(n4438), .op(n4439) );
  and4_1 U4733 ( .ip1(n4442), .ip2(n4441), .ip3(n4440), .ip4(n4439), .op(n4479) );
  nor3_1 U4734 ( .ip1(n4453), .ip2(n4465), .ip3(n4464), .op(n18821) );
  mux2_1 U4735 ( .ip1(\ANSWER/mem[0][6][1] ), .ip2(\ANSWER/mem[1][6][1] ), .s(
        n17401), .op(n4444) );
  mux2_1 U4736 ( .ip1(\ANSWER/mem[2][6][1] ), .ip2(\ANSWER/mem[3][6][1] ), .s(
        n17401), .op(n4443) );
  mux2_1 U4737 ( .ip1(n4444), .ip2(n4443), .s(n4456), .op(n4448) );
  mux2_1 U4738 ( .ip1(\ANSWER/mem[4][6][1] ), .ip2(\ANSWER/mem[5][6][1] ), .s(
        n17401), .op(n4446) );
  mux2_1 U4739 ( .ip1(\ANSWER/mem[6][6][1] ), .ip2(\ANSWER/mem[7][6][1] ), .s(
        n17401), .op(n4445) );
  mux2_1 U4740 ( .ip1(n4446), .ip2(n4445), .s(n15636), .op(n4447) );
  mux2_1 U4741 ( .ip1(n4448), .ip2(n4447), .s(n18859), .op(n4450) );
  mux2_1 U4742 ( .ip1(\ANSWER/mem[8][6][1] ), .ip2(\ANSWER/mem[9][6][1] ), .s(
        n17401), .op(n4449) );
  mux2_1 U4743 ( .ip1(n4450), .ip2(n4449), .s(n18227), .op(n4451) );
  nand2_1 U4744 ( .ip1(n18821), .ip2(n4451), .op(n4478) );
  nor3_1 U4745 ( .ip1(n4453), .ip2(n4452), .ip3(n4465), .op(n18884) );
  mux2_1 U4746 ( .ip1(\ANSWER/mem[0][2][1] ), .ip2(\ANSWER/mem[1][2][1] ), .s(
        n17536), .op(n4455) );
  mux2_1 U4747 ( .ip1(\ANSWER/mem[2][2][1] ), .ip2(\ANSWER/mem[3][2][1] ), .s(
        n17536), .op(n4454) );
  mux2_1 U4748 ( .ip1(n4455), .ip2(n4454), .s(n4456), .op(n4460) );
  mux2_1 U4749 ( .ip1(\ANSWER/mem[4][2][1] ), .ip2(\ANSWER/mem[5][2][1] ), .s(
        n17536), .op(n4458) );
  mux2_1 U4750 ( .ip1(\ANSWER/mem[6][2][1] ), .ip2(\ANSWER/mem[7][2][1] ), .s(
        n17401), .op(n4457) );
  mux2_1 U4751 ( .ip1(n4458), .ip2(n4457), .s(n4456), .op(n4459) );
  mux2_1 U4752 ( .ip1(n4460), .ip2(n4459), .s(n18859), .op(n4462) );
  mux2_1 U4753 ( .ip1(\ANSWER/mem[8][2][1] ), .ip2(\ANSWER/mem[9][2][1] ), .s(
        n15643), .op(n4461) );
  mux2_1 U4754 ( .ip1(n4462), .ip2(n4461), .s(n18227), .op(n4463) );
  nand2_1 U4755 ( .ip1(n18884), .ip2(n4463), .op(n4477) );
  nor3_1 U4756 ( .ip1(n4466), .ip2(n4465), .ip3(n4464), .op(n18865) );
  mux2_1 U4757 ( .ip1(\ANSWER/mem[0][7][1] ), .ip2(\ANSWER/mem[1][7][1] ), .s(
        n17401), .op(n4468) );
  mux2_1 U4758 ( .ip1(\ANSWER/mem[2][7][1] ), .ip2(\ANSWER/mem[3][7][1] ), .s(
        n17401), .op(n4467) );
  mux2_1 U4759 ( .ip1(n4468), .ip2(n4467), .s(n15636), .op(n4472) );
  mux2_1 U4760 ( .ip1(\ANSWER/mem[4][7][1] ), .ip2(\ANSWER/mem[5][7][1] ), .s(
        n17401), .op(n4470) );
  mux2_1 U4761 ( .ip1(\ANSWER/mem[6][7][1] ), .ip2(\ANSWER/mem[7][7][1] ), .s(
        n15643), .op(n4469) );
  mux2_1 U4762 ( .ip1(n4470), .ip2(n4469), .s(n15636), .op(n4471) );
  mux2_1 U4763 ( .ip1(n4472), .ip2(n4471), .s(n18859), .op(n4474) );
  mux2_1 U4764 ( .ip1(\ANSWER/mem[8][7][1] ), .ip2(\ANSWER/mem[9][7][1] ), .s(
        n15643), .op(n4473) );
  mux2_1 U4765 ( .ip1(n4474), .ip2(n4473), .s(n18227), .op(n4475) );
  nand2_1 U4766 ( .ip1(n18865), .ip2(n4475), .op(n4476) );
  nand4_1 U4767 ( .ip1(n4479), .ip2(n4478), .ip3(n4477), .ip4(n4476), .op(
        n4480) );
  nand2_1 U4768 ( .ip1(n18888), .ip2(n4480), .op(n4481) );
  nand4_1 U4769 ( .ip1(n4484), .ip2(n4483), .ip3(n4482), .ip4(n4481), .op(
        \ANSWER/N486 ) );
  inv_1 U4770 ( .ip(\CNTRL/currentState [1]), .op(n15086) );
  nor3_1 U4771 ( .ip1(\CNTRL/currentState [0]), .ip2(n15086), .ip3(n15083), 
        .op(n4495) );
  mux2_1 U4772 ( .ip1(m2DataIn[8]), .ip2(rdata[8]), .s(n4495), .op(n4488) );
  mux2_1 U4773 ( .ip1(m2DataIn[7]), .ip2(rdata[7]), .s(n4495), .op(n4535) );
  inv_1 U4774 ( .ip(m2DataIn[6]), .op(n16273) );
  inv_1 U4775 ( .ip(rdata[6]), .op(n16027) );
  mux2_1 U4776 ( .ip1(n16273), .ip2(n16027), .s(n4495), .op(n4527) );
  mux2_1 U4777 ( .ip1(m2DataIn[5]), .ip2(rdata[5]), .s(n4495), .op(n4522) );
  inv_1 U4778 ( .ip(m2DataIn[4]), .op(n16445) );
  inv_1 U4779 ( .ip(rdata[4]), .op(n15989) );
  mux2_1 U4780 ( .ip1(n16445), .ip2(n15989), .s(n4495), .op(n4519) );
  mux2_1 U4781 ( .ip1(m2DataIn[3]), .ip2(rdata[3]), .s(n4495), .op(n4515) );
  mux2_1 U4782 ( .ip1(m2DataIn[2]), .ip2(rdata[2]), .s(n4495), .op(n4512) );
  mux2_1 U4783 ( .ip1(m2DataIn[1]), .ip2(rdata[1]), .s(n4495), .op(n4509) );
  mux2_1 U4784 ( .ip1(m2DataIn[0]), .ip2(rdata[0]), .s(n4495), .op(n4516) );
  nor2_1 U4785 ( .ip1(n4509), .ip2(n4516), .op(n4510) );
  inv_1 U4786 ( .ip(n4510), .op(n4529) );
  nor2_1 U4787 ( .ip1(n4512), .ip2(n4529), .op(n4513) );
  inv_1 U4788 ( .ip(n4513), .op(n4485) );
  nor2_1 U4789 ( .ip1(n4515), .ip2(n4485), .op(n4517) );
  nand2_1 U4790 ( .ip1(n4519), .ip2(n4517), .op(n4520) );
  nor2_1 U4791 ( .ip1(n4522), .ip2(n4520), .op(n4524) );
  nand2_1 U4792 ( .ip1(n4527), .ip2(n4524), .op(n4533) );
  or2_1 U4793 ( .ip1(n4535), .ip2(n4533), .op(n4487) );
  mux2_1 U4794 ( .ip1(m2DataIn[15]), .ip2(rdata[15]), .s(n4495), .op(n18918)
         );
  nand2_1 U4795 ( .ip1(n4487), .ip2(n18918), .op(n4486) );
  xor2_1 U4796 ( .ip1(n4488), .ip2(n4486), .op(n4557) );
  inv_1 U4797 ( .ip(n4557), .op(n4588) );
  or2_1 U4798 ( .ip1(n4488), .ip2(n4487), .op(n15445) );
  nand2_1 U4799 ( .ip1(n18918), .ip2(n15445), .op(n4496) );
  inv_1 U4800 ( .ip(m2DataIn[9]), .op(n16690) );
  inv_1 U4801 ( .ip(rdata[9]), .op(n4489) );
  mux2_1 U4802 ( .ip1(n16690), .ip2(n4489), .s(n4495), .op(n4497) );
  xor2_1 U4803 ( .ip1(n4496), .ip2(n4497), .op(n15444) );
  mux2_1 U4804 ( .ip1(m2DataIn[11]), .ip2(rdata[11]), .s(n4495), .op(n4501) );
  mux2_1 U4805 ( .ip1(m2DataIn[12]), .ip2(rdata[12]), .s(n4495), .op(n4500) );
  or2_1 U4806 ( .ip1(n4501), .ip2(n4500), .op(n4494) );
  mux2_1 U4807 ( .ip1(m2DataIn[14]), .ip2(rdata[14]), .s(n4495), .op(n4491) );
  mux2_1 U4808 ( .ip1(m2DataIn[13]), .ip2(rdata[13]), .s(n4495), .op(n4490) );
  and3_1 U4809 ( .ip1(n4491), .ip2(n4494), .ip3(n4490), .op(n4493) );
  nor3_1 U4810 ( .ip1(n18918), .ip2(n4491), .ip3(n4490), .op(n4492) );
  nor2_1 U4811 ( .ip1(n4493), .ip2(n4492), .op(n4502) );
  or2_1 U4812 ( .ip1(n4494), .ip2(n4502), .op(n4505) );
  inv_1 U4813 ( .ip(m2DataIn[10]), .op(n16600) );
  inv_1 U4814 ( .ip(rdata[10]), .op(n16358) );
  mux2_1 U4815 ( .ip1(n16600), .ip2(n16358), .s(n4495), .op(n4506) );
  nand2_1 U4816 ( .ip1(n4497), .ip2(n4496), .op(n4498) );
  nand2_1 U4817 ( .ip1(n18918), .ip2(n4498), .op(n4507) );
  nand2_1 U4818 ( .ip1(n4506), .ip2(n4507), .op(n4499) );
  nand4_1 U4819 ( .ip1(n18918), .ip2(n4501), .ip3(n4500), .ip4(n4499), .op(
        n4503) );
  or2_1 U4820 ( .ip1(n4503), .ip2(n4502), .op(n4504) );
  nand2_1 U4821 ( .ip1(n4505), .ip2(n4504), .op(n15447) );
  inv_1 U4822 ( .ip(n15447), .op(n4559) );
  xor2_1 U4823 ( .ip1(n4507), .ip2(n4506), .op(n15443) );
  nor2_1 U4824 ( .ip1(n4559), .ip2(n15443), .op(n4562) );
  nand2_1 U4825 ( .ip1(n15444), .ip2(n4562), .op(n15428) );
  nor2_1 U4826 ( .ip1(n4588), .ip2(n15428), .op(n4570) );
  nand2_1 U4827 ( .ip1(n18918), .ip2(n4516), .op(n4508) );
  xnor2_1 U4828 ( .ip1(n4509), .ip2(n4508), .op(n4542) );
  inv_1 U4829 ( .ip(n18918), .op(n4525) );
  nor2_1 U4830 ( .ip1(n4525), .ip2(n4510), .op(n4511) );
  xor2_1 U4831 ( .ip1(n4512), .ip2(n4511), .op(n4543) );
  nor2_1 U4832 ( .ip1(n4525), .ip2(n4513), .op(n4514) );
  xor2_1 U4833 ( .ip1(n4515), .ip2(n4514), .op(n4545) );
  not_ab_or_c_or_d U4834 ( .ip1(n4516), .ip2(n4542), .ip3(n4543), .ip4(n4545), 
        .op(n4523) );
  or2_1 U4835 ( .ip1(n4517), .ip2(n4525), .op(n4518) );
  xor2_1 U4836 ( .ip1(n4519), .ip2(n4518), .op(n4546) );
  inv_1 U4837 ( .ip(n4546), .op(n4531) );
  nand2_1 U4838 ( .ip1(n4520), .ip2(n18918), .op(n4521) );
  xor2_1 U4839 ( .ip1(n4522), .ip2(n4521), .op(n4548) );
  nor3_1 U4840 ( .ip1(n4523), .ip2(n4531), .ip3(n4548), .op(n4528) );
  nor2_1 U4841 ( .ip1(n4525), .ip2(n4524), .op(n4526) );
  xnor2_1 U4842 ( .ip1(n4527), .ip2(n4526), .op(n4553) );
  nor2_1 U4843 ( .ip1(n4528), .ip2(n4553), .op(n4583) );
  inv_1 U4844 ( .ip(n4583), .op(n4563) );
  nand3_1 U4845 ( .ip1(n4529), .ip2(n4543), .ip3(n4545), .op(n4530) );
  nand3_1 U4846 ( .ip1(n4531), .ip2(n4548), .ip3(n4530), .op(n4532) );
  nand2_1 U4847 ( .ip1(n4553), .ip2(n4532), .op(n15465) );
  nand2_1 U4848 ( .ip1(n4563), .ip2(n15465), .op(n4549) );
  inv_1 U4849 ( .ip(n4549), .op(n15474) );
  nand2_1 U4850 ( .ip1(n4533), .ip2(n18918), .op(n4534) );
  xor2_1 U4851 ( .ip1(n4535), .ip2(n4534), .op(n4589) );
  inv_1 U4852 ( .ip(n4589), .op(n15468) );
  inv_1 U4853 ( .ip(n4570), .op(n4568) );
  nor2_1 U4854 ( .ip1(n15468), .ip2(n4568), .op(n15464) );
  nand2_1 U4855 ( .ip1(n15468), .ip2(n4563), .op(n4536) );
  nand2_1 U4856 ( .ip1(n4557), .ip2(n4536), .op(n15420) );
  nor3_1 U4857 ( .ip1(n4589), .ip2(n15428), .ip3(n15420), .op(n15454) );
  not_ab_or_c_or_d U4858 ( .ip1(n4570), .ip2(n15474), .ip3(n15464), .ip4(
        n15454), .op(n15493) );
  inv_1 U4859 ( .ip(n15444), .op(n4558) );
  and2_1 U4860 ( .ip1(n4558), .ip2(n4562), .op(n4592) );
  nand2_1 U4861 ( .ip1(n4592), .ip2(n4588), .op(n4576) );
  inv_1 U4862 ( .ip(n4576), .op(n15475) );
  nand2_1 U4863 ( .ip1(n4589), .ip2(n15474), .op(n4551) );
  not_ab_or_c_or_d U4864 ( .ip1(n4543), .ip2(n4542), .ip3(n4546), .ip4(n4545), 
        .op(n4537) );
  nor2_1 U4865 ( .ip1(n4548), .ip2(n4537), .op(n4538) );
  nand2_1 U4866 ( .ip1(n4538), .ip2(n4553), .op(n4587) );
  inv_1 U4867 ( .ip(n4587), .op(n15437) );
  nand2_1 U4868 ( .ip1(n4589), .ip2(n15437), .op(n4574) );
  nor2_1 U4869 ( .ip1(n15465), .ip2(n4538), .op(n4584) );
  inv_1 U4870 ( .ip(n4584), .op(n4539) );
  nor2_1 U4871 ( .ip1(n15468), .ip2(n4539), .op(n15427) );
  inv_1 U4872 ( .ip(n15427), .op(n4540) );
  nand3_1 U4873 ( .ip1(n4551), .ip2(n4574), .ip3(n4540), .op(n4541) );
  nand2_1 U4874 ( .ip1(n15475), .ip2(n4541), .op(n15419) );
  or2_1 U4875 ( .ip1(n4543), .ip2(n4542), .op(n4544) );
  nand3_1 U4876 ( .ip1(n4546), .ip2(n4545), .ip3(n4544), .op(n4547) );
  nand2_1 U4877 ( .ip1(n4548), .ip2(n4547), .op(n4554) );
  nand2_1 U4878 ( .ip1(n4583), .ip2(n4554), .op(n4550) );
  nor2_1 U4879 ( .ip1(n4589), .ip2(n4550), .op(n15417) );
  nand2_1 U4880 ( .ip1(n4557), .ip2(n4592), .op(n15467) );
  inv_1 U4881 ( .ip(n15467), .op(n4573) );
  nand2_1 U4882 ( .ip1(n15417), .ip2(n4573), .op(n15415) );
  nor2_1 U4883 ( .ip1(n4549), .ip2(n15467), .op(n15442) );
  nand2_1 U4884 ( .ip1(n15442), .ip2(n15468), .op(n4594) );
  and2_1 U4885 ( .ip1(n15415), .ip2(n4594), .op(n4552) );
  nor2_1 U4886 ( .ip1(n15468), .ip2(n4550), .op(n15435) );
  inv_1 U4887 ( .ip(n15435), .op(n15466) );
  nand2_1 U4888 ( .ip1(n4551), .ip2(n15466), .op(n15455) );
  nand2_1 U4889 ( .ip1(n4573), .ip2(n15455), .op(n15485) );
  nand4_1 U4890 ( .ip1(n15493), .ip2(n15419), .ip3(n4552), .ip4(n15485), .op(
        n3906) );
  nor2_1 U4891 ( .ip1(n4554), .ip2(n4553), .op(n4578) );
  nand2_1 U4892 ( .ip1(n4589), .ip2(n4578), .op(n4575) );
  nor2_1 U4893 ( .ip1(n4588), .ip2(n4575), .op(n15429) );
  inv_1 U4894 ( .ip(n15443), .op(n15423) );
  or2_1 U4895 ( .ip1(n15429), .ip2(n15423), .op(n4556) );
  or2_1 U4896 ( .ip1(n4558), .ip2(n15423), .op(n4555) );
  nand2_1 U4897 ( .ip1(n4556), .ip2(n4555), .op(n4566) );
  nand3_1 U4898 ( .ip1(n4557), .ip2(n4589), .ip3(n15465), .op(n15421) );
  nor3_1 U4899 ( .ip1(n15444), .ip2(n4559), .ip3(n15421), .op(n4565) );
  nor2_1 U4900 ( .ip1(n4558), .ip2(n4557), .op(n4561) );
  nor2_1 U4901 ( .ip1(n4589), .ip2(n4587), .op(n4569) );
  nand2_1 U4902 ( .ip1(n4561), .ip2(n4569), .op(n4560) );
  not_ab_or_c_or_d U4903 ( .ip1(n15423), .ip2(n4560), .ip3(n4566), .ip4(n4559), 
        .op(n15426) );
  and2_1 U4904 ( .ip1(n4562), .ip2(n4561), .op(n15470) );
  nand2_1 U4905 ( .ip1(n15417), .ip2(n15470), .op(n15431) );
  nand4_1 U4906 ( .ip1(n15470), .ip2(n15468), .ip3(n4563), .ip4(n4587), .op(
        n4564) );
  nand2_1 U4907 ( .ip1(n15431), .ip2(n4564), .op(n15462) );
  not_ab_or_c_or_d U4908 ( .ip1(n4566), .ip2(n4565), .ip3(n15426), .ip4(n15462), .op(n15491) );
  and2_1 U4909 ( .ip1(n4584), .ip2(n15464), .op(n15456) );
  or2_1 U4910 ( .ip1(n15437), .ip2(n15456), .op(n4567) );
  nand2_1 U4911 ( .ip1(n15464), .ip2(n4567), .op(n15433) );
  nand2_1 U4912 ( .ip1(n15468), .ip2(n4584), .op(n4577) );
  nor2_1 U4913 ( .ip1(n4577), .ip2(n4568), .op(n15463) );
  or2_1 U4914 ( .ip1(n4569), .ip2(n15463), .op(n4571) );
  nand2_1 U4915 ( .ip1(n4571), .ip2(n4570), .op(n15472) );
  nand3_1 U4916 ( .ip1(n4578), .ip2(n15470), .ip3(n4589), .op(n4572) );
  nand2_1 U4917 ( .ip1(n15472), .ip2(n4572), .op(n4582) );
  nand2_1 U4918 ( .ip1(n15427), .ip2(n4573), .op(n15476) );
  or2_1 U4919 ( .ip1(n4574), .ip2(n15467), .op(n15449) );
  nand2_1 U4920 ( .ip1(n15476), .ip2(n15449), .op(n4590) );
  inv_1 U4921 ( .ip(n4590), .op(n4580) );
  nor2_1 U4922 ( .ip1(n4576), .ip2(n4575), .op(n15441) );
  nor2_1 U4923 ( .ip1(n15467), .ip2(n4577), .op(n15413) );
  nor2_1 U4924 ( .ip1(n15441), .ip2(n15413), .op(n4596) );
  inv_1 U4925 ( .ip(n4578), .op(n15469) );
  nand2_1 U4926 ( .ip1(n15475), .ip2(n15468), .op(n15436) );
  nor2_1 U4927 ( .ip1(n15469), .ip2(n15436), .op(n15416) );
  inv_1 U4928 ( .ip(n15416), .op(n4579) );
  nand4_1 U4929 ( .ip1(n4580), .ip2(n4596), .ip3(n4579), .ip4(n4594), .op(
        n4581) );
  not_ab_or_c_or_d U4930 ( .ip1(n4583), .ip2(n15464), .ip3(n4582), .ip4(n4581), 
        .op(n4586) );
  nand2_1 U4931 ( .ip1(n15475), .ip2(n4584), .op(n4585) );
  nand4_1 U4932 ( .ip1(n15491), .ip2(n15433), .ip3(n4586), .ip4(n4585), .op(
        n3908) );
  nor3_1 U4933 ( .ip1(n4589), .ip2(n4587), .ip3(n15467), .op(n15451) );
  nor3_1 U4934 ( .ip1(n4589), .ip2(n4588), .ip3(n15469), .op(n15425) );
  or2_1 U4935 ( .ip1(n15425), .ip2(n4590), .op(n4591) );
  nand2_1 U4936 ( .ip1(n4592), .ip2(n4591), .op(n15486) );
  nand2_1 U4937 ( .ip1(n15486), .ip2(n15485), .op(n4593) );
  not_ab_or_c_or_d U4938 ( .ip1(n15435), .ip2(n15475), .ip3(n15451), .ip4(
        n4593), .op(n4595) );
  nand4_1 U4939 ( .ip1(n4596), .ip2(n4595), .ip3(n15415), .ip4(n4594), .op(
        n3904) );
  nand2_1 U4940 ( .ip1(\CNTRL/currentState [0]), .ip2(\CNTRL/currentState [1]), 
        .op(n15094) );
  nor2_1 U4941 ( .ip1(n15083), .ip2(n15094), .op(n16714) );
  nor2_1 U4942 ( .ip1(\CNTRL/count_20Q [2]), .ip2(\CNTRL/count_20Q [3]), .op(
        n15185) );
  nand2_1 U4943 ( .ip1(\CNTRL/count_20Q [4]), .ip2(n15185), .op(n15167) );
  nand2_1 U4944 ( .ip1(\CNTRL/count_20Q [0]), .ip2(\CNTRL/count_20Q [1]), .op(
        n15100) );
  nor2_1 U4945 ( .ip1(n15167), .ip2(n15100), .op(n15091) );
  inv_1 U4946 ( .ip(n15091), .op(n4597) );
  nor2_1 U4947 ( .ip1(n15094), .ip2(n4597), .op(n4598) );
  nor4_1 U4948 ( .ip1(n15092), .ip2(n16714), .ip3(reset), .ip4(n4598), .op(
        n4108) );
  inv_1 U4949 ( .ip(\CNTRL/currentState [0]), .op(n15058) );
  nor2_1 U4950 ( .ip1(\CNTRL/currentState [2]), .ip2(n15058), .op(n4599) );
  nor3_1 U4951 ( .ip1(n15624), .ip2(reset), .ip3(n4599), .op(n15099) );
  inv_1 U4952 ( .ip(reset), .op(n15159) );
  nand3_1 U4953 ( .ip1(\CNTRL/currentState [1]), .ip2(\CNTRL/currentState [0]), 
        .ip3(n15083), .op(n4600) );
  nand2_1 U4954 ( .ip1(n15087), .ip2(n4600), .op(n4601) );
  nand2_1 U4955 ( .ip1(n15159), .ip2(n4601), .op(n15098) );
  nor2_1 U4956 ( .ip1(n15091), .ip2(n15098), .op(n15108) );
  or2_1 U4957 ( .ip1(n15099), .ip2(n15108), .op(n4603) );
  or2_1 U4958 ( .ip1(n15094), .ip2(n15108), .op(n4602) );
  nand2_1 U4959 ( .ip1(n4603), .ip2(n4602), .op(n15140) );
  inv_1 U4960 ( .ip(n16714), .op(n15052) );
  nand2_1 U4961 ( .ip1(n15624), .ip2(n15091), .op(n15051) );
  inv_1 U4962 ( .ip(\CNTRL/count_10Q [3]), .op(n15139) );
  nor4_1 U4963 ( .ip1(\CNTRL/count_10Q [2]), .ip2(\CNTRL/count_10Q [1]), .ip3(
        n15132), .ip4(n15139), .op(n15113) );
  not_ab_or_c_or_d U4964 ( .ip1(n15052), .ip2(n15051), .ip3(n15113), .ip4(
        reset), .op(n15131) );
  nand2_1 U4965 ( .ip1(n15131), .ip2(n15132), .op(n4605) );
  nand2_1 U4966 ( .ip1(n15140), .ip2(n4605), .op(n15133) );
  inv_1 U4967 ( .ip(n15133), .op(n4604) );
  or2_1 U4968 ( .ip1(n15132), .ip2(n4604), .op(n4606) );
  nand2_1 U4969 ( .ip1(n4606), .ip2(n4605), .op(n4098) );
  inv_1 U4970 ( .ip(n15099), .op(n15102) );
  inv_1 U4971 ( .ip(n15100), .op(n15109) );
  nand3_1 U4972 ( .ip1(\CNTRL/count_20Q [2]), .ip2(\CNTRL/count_20Q [3]), 
        .ip3(n15109), .op(n4607) );
  nand2_1 U4973 ( .ip1(n15108), .ip2(n4607), .op(n4608) );
  nand2_1 U4974 ( .ip1(n15102), .ip2(n4608), .op(n15089) );
  inv_1 U4975 ( .ip(n15089), .op(n4609) );
  or2_1 U4976 ( .ip1(n15174), .ip2(n4609), .op(n4612) );
  nand3_1 U4977 ( .ip1(\CNTRL/count_20Q [2]), .ip2(n15109), .ip3(n15108), .op(
        n4610) );
  or2_1 U4978 ( .ip1(n4610), .ip2(n4609), .op(n4611) );
  nand2_1 U4979 ( .ip1(n4612), .ip2(n4611), .op(n4103) );
  buf_1 U4980 ( .ip(\STAGE_1/weightReg [1]), .op(n13707) );
  buf_1 U4981 ( .ip(n13707), .op(n10507) );
  inv_1 U4982 ( .ip(\STAGE_1/weightReg [0]), .op(n10476) );
  buf_1 U4983 ( .ip(n10476), .op(n13646) );
  inv_1 U4984 ( .ip(\STAGE_1/weightReg [3]), .op(n13801) );
  inv_1 U4985 ( .ip(m1Inputs[130]), .op(n9461) );
  inv_1 U4986 ( .ip(m1Inputs[133]), .op(n9299) );
  nor4_1 U4987 ( .ip1(n10476), .ip2(n13801), .ip3(n9461), .ip4(n9299), .op(
        n4613) );
  inv_1 U4988 ( .ip(n4613), .op(n4618) );
  nand2_1 U4989 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[133]), .op(n4652) );
  or2_1 U4990 ( .ip1(n4652), .ip2(n4613), .op(n4616) );
  buf_1 U4991 ( .ip(\STAGE_1/weightReg [3]), .op(n9733) );
  nand2_1 U4992 ( .ip1(n9733), .ip2(m1Inputs[130]), .op(n4614) );
  or2_1 U4993 ( .ip1(n4614), .ip2(n4613), .op(n4615) );
  nand2_1 U4994 ( .ip1(n4616), .ip2(n4615), .op(n4690) );
  inv_1 U4995 ( .ip(m1Inputs[128]), .op(n9509) );
  nor2_1 U4996 ( .ip1(n9509), .ip2(n13835), .op(n4689) );
  nand2_1 U4997 ( .ip1(n4690), .ip2(n4689), .op(n4617) );
  nand2_1 U4998 ( .ip1(n4618), .ip2(n4617), .op(n4681) );
  nand2_1 U4999 ( .ip1(n4672), .ip2(m1Inputs[132]), .op(n4620) );
  buf_1 U5000 ( .ip(\STAGE_1/weightReg [2]), .op(n4619) );
  inv_1 U5001 ( .ip(n4619), .op(n6745) );
  inv_1 U5002 ( .ip(\STAGE_1/weightReg [1]), .op(n9047) );
  inv_1 U5003 ( .ip(m1Inputs[132]), .op(n9530) );
  nor4_1 U5004 ( .ip1(n6745), .ip2(n9047), .ip3(n9530), .ip4(n9299), .op(n4670) );
  or2_1 U5005 ( .ip1(n4620), .ip2(n4670), .op(n4623) );
  nand2_1 U5006 ( .ip1(n13707), .ip2(m1Inputs[133]), .op(n4621) );
  or2_1 U5007 ( .ip1(n4621), .ip2(n4670), .op(n4622) );
  nand2_1 U5008 ( .ip1(n4623), .ip2(n4622), .op(n4680) );
  inv_1 U5009 ( .ip(m1Inputs[129]), .op(n9540) );
  nor2_1 U5010 ( .ip1(n9540), .ip2(n4624), .op(n4647) );
  inv_1 U5011 ( .ip(m1Inputs[134]), .op(n14587) );
  nor2_1 U5012 ( .ip1(n10476), .ip2(n14587), .op(n8946) );
  inv_1 U5013 ( .ip(\STAGE_1/weightReg [6]), .op(n14289) );
  nor2_1 U5014 ( .ip1(n9509), .ip2(n14289), .op(n4646) );
  and3_1 U5015 ( .ip1(n13707), .ip2(m1Inputs[134]), .ip3(n4666), .op(n8984) );
  inv_1 U5016 ( .ip(m1Inputs[131]), .op(n9154) );
  nand2_1 U5017 ( .ip1(m1Inputs[130]), .ip2(\STAGE_1/weightReg [4]), .op(n4683) );
  inv_1 U5018 ( .ip(\STAGE_1/weightReg [5]), .op(n4624) );
  inv_1 U5019 ( .ip(n4624), .op(n12699) );
  inv_1 U5020 ( .ip(n12699), .op(n8942) );
  nor3_1 U5021 ( .ip1(n9154), .ip2(n4683), .ip3(n8942), .op(n4637) );
  nor2_1 U5022 ( .ip1(n9154), .ip2(n14783), .op(n4648) );
  or2_1 U5023 ( .ip1(n14369), .ip2(n4648), .op(n4626) );
  or2_1 U5024 ( .ip1(m1Inputs[130]), .ip2(n4648), .op(n4625) );
  nand2_1 U5025 ( .ip1(n4626), .ip2(n4625), .op(n4636) );
  inv_1 U5026 ( .ip(\STAGE_1/weightReg [7]), .op(n12156) );
  buf_1 U5027 ( .ip(n12156), .op(n14384) );
  inv_1 U5028 ( .ip(n14384), .op(n4627) );
  buf_1 U5029 ( .ip(n12156), .op(n14368) );
  inv_1 U5030 ( .ip(n14368), .op(n14835) );
  nand2_1 U5031 ( .ip1(m1Inputs[128]), .ip2(n14835), .op(n4638) );
  nor2_1 U5032 ( .ip1(n4636), .ip2(n4638), .op(n4628) );
  nor2_1 U5033 ( .ip1(n4637), .ip2(n4628), .op(n8953) );
  nand2_1 U5034 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[135]), .op(n9504) );
  buf_1 U5035 ( .ip(\STAGE_1/weightReg [3]), .op(n12578) );
  nor2_1 U5036 ( .ip1(n10476), .ip2(n9530), .op(n4701) );
  and3_1 U5037 ( .ip1(n12578), .ip2(m1Inputs[135]), .ip3(n4701), .op(n4632) );
  or2_1 U5038 ( .ip1(n9504), .ip2(n4632), .op(n4631) );
  nand2_1 U5039 ( .ip1(n12578), .ip2(m1Inputs[132]), .op(n4629) );
  or2_1 U5040 ( .ip1(n4629), .ip2(n4632), .op(n4630) );
  nand2_1 U5041 ( .ip1(n4631), .ip2(n4630), .op(n4644) );
  or2_1 U5042 ( .ip1(n4644), .ip2(n4632), .op(n4634) );
  nor2_1 U5043 ( .ip1(n6745), .ip2(n9299), .op(n4643) );
  or2_1 U5044 ( .ip1(n4643), .ip2(n4632), .op(n4633) );
  nand2_1 U5045 ( .ip1(n4634), .ip2(n4633), .op(n8952) );
  nand2_1 U5046 ( .ip1(m1Inputs[130]), .ip2(\STAGE_1/weightReg [6]), .op(n8951) );
  inv_1 U5047 ( .ip(n4635), .op(n8981) );
  nor2_1 U5048 ( .ip1(n4637), .ip2(n4636), .op(n4639) );
  xor2_1 U5049 ( .ip1(n4639), .ip2(n4638), .op(n4664) );
  inv_1 U5050 ( .ip(\STAGE_1/weightReg [3]), .op(n13082) );
  nand4_1 U5051 ( .ip1(n4619), .ip2(\STAGE_1/weightReg [1]), .ip3(
        m1Inputs[131]), .ip4(m1Inputs[132]), .op(n4673) );
  nor2_1 U5052 ( .ip1(n13082), .ip2(n4673), .op(n4642) );
  nand2_1 U5053 ( .ip1(n4673), .ip2(m1Inputs[131]), .op(n4640) );
  mux2_1 U5054 ( .ip1(n4673), .ip2(n4640), .s(n9733), .op(n4682) );
  nor2_1 U5055 ( .ip1(n4683), .ip2(n4682), .op(n4641) );
  nor2_1 U5056 ( .ip1(n4642), .ip2(n4641), .op(n4663) );
  xnor2_1 U5057 ( .ip1(n4644), .ip2(n4643), .op(n4662) );
  inv_1 U5058 ( .ip(n4645), .op(n8980) );
  buf_1 U5059 ( .ip(n14289), .op(n14836) );
  nor2_1 U5060 ( .ip1(n9540), .ip2(n14836), .op(n4671) );
  fulladder U5061 ( .a(n4647), .b(n8946), .ci(n4646), .co(n4669), .s(n4679) );
  nand2_1 U5062 ( .ip1(m1Inputs[131]), .ip2(\STAGE_1/weightReg [5]), .op(n4649) );
  and3_1 U5063 ( .ip1(m1Inputs[132]), .ip2(\STAGE_1/weightReg [5]), .ip3(n4648), .op(n8967) );
  or2_1 U5064 ( .ip1(n4649), .ip2(n8967), .op(n4651) );
  nand2_1 U5065 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[132]), .op(n8941) );
  or2_1 U5066 ( .ip1(n8941), .ip2(n8967), .op(n4650) );
  nand2_1 U5067 ( .ip1(n4651), .ip2(n4650), .op(n8966) );
  nor2_1 U5068 ( .ip1(n9540), .ip2(n14384), .op(n8968) );
  xor2_1 U5069 ( .ip1(n8966), .ip2(n8968), .op(n8978) );
  nand2_1 U5070 ( .ip1(n9733), .ip2(m1Inputs[133]), .op(n4653) );
  inv_1 U5071 ( .ip(m1Inputs[136]), .op(n14635) );
  nor3_1 U5072 ( .ip1(n13801), .ip2(n14635), .ip3(n4652), .op(n8962) );
  or2_1 U5073 ( .ip1(n4653), .ip2(n8962), .op(n4655) );
  nand2_1 U5074 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[136]), .op(n9448) );
  or2_1 U5075 ( .ip1(n9448), .ip2(n8962), .op(n4654) );
  nand2_1 U5076 ( .ip1(n4655), .ip2(n4654), .op(n8961) );
  inv_1 U5077 ( .ip(\STAGE_1/weightReg [8]), .op(n6503) );
  nor2_1 U5078 ( .ip1(n9509), .ip2(n6503), .op(n8963) );
  xor2_1 U5079 ( .ip1(n8961), .ip2(n8963), .op(n8977) );
  nand2_1 U5080 ( .ip1(m1Inputs[134]), .ip2(n4672), .op(n4656) );
  nand2_1 U5081 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[135]), .op(n8971) );
  nand2_1 U5082 ( .ip1(n4656), .ip2(n8971), .op(n4657) );
  nand4_1 U5083 ( .ip1(\STAGE_1/weightReg [2]), .ip2(\STAGE_1/weightReg [1]), 
        .ip3(m1Inputs[135]), .ip4(m1Inputs[134]), .op(n8955) );
  nand2_1 U5084 ( .ip1(n4657), .ip2(n8955), .op(n8957) );
  nor3_1 U5085 ( .ip1(n15058), .ip2(\CNTRL/currentState [1]), .ip3(
        \CNTRL/currentState [2]), .op(n17289) );
  buf_1 U5086 ( .ip(n17289), .op(n17229) );
  inv_1 U5087 ( .ip(\CNTRL/count_layer1_784Q [6]), .op(n15074) );
  nand3_1 U5088 ( .ip1(n15092), .ip2(n15083), .ip3(n15074), .op(n4658) );
  nor4_1 U5089 ( .ip1(\CNTRL/count_layer1_784Q [4]), .ip2(
        \CNTRL/count_layer1_784Q [7]), .ip3(\CNTRL/count_layer1_784Q [5]), 
        .ip4(n4658), .op(n15047) );
  nor2_1 U5090 ( .ip1(\CNTRL/count_layer1_784Q [0]), .ip2(
        \CNTRL/count_layer1_784Q [1]), .op(n15061) );
  inv_1 U5091 ( .ip(\CNTRL/count_layer1_784Q [8]), .op(n15079) );
  inv_1 U5092 ( .ip(\CNTRL/count_layer1_784Q [9]), .op(n4659) );
  nand4_1 U5093 ( .ip1(n15047), .ip2(n15061), .ip3(n15079), .ip4(n4659), .op(
        n4660) );
  nor3_1 U5094 ( .ip1(\CNTRL/count_layer1_784Q [3]), .ip2(n4660), .ip3(
        \CNTRL/count_layer1_784Q [2]), .op(n4661) );
  nor2_1 U5095 ( .ip1(n17229), .ip2(n4661), .op(n14768) );
  nand2_1 U5096 ( .ip1(column[128]), .ip2(n13498), .op(n8956) );
  xor2_1 U5097 ( .ip1(n8957), .ip2(n8956), .op(n8976) );
  fulladder U5098 ( .a(n4664), .b(n4663), .ci(n4662), .co(n4645), .s(n4665) );
  inv_1 U5099 ( .ip(n4665), .op(n4748) );
  nor2_1 U5100 ( .ip1(n9047), .ip2(n14587), .op(n4667) );
  nor2_1 U5101 ( .ip1(n4667), .ip2(n4666), .op(n4668) );
  nor2_1 U5102 ( .ip1(n8984), .ip2(n4668), .op(n4747) );
  fulladder U5103 ( .a(n4671), .b(n4670), .ci(n4669), .co(n8979), .s(n4746) );
  buf_1 U5104 ( .ip(\STAGE_1/weightReg [2]), .op(n4672) );
  inv_1 U5105 ( .ip(n4672), .op(n10555) );
  nand2_1 U5106 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[130]), .op(n4702) );
  nor3_1 U5107 ( .ip1(n10555), .ip2(n9154), .ip3(n4702), .op(n4698) );
  inv_1 U5108 ( .ip(n4673), .op(n4678) );
  nor2_1 U5109 ( .ip1(n6745), .ip2(n9154), .op(n4674) );
  or2_1 U5110 ( .ip1(m1Inputs[132]), .ip2(n4674), .op(n4676) );
  or2_1 U5111 ( .ip1(n13707), .ip2(n4674), .op(n4675) );
  nand2_1 U5112 ( .ip1(n4676), .ip2(n4675), .op(n4677) );
  nor2_1 U5113 ( .ip1(n4678), .ip2(n4677), .op(n4688) );
  nor2_1 U5114 ( .ip1(n9540), .ip2(n14783), .op(n4687) );
  fulladder U5115 ( .a(n4681), .b(n4680), .ci(n4679), .co(n4666), .s(n4685) );
  xor2_1 U5116 ( .ip1(n4683), .ip2(n4682), .op(n4684) );
  nand2_1 U5117 ( .ip1(n4740), .ip2(n4739), .op(n4745) );
  fulladder U5118 ( .a(n4686), .b(n4685), .ci(n4684), .co(n4739), .s(n4734) );
  fulladder U5119 ( .a(n4698), .b(n4688), .ci(n4687), .co(n4686), .s(n4693) );
  nor2_1 U5120 ( .ip1(n13082), .ip2(n9540), .op(n4700) );
  inv_1 U5121 ( .ip(\STAGE_1/weightReg [4]), .op(n14783) );
  nor2_1 U5122 ( .ip1(n9509), .ip2(n14783), .op(n4699) );
  xor2_1 U5123 ( .ip1(n4690), .ip2(n4689), .op(n4691) );
  or2_1 U5124 ( .ip1(n4734), .ip2(n4733), .op(n4743) );
  fulladder U5125 ( .a(n4693), .b(n4692), .ci(n4691), .co(n4733), .s(n4732) );
  inv_1 U5126 ( .ip(\STAGE_1/weightReg [1]), .op(n13570) );
  nor4_1 U5127 ( .ip1(n13570), .ip2(n13082), .ip3(n9509), .ip4(n9461), .op(
        n4729) );
  nor2_1 U5128 ( .ip1(n13570), .ip2(n9154), .op(n4694) );
  or2_1 U5129 ( .ip1(m1Inputs[130]), .ip2(n4694), .op(n4696) );
  or2_1 U5130 ( .ip1(n4619), .ip2(n4694), .op(n4695) );
  nand2_1 U5131 ( .ip1(n4696), .ip2(n4695), .op(n4697) );
  nor2_1 U5132 ( .ip1(n4698), .ip2(n4697), .op(n4728) );
  fulladder U5133 ( .a(n4701), .b(n4700), .ci(n4699), .co(n4692), .s(n4727) );
  or2_1 U5134 ( .ip1(n4702), .ip2(n4729), .op(n4705) );
  nand2_1 U5135 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[128]), .op(n4703) );
  or2_1 U5136 ( .ip1(n4703), .ip2(n4729), .op(n4704) );
  nand2_1 U5137 ( .ip1(n4705), .ip2(n4704), .op(n4712) );
  nand2_1 U5138 ( .ip1(n4619), .ip2(m1Inputs[128]), .op(n4707) );
  nand2_1 U5139 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[129]), .op(n4706) );
  not_ab_or_c_or_d U5140 ( .ip1(n4707), .ip2(n4706), .ip3(n13646), .ip4(n9461), 
        .op(n4709) );
  buf_1 U5141 ( .ip(\STAGE_1/weightReg [0]), .op(n13803) );
  nand2_1 U5142 ( .ip1(n13803), .ip2(n6745), .op(n5739) );
  nor4_1 U5143 ( .ip1(n13570), .ip2(n5739), .ip3(n9509), .ip4(n9540), .op(
        n4708) );
  or2_1 U5144 ( .ip1(n4709), .ip2(n4708), .op(n4714) );
  nand2_1 U5145 ( .ip1(n4712), .ip2(n4714), .op(n4717) );
  nand2_1 U5146 ( .ip1(n4619), .ip2(m1Inputs[129]), .op(n4711) );
  nor2_1 U5147 ( .ip1(n10476), .ip2(n9154), .op(n4719) );
  nor4_1 U5148 ( .ip1(n6745), .ip2(n13570), .ip3(n9509), .ip4(n9540), .op(
        n4718) );
  xnor2_1 U5149 ( .ip1(n4719), .ip2(n4718), .op(n4710) );
  xor2_1 U5150 ( .ip1(n4711), .ip2(n4710), .op(n4713) );
  nand2_1 U5151 ( .ip1(n4712), .ip2(n4713), .op(n4716) );
  nand2_1 U5152 ( .ip1(n4714), .ip2(n4713), .op(n4715) );
  nand3_1 U5153 ( .ip1(n4717), .ip2(n4716), .ip3(n4715), .op(n4723) );
  nand2_1 U5154 ( .ip1(n4721), .ip2(n4723), .op(n4726) );
  nor2_1 U5155 ( .ip1(n4719), .ip2(n4718), .op(n4720) );
  nor3_1 U5156 ( .ip1(n4720), .ip2(n9540), .ip3(n13854), .op(n4722) );
  nand2_1 U5157 ( .ip1(n4721), .ip2(n4722), .op(n4725) );
  nand2_1 U5158 ( .ip1(n4723), .ip2(n4722), .op(n4724) );
  nand3_1 U5159 ( .ip1(n4726), .ip2(n4725), .ip3(n4724), .op(n4730) );
  nand2_1 U5160 ( .ip1(n4732), .ip2(n4730), .op(n4738) );
  fulladder U5161 ( .a(n4729), .b(n4728), .ci(n4727), .co(n4731), .s(n4721) );
  nand2_1 U5162 ( .ip1(n4730), .ip2(n4731), .op(n4737) );
  nand2_1 U5163 ( .ip1(n4732), .ip2(n4731), .op(n4736) );
  nand2_1 U5164 ( .ip1(n4734), .ip2(n4733), .op(n4735) );
  nand4_1 U5165 ( .ip1(n4738), .ip2(n4737), .ip3(n4736), .ip4(n4735), .op(
        n4742) );
  or2_1 U5166 ( .ip1(n4740), .ip2(n4739), .op(n4741) );
  nand3_1 U5167 ( .ip1(n4743), .ip2(n4742), .ip3(n4741), .op(n4744) );
  nand2_1 U5168 ( .ip1(n4745), .ip2(n4744), .op(n8986) );
  fulladder U5169 ( .a(n4748), .b(n4747), .ci(n4746), .co(n8985), .s(n4740) );
  inv_1 U5170 ( .ip(m1Inputs[146]), .op(n8721) );
  inv_1 U5171 ( .ip(m1Inputs[149]), .op(n14852) );
  nor4_1 U5172 ( .ip1(n10476), .ip2(n13082), .ip3(n8721), .ip4(n14852), .op(
        n4749) );
  inv_1 U5173 ( .ip(n4749), .op(n4754) );
  nand2_1 U5174 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[149]), .op(n4785) );
  or2_1 U5175 ( .ip1(n4785), .ip2(n4749), .op(n4752) );
  nand2_1 U5176 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[146]), .op(n4750) );
  or2_1 U5177 ( .ip1(n4750), .ip2(n4749), .op(n4751) );
  nand2_1 U5178 ( .ip1(n4752), .ip2(n4751), .op(n4815) );
  inv_1 U5179 ( .ip(m1Inputs[144]), .op(n8767) );
  nor2_1 U5180 ( .ip1(n8767), .ip2(n4624), .op(n4814) );
  nand2_1 U5181 ( .ip1(n4815), .ip2(n4814), .op(n4753) );
  nand2_1 U5182 ( .ip1(n4754), .ip2(n4753), .op(n4793) );
  nand2_1 U5183 ( .ip1(n4672), .ip2(m1Inputs[148]), .op(n4755) );
  inv_1 U5184 ( .ip(m1Inputs[148]), .op(n14785) );
  nor4_1 U5185 ( .ip1(n6745), .ip2(n9047), .ip3(n14785), .ip4(n14852), .op(
        n4810) );
  or2_1 U5186 ( .ip1(n4755), .ip2(n4810), .op(n4758) );
  nand2_1 U5187 ( .ip1(n12809), .ip2(m1Inputs[149]), .op(n4756) );
  or2_1 U5188 ( .ip1(n4756), .ip2(n4810), .op(n4757) );
  nand2_1 U5189 ( .ip1(n4758), .ip2(n4757), .op(n4792) );
  inv_1 U5190 ( .ip(m1Inputs[145]), .op(n8797) );
  nor2_1 U5191 ( .ip1(n8797), .ip2(n4624), .op(n4780) );
  inv_1 U5192 ( .ip(m1Inputs[150]), .op(n14841) );
  nor2_1 U5193 ( .ip1(n10476), .ip2(n14841), .op(n8325) );
  nor2_1 U5194 ( .ip1(n8767), .ip2(n14289), .op(n4779) );
  and3_1 U5195 ( .ip1(n10507), .ip2(m1Inputs[150]), .ip3(n4806), .op(n8363) );
  inv_1 U5196 ( .ip(m1Inputs[147]), .op(n8408) );
  nand2_1 U5197 ( .ip1(m1Inputs[146]), .ip2(\STAGE_1/weightReg [4]), .op(n4801) );
  nor3_1 U5198 ( .ip1(n8408), .ip2(n4801), .ip3(n4624), .op(n4770) );
  nor2_1 U5199 ( .ip1(n8408), .ip2(n14783), .op(n4781) );
  or2_1 U5200 ( .ip1(n14369), .ip2(n4781), .op(n4760) );
  or2_1 U5201 ( .ip1(m1Inputs[146]), .ip2(n4781), .op(n4759) );
  nand2_1 U5202 ( .ip1(n4760), .ip2(n4759), .op(n4769) );
  nand2_1 U5203 ( .ip1(m1Inputs[144]), .ip2(n14835), .op(n4771) );
  nor2_1 U5204 ( .ip1(n4769), .ip2(n4771), .op(n4761) );
  nor2_1 U5205 ( .ip1(n4770), .ip2(n4761), .op(n8332) );
  nand2_1 U5206 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[151]), .op(n8762) );
  nor2_1 U5207 ( .ip1(n10476), .ip2(n14785), .op(n4844) );
  and3_1 U5208 ( .ip1(n9733), .ip2(m1Inputs[151]), .ip3(n4844), .op(n4765) );
  or2_1 U5209 ( .ip1(n8762), .ip2(n4765), .op(n4764) );
  nand2_1 U5210 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[148]), .op(n4762) );
  or2_1 U5211 ( .ip1(n4762), .ip2(n4765), .op(n4763) );
  nand2_1 U5212 ( .ip1(n4764), .ip2(n4763), .op(n4777) );
  or2_1 U5213 ( .ip1(n4777), .ip2(n4765), .op(n4767) );
  nor2_1 U5214 ( .ip1(n6745), .ip2(n14852), .op(n4776) );
  or2_1 U5215 ( .ip1(n4776), .ip2(n4765), .op(n4766) );
  nand2_1 U5216 ( .ip1(n4767), .ip2(n4766), .op(n8331) );
  nand2_1 U5217 ( .ip1(m1Inputs[146]), .ip2(\STAGE_1/weightReg [6]), .op(n8330) );
  inv_1 U5218 ( .ip(n4768), .op(n8360) );
  nor2_1 U5219 ( .ip1(n4770), .ip2(n4769), .op(n4772) );
  xor2_1 U5220 ( .ip1(n4772), .ip2(n4771), .op(n4804) );
  nand4_1 U5221 ( .ip1(n4619), .ip2(\STAGE_1/weightReg [1]), .ip3(
        m1Inputs[147]), .ip4(m1Inputs[148]), .op(n4794) );
  nor2_1 U5222 ( .ip1(n13801), .ip2(n4794), .op(n4775) );
  nand2_1 U5223 ( .ip1(n4794), .ip2(m1Inputs[147]), .op(n4773) );
  mux2_1 U5224 ( .ip1(n4794), .ip2(n4773), .s(n9733), .op(n4800) );
  nor2_1 U5225 ( .ip1(n4801), .ip2(n4800), .op(n4774) );
  nor2_1 U5226 ( .ip1(n4775), .ip2(n4774), .op(n4803) );
  xnor2_1 U5227 ( .ip1(n4777), .ip2(n4776), .op(n4802) );
  inv_1 U5228 ( .ip(n4778), .op(n8359) );
  nor2_1 U5229 ( .ip1(n8797), .ip2(n14836), .op(n4811) );
  fulladder U5230 ( .a(n4780), .b(n8325), .ci(n4779), .co(n4809), .s(n4791) );
  nand2_1 U5231 ( .ip1(m1Inputs[147]), .ip2(\STAGE_1/weightReg [5]), .op(n4782) );
  and3_1 U5232 ( .ip1(m1Inputs[148]), .ip2(\STAGE_1/weightReg [5]), .ip3(n4781), .op(n8346) );
  or2_1 U5233 ( .ip1(n4782), .ip2(n8346), .op(n4784) );
  nand2_1 U5234 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[148]), .op(n8321) );
  or2_1 U5235 ( .ip1(n8321), .ip2(n8346), .op(n4783) );
  nand2_1 U5236 ( .ip1(n4784), .ip2(n4783), .op(n8345) );
  nor2_1 U5237 ( .ip1(n8797), .ip2(n14368), .op(n8347) );
  xor2_1 U5238 ( .ip1(n8345), .ip2(n8347), .op(n8357) );
  nand2_1 U5239 ( .ip1(n9733), .ip2(m1Inputs[149]), .op(n4786) );
  inv_1 U5240 ( .ip(m1Inputs[152]), .op(n14882) );
  nor3_1 U5241 ( .ip1(n13082), .ip2(n14882), .ip3(n4785), .op(n8341) );
  or2_1 U5242 ( .ip1(n4786), .ip2(n8341), .op(n4788) );
  nand2_1 U5243 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[152]), .op(n8708) );
  or2_1 U5244 ( .ip1(n8708), .ip2(n8341), .op(n4787) );
  nand2_1 U5245 ( .ip1(n4788), .ip2(n4787), .op(n8340) );
  nor2_1 U5246 ( .ip1(n8767), .ip2(n6504), .op(n8342) );
  xor2_1 U5247 ( .ip1(n8340), .ip2(n8342), .op(n8356) );
  nand2_1 U5248 ( .ip1(m1Inputs[150]), .ip2(n4619), .op(n4789) );
  nand2_1 U5249 ( .ip1(n10507), .ip2(m1Inputs[151]), .op(n8350) );
  nand2_1 U5250 ( .ip1(n4789), .ip2(n8350), .op(n4790) );
  nand4_1 U5251 ( .ip1(n4619), .ip2(\STAGE_1/weightReg [1]), .ip3(
        m1Inputs[151]), .ip4(m1Inputs[150]), .op(n8334) );
  nand2_1 U5252 ( .ip1(n4790), .ip2(n8334), .op(n8336) );
  buf_1 U5253 ( .ip(n14768), .op(n13498) );
  nand2_1 U5254 ( .ip1(column[144]), .ip2(n13498), .op(n8335) );
  xor2_1 U5255 ( .ip1(n8336), .ip2(n8335), .op(n8355) );
  fulladder U5256 ( .a(n4793), .b(n4792), .ci(n4791), .co(n4806), .s(n4862) );
  nand2_1 U5257 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[146]), .op(n4827) );
  nor3_1 U5258 ( .ip1(n10555), .ip2(n8408), .ip3(n4827), .op(n4838) );
  inv_1 U5259 ( .ip(n4794), .op(n4799) );
  nor2_1 U5260 ( .ip1(n6745), .ip2(n8408), .op(n4795) );
  or2_1 U5261 ( .ip1(m1Inputs[148]), .ip2(n4795), .op(n4797) );
  or2_1 U5262 ( .ip1(n13707), .ip2(n4795), .op(n4796) );
  nand2_1 U5263 ( .ip1(n4797), .ip2(n4796), .op(n4798) );
  nor2_1 U5264 ( .ip1(n4799), .ip2(n4798), .op(n4813) );
  nor2_1 U5265 ( .ip1(n8797), .ip2(n14783), .op(n4812) );
  xor2_1 U5266 ( .ip1(n4801), .ip2(n4800), .op(n4860) );
  fulladder U5267 ( .a(n4804), .b(n4803), .ci(n4802), .co(n4778), .s(n4805) );
  inv_1 U5268 ( .ip(n4805), .op(n4878) );
  nor2_1 U5269 ( .ip1(n13570), .ip2(n14841), .op(n4807) );
  nor2_1 U5270 ( .ip1(n4807), .ip2(n4806), .op(n4808) );
  nor2_1 U5271 ( .ip1(n8363), .ip2(n4808), .op(n4877) );
  fulladder U5272 ( .a(n4811), .b(n4810), .ci(n4809), .co(n8358), .s(n4876) );
  nand2_1 U5273 ( .ip1(n4870), .ip2(n4869), .op(n4875) );
  fulladder U5274 ( .a(n4838), .b(n4813), .ci(n4812), .co(n4861), .s(n4859) );
  nor2_1 U5275 ( .ip1(n13082), .ip2(n8797), .op(n4843) );
  nor2_1 U5276 ( .ip1(n8767), .ip2(n14783), .op(n4842) );
  xor2_1 U5277 ( .ip1(n4815), .ip2(n4814), .op(n4857) );
  nor2_1 U5278 ( .ip1(n10476), .ip2(n8408), .op(n4824) );
  nor4_1 U5279 ( .ip1(n6745), .ip2(n13570), .ip3(n8797), .ip4(n8767), .op(
        n4823) );
  nor2_1 U5280 ( .ip1(n4824), .ip2(n4823), .op(n4816) );
  nor3_1 U5281 ( .ip1(n4816), .ip2(n8797), .ip3(n6745), .op(n4845) );
  nor2_1 U5282 ( .ip1(n13570), .ip2(n8797), .op(n4817) );
  nor3_1 U5283 ( .ip1(n8721), .ip2(n6745), .ip3(n8767), .op(n4818) );
  or2_1 U5284 ( .ip1(n4817), .ip2(n4818), .op(n4821) );
  nand2_1 U5285 ( .ip1(n5056), .ip2(m1Inputs[144]), .op(n4819) );
  or2_1 U5286 ( .ip1(n4819), .ip2(n4818), .op(n4820) );
  nand2_1 U5287 ( .ip1(n4821), .ip2(n4820), .op(n4822) );
  not_ab_or_c_or_d U5288 ( .ip1(n8767), .ip2(n8721), .ip3(n4822), .ip4(n13646), 
        .op(n4831) );
  nand2_1 U5289 ( .ip1(n4619), .ip2(m1Inputs[145]), .op(n4826) );
  xnor2_1 U5290 ( .ip1(n4824), .ip2(n4823), .op(n4825) );
  xor2_1 U5291 ( .ip1(n4826), .ip2(n4825), .op(n4833) );
  nand2_1 U5292 ( .ip1(n4831), .ip2(n4833), .op(n4836) );
  inv_1 U5293 ( .ip(\STAGE_1/weightReg [3]), .op(n13487) );
  nor4_1 U5294 ( .ip1(n13570), .ip2(n13487), .ip3(n8767), .ip4(n8721), .op(
        n4853) );
  or2_1 U5295 ( .ip1(n4827), .ip2(n4853), .op(n4830) );
  buf_1 U5296 ( .ip(n9733), .op(n13614) );
  nand2_1 U5297 ( .ip1(n13614), .ip2(m1Inputs[144]), .op(n4828) );
  or2_1 U5298 ( .ip1(n4828), .ip2(n4853), .op(n4829) );
  nand2_1 U5299 ( .ip1(n4830), .ip2(n4829), .op(n4832) );
  nand2_1 U5300 ( .ip1(n4831), .ip2(n4832), .op(n4835) );
  nand2_1 U5301 ( .ip1(n4833), .ip2(n4832), .op(n4834) );
  nand3_1 U5302 ( .ip1(n4836), .ip2(n4835), .ip3(n4834), .op(n4847) );
  nand2_1 U5303 ( .ip1(n4845), .ip2(n4847), .op(n4850) );
  nand2_1 U5304 ( .ip1(n5056), .ip2(m1Inputs[146]), .op(n4837) );
  or2_1 U5305 ( .ip1(n4837), .ip2(n4838), .op(n4841) );
  nand2_1 U5306 ( .ip1(n13707), .ip2(m1Inputs[147]), .op(n4839) );
  or2_1 U5307 ( .ip1(n4839), .ip2(n4838), .op(n4840) );
  nand2_1 U5308 ( .ip1(n4841), .ip2(n4840), .op(n4852) );
  fulladder U5309 ( .a(n4844), .b(n4843), .ci(n4842), .co(n4858), .s(n4851) );
  nand2_1 U5310 ( .ip1(n4845), .ip2(n4846), .op(n4849) );
  nand2_1 U5311 ( .ip1(n4847), .ip2(n4846), .op(n4848) );
  nand3_1 U5312 ( .ip1(n4850), .ip2(n4849), .ip3(n4848), .op(n4854) );
  nand2_1 U5313 ( .ip1(n4856), .ip2(n4854), .op(n4866) );
  fulladder U5314 ( .a(n4853), .b(n4852), .ci(n4851), .co(n4855), .s(n4846) );
  nand2_1 U5315 ( .ip1(n4854), .ip2(n4855), .op(n4865) );
  nand2_1 U5316 ( .ip1(n4856), .ip2(n4855), .op(n4864) );
  fulladder U5317 ( .a(n4859), .b(n4858), .ci(n4857), .co(n4868), .s(n4856) );
  fulladder U5318 ( .a(n4862), .b(n4861), .ci(n4860), .co(n4870), .s(n4867) );
  nand2_1 U5319 ( .ip1(n4868), .ip2(n4867), .op(n4863) );
  nand4_1 U5320 ( .ip1(n4866), .ip2(n4865), .ip3(n4864), .ip4(n4863), .op(
        n4873) );
  or2_1 U5321 ( .ip1(n4868), .ip2(n4867), .op(n4872) );
  or2_1 U5322 ( .ip1(n4870), .ip2(n4869), .op(n4871) );
  nand3_1 U5323 ( .ip1(n4873), .ip2(n4872), .ip3(n4871), .op(n4874) );
  nand2_1 U5324 ( .ip1(n4875), .ip2(n4874), .op(n8365) );
  fulladder U5325 ( .a(n4878), .b(n4877), .ci(n4876), .co(n8364), .s(n4869) );
  inv_1 U5326 ( .ip(m1Inputs[114]), .op(n8099) );
  nor2_1 U5327 ( .ip1(n10476), .ip2(n8099), .op(n4955) );
  and3_1 U5328 ( .ip1(n12578), .ip2(n4955), .ip3(m1Inputs[117]), .op(n4879) );
  inv_1 U5329 ( .ip(n4879), .op(n4884) );
  nand2_1 U5330 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[117]), .op(n4916) );
  or2_1 U5331 ( .ip1(n4916), .ip2(n4879), .op(n4882) );
  nand2_1 U5332 ( .ip1(n9733), .ip2(m1Inputs[114]), .op(n4880) );
  or2_1 U5333 ( .ip1(n4880), .ip2(n4879), .op(n4881) );
  nand2_1 U5334 ( .ip1(n4882), .ip2(n4881), .op(n4980) );
  inv_1 U5335 ( .ip(m1Inputs[112]), .op(n8145) );
  nor2_1 U5336 ( .ip1(n8145), .ip2(n12746), .op(n4979) );
  nand2_1 U5337 ( .ip1(n4980), .ip2(n4979), .op(n4883) );
  nand2_1 U5338 ( .ip1(n4884), .ip2(n4883), .op(n4940) );
  nand2_1 U5339 ( .ip1(n4619), .ip2(m1Inputs[116]), .op(n4885) );
  inv_1 U5340 ( .ip(m1Inputs[116]), .op(n8166) );
  inv_1 U5341 ( .ip(m1Inputs[117]), .op(n14286) );
  nor4_1 U5342 ( .ip1(n6745), .ip2(n9047), .ip3(n8166), .ip4(n14286), .op(
        n4930) );
  or2_1 U5343 ( .ip1(n4885), .ip2(n4930), .op(n4888) );
  nand2_1 U5344 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[117]), .op(n4886) );
  or2_1 U5345 ( .ip1(n4886), .ip2(n4930), .op(n4887) );
  nand2_1 U5346 ( .ip1(n4888), .ip2(n4887), .op(n4939) );
  inv_1 U5347 ( .ip(m1Inputs[113]), .op(n8177) );
  nor2_1 U5348 ( .ip1(n8177), .ip2(n13835), .op(n4911) );
  inv_1 U5349 ( .ip(m1Inputs[118]), .op(n8172) );
  nor2_1 U5350 ( .ip1(n10476), .ip2(n8172), .op(n7706) );
  nor2_1 U5351 ( .ip1(n8145), .ip2(n14289), .op(n4910) );
  and3_1 U5352 ( .ip1(n10507), .ip2(m1Inputs[118]), .ip3(n4926), .op(n7744) );
  inv_1 U5353 ( .ip(m1Inputs[115]), .op(n7790) );
  inv_1 U5354 ( .ip(n14783), .op(n13637) );
  nand2_1 U5355 ( .ip1(m1Inputs[114]), .ip2(n13637), .op(n4942) );
  nor3_1 U5356 ( .ip1(n7790), .ip2(n4942), .ip3(n4624), .op(n4901) );
  nor2_1 U5357 ( .ip1(n7790), .ip2(n14783), .op(n4889) );
  or2_1 U5358 ( .ip1(n14369), .ip2(n4889), .op(n4891) );
  or2_1 U5359 ( .ip1(m1Inputs[114]), .ip2(n4889), .op(n4890) );
  nand2_1 U5360 ( .ip1(n4891), .ip2(n4890), .op(n4900) );
  nand2_1 U5361 ( .ip1(m1Inputs[112]), .ip2(n14835), .op(n4902) );
  nor2_1 U5362 ( .ip1(n4900), .ip2(n4902), .op(n4892) );
  nor2_1 U5363 ( .ip1(n4901), .ip2(n4892), .op(n7713) );
  nand2_1 U5364 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[119]), .op(n8140) );
  nor2_1 U5365 ( .ip1(n10476), .ip2(n8166), .op(n4978) );
  and3_1 U5366 ( .ip1(n12578), .ip2(m1Inputs[119]), .ip3(n4978), .op(n4896) );
  or2_1 U5367 ( .ip1(n8140), .ip2(n4896), .op(n4895) );
  nand2_1 U5368 ( .ip1(n13614), .ip2(m1Inputs[116]), .op(n4893) );
  or2_1 U5369 ( .ip1(n4893), .ip2(n4896), .op(n4894) );
  nand2_1 U5370 ( .ip1(n4895), .ip2(n4894), .op(n4908) );
  or2_1 U5371 ( .ip1(n4908), .ip2(n4896), .op(n4898) );
  inv_1 U5372 ( .ip(\STAGE_1/weightReg [2]), .op(n13854) );
  nor2_1 U5373 ( .ip1(n13854), .ip2(n14286), .op(n4907) );
  or2_1 U5374 ( .ip1(n4907), .ip2(n4896), .op(n4897) );
  nand2_1 U5375 ( .ip1(n4898), .ip2(n4897), .op(n7712) );
  nand2_1 U5376 ( .ip1(m1Inputs[114]), .ip2(n12981), .op(n7711) );
  inv_1 U5377 ( .ip(n4899), .op(n7741) );
  nor2_1 U5378 ( .ip1(n4901), .ip2(n4900), .op(n4903) );
  xor2_1 U5379 ( .ip1(n4903), .ip2(n4902), .op(n4924) );
  nand4_1 U5380 ( .ip1(\STAGE_1/weightReg [2]), .ip2(n10507), .ip3(
        m1Inputs[115]), .ip4(m1Inputs[116]), .op(n4932) );
  nor2_1 U5381 ( .ip1(n13801), .ip2(n4932), .op(n4906) );
  nand2_1 U5382 ( .ip1(n4932), .ip2(m1Inputs[115]), .op(n4904) );
  mux2_1 U5383 ( .ip1(n4932), .ip2(n4904), .s(n13614), .op(n4941) );
  nor2_1 U5384 ( .ip1(n4942), .ip2(n4941), .op(n4905) );
  nor2_1 U5385 ( .ip1(n4906), .ip2(n4905), .op(n4923) );
  xnor2_1 U5386 ( .ip1(n4908), .ip2(n4907), .op(n4922) );
  inv_1 U5387 ( .ip(n4909), .op(n7740) );
  nor2_1 U5388 ( .ip1(n8177), .ip2(n14836), .op(n4931) );
  fulladder U5389 ( .a(n4911), .b(n7706), .ci(n4910), .co(n4929), .s(n4938) );
  buf_1 U5390 ( .ip(\STAGE_1/weightReg [5]), .op(n14369) );
  nand2_1 U5391 ( .ip1(m1Inputs[115]), .ip2(n14369), .op(n4912) );
  nand2_1 U5392 ( .ip1(m1Inputs[116]), .ip2(n14369), .op(n7703) );
  nor3_1 U5393 ( .ip1(n7790), .ip2(n14783), .ip3(n7703), .op(n7727) );
  or2_1 U5394 ( .ip1(n4912), .ip2(n7727), .op(n4915) );
  nand2_1 U5395 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[116]), .op(n4913) );
  or2_1 U5396 ( .ip1(n4913), .ip2(n7727), .op(n4914) );
  nand2_1 U5397 ( .ip1(n4915), .ip2(n4914), .op(n7726) );
  nor2_1 U5398 ( .ip1(n8177), .ip2(n14368), .op(n7728) );
  xor2_1 U5399 ( .ip1(n7726), .ip2(n7728), .op(n7738) );
  nand2_1 U5400 ( .ip1(n9733), .ip2(m1Inputs[117]), .op(n4917) );
  inv_1 U5401 ( .ip(m1Inputs[120]), .op(n14418) );
  nor3_1 U5402 ( .ip1(n13082), .ip2(n14418), .ip3(n4916), .op(n7722) );
  or2_1 U5403 ( .ip1(n4917), .ip2(n7722), .op(n4919) );
  nand2_1 U5404 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[120]), .op(n8087) );
  or2_1 U5405 ( .ip1(n8087), .ip2(n7722), .op(n4918) );
  nand2_1 U5406 ( .ip1(n4919), .ip2(n4918), .op(n7721) );
  nor2_1 U5407 ( .ip1(n8145), .ip2(n6503), .op(n7723) );
  xor2_1 U5408 ( .ip1(n7721), .ip2(n7723), .op(n7737) );
  nand2_1 U5409 ( .ip1(m1Inputs[118]), .ip2(\STAGE_1/weightReg [2]), .op(n4920) );
  nand2_1 U5410 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[119]), .op(n7731) );
  nand2_1 U5411 ( .ip1(n4920), .ip2(n7731), .op(n4921) );
  nand4_1 U5412 ( .ip1(n4619), .ip2(n10507), .ip3(m1Inputs[119]), .ip4(
        m1Inputs[118]), .op(n7715) );
  nand2_1 U5413 ( .ip1(n4921), .ip2(n7715), .op(n7717) );
  nand2_1 U5414 ( .ip1(column[112]), .ip2(n13498), .op(n7716) );
  xor2_1 U5415 ( .ip1(n7717), .ip2(n7716), .op(n7736) );
  fulladder U5416 ( .a(n4924), .b(n4923), .ci(n4922), .co(n4909), .s(n4925) );
  inv_1 U5417 ( .ip(n4925), .op(n5011) );
  nor2_1 U5418 ( .ip1(n13570), .ip2(n8172), .op(n4927) );
  nor2_1 U5419 ( .ip1(n4927), .ip2(n4926), .op(n4928) );
  nor2_1 U5420 ( .ip1(n7744), .ip2(n4928), .op(n5010) );
  fulladder U5421 ( .a(n4931), .b(n4930), .ci(n4929), .co(n7739), .s(n5009) );
  nand2_1 U5422 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[114]), .op(n4950) );
  nor3_1 U5423 ( .ip1(n10555), .ip2(n7790), .ip3(n4950), .op(n4975) );
  inv_1 U5424 ( .ip(n4932), .op(n4937) );
  nor2_1 U5425 ( .ip1(n6745), .ip2(n7790), .op(n4933) );
  or2_1 U5426 ( .ip1(m1Inputs[116]), .ip2(n4933), .op(n4935) );
  or2_1 U5427 ( .ip1(n10507), .ip2(n4933), .op(n4934) );
  nand2_1 U5428 ( .ip1(n4935), .ip2(n4934), .op(n4936) );
  nor2_1 U5429 ( .ip1(n4937), .ip2(n4936), .op(n4974) );
  nor2_1 U5430 ( .ip1(n8177), .ip2(n14783), .op(n4973) );
  fulladder U5431 ( .a(n4940), .b(n4939), .ci(n4938), .co(n4926), .s(n4944) );
  xor2_1 U5432 ( .ip1(n4942), .ip2(n4941), .op(n4943) );
  nand2_1 U5433 ( .ip1(n5004), .ip2(n5003), .op(n5008) );
  fulladder U5434 ( .a(n4945), .b(n4944), .ci(n4943), .co(n5003), .s(n4998) );
  nor2_1 U5435 ( .ip1(n13487), .ip2(n8177), .op(n4977) );
  nor2_1 U5436 ( .ip1(n8145), .ip2(n14783), .op(n4976) );
  nor4_1 U5437 ( .ip1(n13570), .ip2(n13487), .ip3(n8145), .ip4(n8099), .op(
        n4971) );
  nor2_1 U5438 ( .ip1(n13570), .ip2(n7790), .op(n4946) );
  or2_1 U5439 ( .ip1(m1Inputs[114]), .ip2(n4946), .op(n4948) );
  or2_1 U5440 ( .ip1(n4619), .ip2(n4946), .op(n4947) );
  nand2_1 U5441 ( .ip1(n4948), .ip2(n4947), .op(n4949) );
  nor2_1 U5442 ( .ip1(n4975), .ip2(n4949), .op(n4970) );
  or2_1 U5443 ( .ip1(n4950), .ip2(n4971), .op(n4953) );
  nand2_1 U5444 ( .ip1(n12578), .ip2(m1Inputs[112]), .op(n4951) );
  or2_1 U5445 ( .ip1(n4951), .ip2(n4971), .op(n4952) );
  nand2_1 U5446 ( .ip1(n4953), .ip2(n4952), .op(n4964) );
  not_ab_or_c_or_d U5447 ( .ip1(n10507), .ip2(m1Inputs[112]), .ip3(n10555), 
        .ip4(n8177), .op(n4981) );
  nor2_1 U5448 ( .ip1(n10476), .ip2(n7790), .op(n4954) );
  xor2_1 U5449 ( .ip1(n4981), .ip2(n4954), .op(n4966) );
  nand2_1 U5450 ( .ip1(n4964), .ip2(n4966), .op(n4969) );
  nand2_1 U5451 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[113]), .op(n4959) );
  or2_1 U5452 ( .ip1(m1Inputs[112]), .ip2(n4955), .op(n4958) );
  inv_1 U5453 ( .ip(n5739), .op(n4956) );
  or2_1 U5454 ( .ip1(n4956), .ip2(n4955), .op(n4957) );
  nand2_1 U5455 ( .ip1(n4958), .ip2(n4957), .op(n4960) );
  or2_1 U5456 ( .ip1(n4959), .ip2(n4960), .op(n4963) );
  nand2_1 U5457 ( .ip1(n4672), .ip2(m1Inputs[112]), .op(n4961) );
  or2_1 U5458 ( .ip1(n4961), .ip2(n4960), .op(n4962) );
  nand2_1 U5459 ( .ip1(n4963), .ip2(n4962), .op(n4965) );
  nand2_1 U5460 ( .ip1(n4964), .ip2(n4965), .op(n4968) );
  nand2_1 U5461 ( .ip1(n4966), .ip2(n4965), .op(n4967) );
  nand3_1 U5462 ( .ip1(n4969), .ip2(n4968), .ip3(n4967), .op(n4987) );
  fulladder U5463 ( .a(n4972), .b(n4971), .ci(n4970), .co(n4994), .s(n4986) );
  fulladder U5464 ( .a(n4975), .b(n4974), .ci(n4973), .co(n4945), .s(n4992) );
  fulladder U5465 ( .a(n4978), .b(n4977), .ci(n4976), .co(n4991), .s(n4972) );
  xor2_1 U5466 ( .ip1(n4980), .ip2(n4979), .op(n4990) );
  and2_1 U5467 ( .ip1(n4994), .ip2(n4993), .op(n4985) );
  nor3_1 U5468 ( .ip1(n4986), .ip2(n4987), .ip3(n4985), .op(n4989) );
  nand4_1 U5469 ( .ip1(n5056), .ip2(\STAGE_1/weightReg [1]), .ip3(
        m1Inputs[113]), .ip4(m1Inputs[112]), .op(n4983) );
  nand3_1 U5470 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n4981), .ip3(
        m1Inputs[115]), .op(n4982) );
  nand2_1 U5471 ( .ip1(n4983), .ip2(n4982), .op(n4984) );
  not_ab_or_c_or_d U5472 ( .ip1(n4987), .ip2(n4986), .ip3(n4985), .ip4(n4984), 
        .op(n4988) );
  or2_1 U5473 ( .ip1(n4989), .ip2(n4988), .op(n4997) );
  fulladder U5474 ( .a(n4992), .b(n4991), .ci(n4990), .co(n5000), .s(n4993) );
  nor2_1 U5475 ( .ip1(n5000), .ip2(n4998), .op(n4996) );
  nor2_1 U5476 ( .ip1(n4994), .ip2(n4993), .op(n4995) );
  nor3_1 U5477 ( .ip1(n4997), .ip2(n4996), .ip3(n4995), .op(n4999) );
  or2_1 U5478 ( .ip1(n4998), .ip2(n4999), .op(n5002) );
  or2_1 U5479 ( .ip1(n5000), .ip2(n4999), .op(n5001) );
  nand2_1 U5480 ( .ip1(n5002), .ip2(n5001), .op(n5006) );
  nor2_1 U5481 ( .ip1(n5004), .ip2(n5003), .op(n5005) );
  or2_1 U5482 ( .ip1(n5006), .ip2(n5005), .op(n5007) );
  nand2_1 U5483 ( .ip1(n5008), .ip2(n5007), .op(n7746) );
  fulladder U5484 ( .a(n5011), .b(n5010), .ci(n5009), .co(n7745), .s(n5004) );
  inv_1 U5485 ( .ip(m1Inputs[98]), .op(n7486) );
  inv_1 U5486 ( .ip(m1Inputs[101]), .op(n7326) );
  nor4_1 U5487 ( .ip1(n13646), .ip2(n13082), .ip3(n7486), .ip4(n7326), .op(
        n5012) );
  inv_1 U5488 ( .ip(n5012), .op(n5017) );
  nand2_1 U5489 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[101]), .op(n5050) );
  or2_1 U5490 ( .ip1(n5050), .ip2(n5012), .op(n5015) );
  nand2_1 U5491 ( .ip1(n13614), .ip2(m1Inputs[98]), .op(n5013) );
  or2_1 U5492 ( .ip1(n5013), .ip2(n5012), .op(n5014) );
  nand2_1 U5493 ( .ip1(n5015), .ip2(n5014), .op(n5115) );
  inv_1 U5494 ( .ip(m1Inputs[96]), .op(n7532) );
  nor2_1 U5495 ( .ip1(n7532), .ip2(n4624), .op(n5114) );
  nand2_1 U5496 ( .ip1(n5115), .ip2(n5114), .op(n5016) );
  nand2_1 U5497 ( .ip1(n5017), .ip2(n5016), .op(n5065) );
  nand2_1 U5498 ( .ip1(n4619), .ip2(m1Inputs[100]), .op(n5018) );
  inv_1 U5499 ( .ip(m1Inputs[100]), .op(n7553) );
  nor4_1 U5500 ( .ip1(n6745), .ip2(n13570), .ip3(n7553), .ip4(n7326), .op(
        n5076) );
  or2_1 U5501 ( .ip1(n5018), .ip2(n5076), .op(n5021) );
  nand2_1 U5502 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[101]), .op(n5019) );
  or2_1 U5503 ( .ip1(n5019), .ip2(n5076), .op(n5020) );
  nand2_1 U5504 ( .ip1(n5021), .ip2(n5020), .op(n5064) );
  inv_1 U5505 ( .ip(m1Inputs[97]), .op(n7564) );
  nor2_1 U5506 ( .ip1(n7564), .ip2(n12746), .op(n5044) );
  inv_1 U5507 ( .ip(m1Inputs[102]), .op(n7559) );
  nor2_1 U5508 ( .ip1(n10476), .ip2(n7559), .op(n6938) );
  nor2_1 U5509 ( .ip1(n7532), .ip2(n14836), .op(n5043) );
  and3_1 U5510 ( .ip1(n10507), .ip2(m1Inputs[102]), .ip3(n5072), .op(n6976) );
  nand2_1 U5511 ( .ip1(m1Inputs[99]), .ip2(n13637), .op(n5045) );
  inv_1 U5512 ( .ip(m1Inputs[99]), .op(n7184) );
  nand2_1 U5513 ( .ip1(m1Inputs[98]), .ip2(n13637), .op(n5067) );
  nor3_1 U5514 ( .ip1(n7184), .ip2(n5067), .ip3(n12746), .op(n5025) );
  or2_1 U5515 ( .ip1(n5045), .ip2(n5025), .op(n5024) );
  nand2_1 U5516 ( .ip1(m1Inputs[98]), .ip2(n14369), .op(n5022) );
  or2_1 U5517 ( .ip1(n5022), .ip2(n5025), .op(n5023) );
  nand2_1 U5518 ( .ip1(n5024), .ip2(n5023), .op(n5036) );
  or2_1 U5519 ( .ip1(n5036), .ip2(n5025), .op(n5027) );
  nor2_1 U5520 ( .ip1(n7532), .ip2(n14384), .op(n5035) );
  or2_1 U5521 ( .ip1(n5035), .ip2(n5025), .op(n5026) );
  nand2_1 U5522 ( .ip1(n5027), .ip2(n5026), .op(n6945) );
  nand2_1 U5523 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[103]), .op(n7527) );
  nor2_1 U5524 ( .ip1(n10476), .ip2(n7553), .op(n5113) );
  and3_1 U5525 ( .ip1(n12578), .ip2(m1Inputs[103]), .ip3(n5113), .op(n5031) );
  or2_1 U5526 ( .ip1(n7527), .ip2(n5031), .op(n5030) );
  nand2_1 U5527 ( .ip1(n13614), .ip2(m1Inputs[100]), .op(n5028) );
  or2_1 U5528 ( .ip1(n5028), .ip2(n5031), .op(n5029) );
  nand2_1 U5529 ( .ip1(n5030), .ip2(n5029), .op(n5041) );
  or2_1 U5530 ( .ip1(n5041), .ip2(n5031), .op(n5033) );
  nor2_1 U5531 ( .ip1(n13854), .ip2(n7326), .op(n5040) );
  or2_1 U5532 ( .ip1(n5040), .ip2(n5031), .op(n5032) );
  nand2_1 U5533 ( .ip1(n5033), .ip2(n5032), .op(n6944) );
  nand2_1 U5534 ( .ip1(m1Inputs[98]), .ip2(n12981), .op(n6943) );
  inv_1 U5535 ( .ip(n5034), .op(n6973) );
  xnor2_1 U5536 ( .ip1(n5036), .ip2(n5035), .op(n5070) );
  nand4_1 U5537 ( .ip1(n4672), .ip2(\STAGE_1/weightReg [1]), .ip3(m1Inputs[99]), .ip4(m1Inputs[100]), .op(n5057) );
  nor2_1 U5538 ( .ip1(n13801), .ip2(n5057), .op(n5039) );
  nand2_1 U5539 ( .ip1(n5057), .ip2(m1Inputs[99]), .op(n5037) );
  mux2_1 U5540 ( .ip1(n5057), .ip2(n5037), .s(n13614), .op(n5066) );
  nor2_1 U5541 ( .ip1(n5067), .ip2(n5066), .op(n5038) );
  nor2_1 U5542 ( .ip1(n5039), .ip2(n5038), .op(n5069) );
  xnor2_1 U5543 ( .ip1(n5041), .ip2(n5040), .op(n5068) );
  inv_1 U5544 ( .ip(n5042), .op(n6972) );
  nor2_1 U5545 ( .ip1(n7564), .ip2(n14836), .op(n5077) );
  fulladder U5546 ( .a(n5044), .b(n6938), .ci(n5043), .co(n5075), .s(n5063) );
  nand2_1 U5547 ( .ip1(m1Inputs[99]), .ip2(n14369), .op(n5046) );
  nand2_1 U5548 ( .ip1(m1Inputs[100]), .ip2(\STAGE_1/weightReg [5]), .op(n6935) );
  nor2_1 U5549 ( .ip1(n5045), .ip2(n6935), .op(n6959) );
  or2_1 U5550 ( .ip1(n5046), .ip2(n6959), .op(n5049) );
  nand2_1 U5551 ( .ip1(n13637), .ip2(m1Inputs[100]), .op(n5047) );
  or2_1 U5552 ( .ip1(n5047), .ip2(n6959), .op(n5048) );
  nand2_1 U5553 ( .ip1(n5049), .ip2(n5048), .op(n6958) );
  nor2_1 U5554 ( .ip1(n7564), .ip2(n14368), .op(n6960) );
  xor2_1 U5555 ( .ip1(n6958), .ip2(n6960), .op(n6970) );
  nand2_1 U5556 ( .ip1(n13614), .ip2(m1Inputs[101]), .op(n5051) );
  inv_1 U5557 ( .ip(m1Inputs[104]), .op(n14169) );
  nor3_1 U5558 ( .ip1(n13082), .ip2(n14169), .ip3(n5050), .op(n6954) );
  or2_1 U5559 ( .ip1(n5051), .ip2(n6954), .op(n5053) );
  nand2_1 U5560 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[104]), .op(n7473) );
  or2_1 U5561 ( .ip1(n7473), .ip2(n6954), .op(n5052) );
  nand2_1 U5562 ( .ip1(n5053), .ip2(n5052), .op(n6953) );
  nor2_1 U5563 ( .ip1(n7532), .ip2(n6503), .op(n6955) );
  xor2_1 U5564 ( .ip1(n6953), .ip2(n6955), .op(n6969) );
  nand2_1 U5565 ( .ip1(m1Inputs[102]), .ip2(n4672), .op(n5054) );
  nand2_1 U5566 ( .ip1(n10507), .ip2(m1Inputs[103]), .op(n6963) );
  nand2_1 U5567 ( .ip1(n5054), .ip2(n6963), .op(n5055) );
  nand4_1 U5568 ( .ip1(\STAGE_1/weightReg [2]), .ip2(n10507), .ip3(
        m1Inputs[103]), .ip4(m1Inputs[102]), .op(n6947) );
  nand2_1 U5569 ( .ip1(n5055), .ip2(n6947), .op(n6949) );
  nand2_1 U5570 ( .ip1(column[96]), .ip2(n13498), .op(n6948) );
  xor2_1 U5571 ( .ip1(n6949), .ip2(n6948), .op(n6968) );
  buf_1 U5572 ( .ip(\STAGE_1/weightReg [2]), .op(n5056) );
  inv_1 U5573 ( .ip(n5056), .op(n13709) );
  nand2_1 U5574 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[98]), .op(n5088)
         );
  nor3_1 U5575 ( .ip1(n13709), .ip2(n7184), .ip3(n5088), .op(n5110) );
  inv_1 U5576 ( .ip(n5057), .op(n5062) );
  nor2_1 U5577 ( .ip1(n13854), .ip2(n7184), .op(n5058) );
  or2_1 U5578 ( .ip1(m1Inputs[100]), .ip2(n5058), .op(n5060) );
  or2_1 U5579 ( .ip1(n10507), .ip2(n5058), .op(n5059) );
  nand2_1 U5580 ( .ip1(n5060), .ip2(n5059), .op(n5061) );
  nor2_1 U5581 ( .ip1(n5062), .ip2(n5061), .op(n5109) );
  nor2_1 U5582 ( .ip1(n7564), .ip2(n14783), .op(n5108) );
  fulladder U5583 ( .a(n5065), .b(n5064), .ci(n5063), .co(n5072), .s(n5128) );
  xor2_1 U5584 ( .ip1(n5067), .ip2(n5066), .op(n5127) );
  fulladder U5585 ( .a(n5070), .b(n5069), .ci(n5068), .co(n5042), .s(n5071) );
  inv_1 U5586 ( .ip(n5071), .op(n5142) );
  nor2_1 U5587 ( .ip1(n13570), .ip2(n7559), .op(n5073) );
  nor2_1 U5588 ( .ip1(n5073), .ip2(n5072), .op(n5074) );
  nor2_1 U5589 ( .ip1(n6976), .ip2(n5074), .op(n5141) );
  fulladder U5590 ( .a(n5077), .b(n5076), .ci(n5075), .co(n6971), .s(n5140) );
  nand2_1 U5591 ( .ip1(n5131), .ip2(n5130), .op(n5139) );
  nand4_1 U5592 ( .ip1(n4619), .ip2(n10507), .ip3(m1Inputs[97]), .ip4(
        m1Inputs[96]), .op(n5079) );
  not_ab_or_c_or_d U5593 ( .ip1(n10507), .ip2(m1Inputs[96]), .ip3(n10555), 
        .ip4(n7564), .op(n5087) );
  nand3_1 U5594 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n5087), .ip3(m1Inputs[99]), .op(n5078) );
  nand2_1 U5595 ( .ip1(n5079), .ip2(n5078), .op(n5104) );
  nor2_1 U5596 ( .ip1(n13570), .ip2(n7564), .op(n5080) );
  nor3_1 U5597 ( .ip1(n7486), .ip2(n6745), .ip3(n7532), .op(n5081) );
  or2_1 U5598 ( .ip1(n5080), .ip2(n5081), .op(n5084) );
  nand2_1 U5599 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[96]), .op(n5082)
         );
  or2_1 U5600 ( .ip1(n5082), .ip2(n5081), .op(n5083) );
  nand2_1 U5601 ( .ip1(n5084), .ip2(n5083), .op(n5085) );
  not_ab_or_c_or_d U5602 ( .ip1(n7532), .ip2(n7486), .ip3(n5085), .ip4(n10476), 
        .op(n5092) );
  nor2_1 U5603 ( .ip1(n10476), .ip2(n7184), .op(n5086) );
  xor2_1 U5604 ( .ip1(n5087), .ip2(n5086), .op(n5094) );
  nand2_1 U5605 ( .ip1(n5092), .ip2(n5094), .op(n5097) );
  nor4_1 U5606 ( .ip1(n9047), .ip2(n13082), .ip3(n7532), .ip4(n7486), .op(
        n5107) );
  or2_1 U5607 ( .ip1(n5088), .ip2(n5107), .op(n5091) );
  nand2_1 U5608 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[96]), .op(n5089)
         );
  or2_1 U5609 ( .ip1(n5089), .ip2(n5107), .op(n5090) );
  nand2_1 U5610 ( .ip1(n5091), .ip2(n5090), .op(n5093) );
  nand2_1 U5611 ( .ip1(n5092), .ip2(n5093), .op(n5096) );
  nand2_1 U5612 ( .ip1(n5094), .ip2(n5093), .op(n5095) );
  nand3_1 U5613 ( .ip1(n5097), .ip2(n5096), .ip3(n5095), .op(n5102) );
  nand2_1 U5614 ( .ip1(n5104), .ip2(n5102), .op(n5119) );
  nand2_1 U5615 ( .ip1(n4619), .ip2(m1Inputs[98]), .op(n5098) );
  or2_1 U5616 ( .ip1(n5098), .ip2(n5110), .op(n5101) );
  nand2_1 U5617 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[99]), .op(n5099)
         );
  or2_1 U5618 ( .ip1(n5099), .ip2(n5110), .op(n5100) );
  nand2_1 U5619 ( .ip1(n5101), .ip2(n5100), .op(n5106) );
  nor2_1 U5620 ( .ip1(n13487), .ip2(n7564), .op(n5112) );
  nor2_1 U5621 ( .ip1(n7532), .ip2(n14783), .op(n5111) );
  nand2_1 U5622 ( .ip1(n5102), .ip2(n5103), .op(n5118) );
  nand2_1 U5623 ( .ip1(n5104), .ip2(n5103), .op(n5117) );
  fulladder U5624 ( .a(n5107), .b(n5106), .ci(n5105), .co(n5121), .s(n5103) );
  fulladder U5625 ( .a(n5110), .b(n5109), .ci(n5108), .co(n5129), .s(n5126) );
  fulladder U5626 ( .a(n5113), .b(n5112), .ci(n5111), .co(n5125), .s(n5105) );
  xor2_1 U5627 ( .ip1(n5115), .ip2(n5114), .op(n5124) );
  nand2_1 U5628 ( .ip1(n5121), .ip2(n5120), .op(n5116) );
  nand4_1 U5629 ( .ip1(n5119), .ip2(n5118), .ip3(n5117), .ip4(n5116), .op(
        n5123) );
  or2_1 U5630 ( .ip1(n5121), .ip2(n5120), .op(n5122) );
  nand2_1 U5631 ( .ip1(n5123), .ip2(n5122), .op(n5137) );
  fulladder U5632 ( .a(n5126), .b(n5125), .ci(n5124), .co(n5133), .s(n5120) );
  fulladder U5633 ( .a(n5129), .b(n5128), .ci(n5127), .co(n5131), .s(n5132) );
  nand2_1 U5634 ( .ip1(n5133), .ip2(n5132), .op(n5136) );
  nor2_1 U5635 ( .ip1(n5131), .ip2(n5130), .op(n5135) );
  nor2_1 U5636 ( .ip1(n5133), .ip2(n5132), .op(n5134) );
  ab_or_c_or_d U5637 ( .ip1(n5137), .ip2(n5136), .ip3(n5135), .ip4(n5134), 
        .op(n5138) );
  nand2_1 U5638 ( .ip1(n5139), .ip2(n5138), .op(n6978) );
  fulladder U5639 ( .a(n5142), .b(n5141), .ci(n5140), .co(n6977), .s(n5130) );
  inv_1 U5640 ( .ip(m1Inputs[53]), .op(n12255) );
  nor2_1 U5641 ( .ip1(n13646), .ip2(n12255), .op(n5212) );
  inv_1 U5642 ( .ip(m1Inputs[50]), .op(n12032) );
  nor2_1 U5643 ( .ip1(n13082), .ip2(n12032), .op(n5217) );
  inv_1 U5644 ( .ip(m1Inputs[48]), .op(n11858) );
  nor2_1 U5645 ( .ip1(n11858), .ip2(n4624), .op(n11160) );
  nand2_1 U5646 ( .ip1(n4672), .ip2(m1Inputs[52]), .op(n5143) );
  inv_1 U5647 ( .ip(m1Inputs[52]), .op(n12066) );
  nor4_1 U5648 ( .ip1(n6745), .ip2(n9047), .ip3(n12066), .ip4(n12255), .op(
        n5197) );
  or2_1 U5649 ( .ip1(n5143), .ip2(n5197), .op(n5146) );
  buf_1 U5650 ( .ip(n13707), .op(n12809) );
  nand2_1 U5651 ( .ip1(n12809), .ip2(m1Inputs[53]), .op(n5144) );
  or2_1 U5652 ( .ip1(n5144), .ip2(n5197), .op(n5145) );
  nand2_1 U5653 ( .ip1(n5146), .ip2(n5145), .op(n5206) );
  inv_1 U5654 ( .ip(m1Inputs[49]), .op(n12126) );
  inv_1 U5655 ( .ip(\STAGE_1/weightReg [5]), .op(n12746) );
  nor2_1 U5656 ( .ip1(n12126), .ip2(n12746), .op(n5168) );
  inv_1 U5657 ( .ip(m1Inputs[54]), .op(n12063) );
  nor2_1 U5658 ( .ip1(n13646), .ip2(n12063), .op(n6733) );
  nor2_1 U5659 ( .ip1(n11858), .ip2(n14289), .op(n11225) );
  and3_1 U5660 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[54]), .ip3(n5193), 
        .op(n6763) );
  nand2_1 U5661 ( .ip1(m1Inputs[51]), .ip2(\STAGE_1/weightReg [4]), .op(n5169)
         );
  inv_1 U5662 ( .ip(m1Inputs[51]), .op(n12138) );
  nand2_1 U5663 ( .ip1(m1Inputs[50]), .ip2(\STAGE_1/weightReg [4]), .op(n5209)
         );
  nor3_1 U5664 ( .ip1(n12138), .ip2(n5209), .ip3(n4624), .op(n5150) );
  or2_1 U5665 ( .ip1(n5169), .ip2(n5150), .op(n5149) );
  nand2_1 U5666 ( .ip1(m1Inputs[50]), .ip2(n12699), .op(n5147) );
  or2_1 U5667 ( .ip1(n5147), .ip2(n5150), .op(n5148) );
  nand2_1 U5668 ( .ip1(n5149), .ip2(n5148), .op(n5158) );
  or2_1 U5669 ( .ip1(n5158), .ip2(n5150), .op(n5152) );
  nor2_1 U5670 ( .ip1(n11858), .ip2(n12156), .op(n11792) );
  or2_1 U5671 ( .ip1(n11792), .ip2(n5150), .op(n5151) );
  nand2_1 U5672 ( .ip1(n5152), .ip2(n5151), .op(n6740) );
  nand2_1 U5673 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[55]), .op(n6788)
         );
  nor3_1 U5674 ( .ip1(n10476), .ip2(n12066), .ip3(n6788), .op(n5164) );
  inv_1 U5675 ( .ip(m1Inputs[55]), .op(n12155) );
  nor2_1 U5676 ( .ip1(n13646), .ip2(n12155), .op(n5153) );
  or2_1 U5677 ( .ip1(m1Inputs[52]), .ip2(n5153), .op(n5155) );
  or2_1 U5678 ( .ip1(n9733), .ip2(n5153), .op(n5154) );
  nand2_1 U5679 ( .ip1(n5155), .ip2(n5154), .op(n5163) );
  nand2_1 U5680 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[53]), .op(n5165)
         );
  nor2_1 U5681 ( .ip1(n5163), .ip2(n5165), .op(n5156) );
  nor2_1 U5682 ( .ip1(n5164), .ip2(n5156), .op(n6739) );
  inv_1 U5683 ( .ip(n14289), .op(n12981) );
  nand2_1 U5684 ( .ip1(m1Inputs[50]), .ip2(n12981), .op(n6738) );
  inv_1 U5685 ( .ip(n5157), .op(n6760) );
  inv_1 U5686 ( .ip(n11792), .op(n5159) );
  mux2_1 U5687 ( .ip1(n5159), .ip2(n11792), .s(n5158), .op(n5191) );
  nand4_1 U5688 ( .ip1(\STAGE_1/weightReg [2]), .ip2(\STAGE_1/weightReg [1]), 
        .ip3(m1Inputs[51]), .ip4(m1Inputs[52]), .op(n5199) );
  nor2_1 U5689 ( .ip1(n13487), .ip2(n5199), .op(n5162) );
  nand2_1 U5690 ( .ip1(n5199), .ip2(m1Inputs[51]), .op(n5160) );
  mux2_1 U5691 ( .ip1(n5199), .ip2(n5160), .s(n9733), .op(n5208) );
  nor2_1 U5692 ( .ip1(n5209), .ip2(n5208), .op(n5161) );
  nor2_1 U5693 ( .ip1(n5162), .ip2(n5161), .op(n5190) );
  nor2_1 U5694 ( .ip1(n5164), .ip2(n5163), .op(n5166) );
  xor2_1 U5695 ( .ip1(n5166), .ip2(n5165), .op(n5189) );
  inv_1 U5696 ( .ip(n5167), .op(n6759) );
  nor2_1 U5697 ( .ip1(n12126), .ip2(n14836), .op(n5198) );
  fulladder U5698 ( .a(n5168), .b(n6733), .ci(n11225), .co(n5196), .s(n5205)
         );
  inv_1 U5699 ( .ip(\STAGE_1/weightReg [5]), .op(n13835) );
  nor3_1 U5700 ( .ip1(n12066), .ip2(n13835), .ip3(n5169), .op(n6753) );
  inv_1 U5701 ( .ip(n6753), .op(n5172) );
  nand2_1 U5702 ( .ip1(m1Inputs[51]), .ip2(n12699), .op(n5170) );
  nand2_1 U5703 ( .ip1(n13637), .ip2(m1Inputs[52]), .op(n6729) );
  nand2_1 U5704 ( .ip1(n5170), .ip2(n6729), .op(n5171) );
  nand2_1 U5705 ( .ip1(n5172), .ip2(n5171), .op(n5173) );
  nor3_1 U5706 ( .ip1(n12126), .ip2(n14384), .ip3(n5173), .op(n6752) );
  or2_1 U5707 ( .ip1(n5173), .ip2(n6752), .op(n5176) );
  nand2_1 U5708 ( .ip1(m1Inputs[49]), .ip2(n4627), .op(n5174) );
  or2_1 U5709 ( .ip1(n5174), .ip2(n6752), .op(n5175) );
  nand2_1 U5710 ( .ip1(n5176), .ip2(n5175), .op(n6757) );
  inv_1 U5711 ( .ip(n6503), .op(n14975) );
  nand2_1 U5712 ( .ip1(m1Inputs[48]), .ip2(n14975), .op(n11830) );
  nand2_1 U5713 ( .ip1(m1Inputs[53]), .ip2(n12578), .op(n5177) );
  nand2_1 U5714 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[56]), .op(n6835)
         );
  nand2_1 U5715 ( .ip1(n5177), .ip2(n6835), .op(n5178) );
  nand3_1 U5716 ( .ip1(n13614), .ip2(m1Inputs[56]), .ip3(n5212), .op(n6749) );
  nand2_1 U5717 ( .ip1(n5178), .ip2(n6749), .op(n5179) );
  nor3_1 U5718 ( .ip1(n11858), .ip2(n6503), .ip3(n5179), .op(n6750) );
  or2_1 U5719 ( .ip1(n11830), .ip2(n6750), .op(n5181) );
  or2_1 U5720 ( .ip1(n5179), .ip2(n6750), .op(n5180) );
  nand2_1 U5721 ( .ip1(n5181), .ip2(n5180), .op(n6756) );
  nand2_1 U5722 ( .ip1(n12809), .ip2(m1Inputs[55]), .op(n5182) );
  nand4_1 U5723 ( .ip1(\STAGE_1/weightReg [2]), .ip2(n10507), .ip3(
        m1Inputs[55]), .ip4(m1Inputs[54]), .op(n6744) );
  inv_1 U5724 ( .ip(n6744), .op(n5183) );
  or2_1 U5725 ( .ip1(n5182), .ip2(n5183), .op(n5186) );
  nand2_1 U5726 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[54]), .op(n5184)
         );
  or2_1 U5727 ( .ip1(n5184), .ip2(n5183), .op(n5185) );
  nand2_1 U5728 ( .ip1(n5186), .ip2(n5185), .op(n6742) );
  inv_1 U5729 ( .ip(n6742), .op(n5188) );
  nand2_1 U5730 ( .ip1(column[48]), .ip2(n14768), .op(n5187) );
  mux2_1 U5731 ( .ip1(n5188), .ip2(n6742), .s(n5187), .op(n6755) );
  fulladder U5732 ( .a(n5191), .b(n5190), .ci(n5189), .co(n5167), .s(n5192) );
  inv_1 U5733 ( .ip(n5192), .op(n5272) );
  nor2_1 U5734 ( .ip1(n9047), .ip2(n12063), .op(n5194) );
  nor2_1 U5735 ( .ip1(n5194), .ip2(n5193), .op(n5195) );
  nor2_1 U5736 ( .ip1(n6763), .ip2(n5195), .op(n5271) );
  fulladder U5737 ( .a(n5198), .b(n5197), .ci(n5196), .co(n6758), .s(n5270) );
  nor2_1 U5738 ( .ip1(n13570), .ip2(n12032), .op(n5237) );
  and3_1 U5739 ( .ip1(n4672), .ip2(n5237), .ip3(m1Inputs[51]), .op(n5219) );
  inv_1 U5740 ( .ip(n5199), .op(n5204) );
  nor2_1 U5741 ( .ip1(n13854), .ip2(n12138), .op(n5200) );
  or2_1 U5742 ( .ip1(m1Inputs[52]), .ip2(n5200), .op(n5202) );
  or2_1 U5743 ( .ip1(n10507), .ip2(n5200), .op(n5201) );
  nand2_1 U5744 ( .ip1(n5202), .ip2(n5201), .op(n5203) );
  nor2_1 U5745 ( .ip1(n5204), .ip2(n5203), .op(n5211) );
  nor2_1 U5746 ( .ip1(n12126), .ip2(n14783), .op(n5210) );
  fulladder U5747 ( .a(n5207), .b(n5206), .ci(n5205), .co(n5193), .s(n5215) );
  xor2_1 U5748 ( .ip1(n5209), .ip2(n5208), .op(n5214) );
  nand2_1 U5749 ( .ip1(n5261), .ip2(n5260), .op(n5269) );
  fulladder U5750 ( .a(n5219), .b(n5211), .ci(n5210), .co(n5216), .s(n5227) );
  nor2_1 U5751 ( .ip1(n13646), .ip2(n12066), .op(n5224) );
  nor2_1 U5752 ( .ip1(n13082), .ip2(n12126), .op(n5223) );
  nor2_1 U5753 ( .ip1(n11858), .ip2(n14783), .op(n11207) );
  fulladder U5754 ( .a(n5212), .b(n5217), .ci(n11160), .co(n5207), .s(n5225)
         );
  inv_1 U5755 ( .ip(n5213), .op(n5267) );
  fulladder U5756 ( .a(n5216), .b(n5215), .ci(n5214), .co(n5260), .s(n5263) );
  nor2_1 U5757 ( .ip1(n9047), .ip2(n11858), .op(n11421) );
  and2_1 U5758 ( .ip1(n5217), .ip2(n11421), .op(n5247) );
  nand2_1 U5759 ( .ip1(n12809), .ip2(m1Inputs[51]), .op(n5218) );
  or2_1 U5760 ( .ip1(n5218), .ip2(n5219), .op(n5222) );
  nand2_1 U5761 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[50]), .op(n5220)
         );
  or2_1 U5762 ( .ip1(n5220), .ip2(n5219), .op(n5221) );
  nand2_1 U5763 ( .ip1(n5222), .ip2(n5221), .op(n5246) );
  fulladder U5764 ( .a(n5224), .b(n5223), .ci(n11207), .co(n5226), .s(n5245)
         );
  fulladder U5765 ( .a(n5227), .b(n5226), .ci(n5225), .co(n5213), .s(n5256) );
  nand2_1 U5766 ( .ip1(n5254), .ip2(n5256), .op(n5259) );
  inv_1 U5767 ( .ip(n11421), .op(n5228) );
  nand2_1 U5768 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[51]), .op(n5236)
         );
  not_ab_or_c_or_d U5769 ( .ip1(n5228), .ip2(n5236), .ip3(n12126), .ip4(n6745), 
        .op(n5248) );
  nor2_1 U5770 ( .ip1(n6745), .ip2(n11858), .op(n11386) );
  or2_1 U5771 ( .ip1(m1Inputs[49]), .ip2(n11386), .op(n5230) );
  or2_1 U5772 ( .ip1(n13707), .ip2(n11386), .op(n5229) );
  nand2_1 U5773 ( .ip1(n5230), .ip2(n5229), .op(n5234) );
  nor2_1 U5774 ( .ip1(n5739), .ip2(n11858), .op(n5231) );
  or2_1 U5775 ( .ip1(m1Inputs[50]), .ip2(n5231), .op(n5232) );
  nand2_1 U5776 ( .ip1(n5232), .ip2(n13803), .op(n5233) );
  nor2_1 U5777 ( .ip1(n5234), .ip2(n5233), .op(n5239) );
  nor3_1 U5778 ( .ip1(n11421), .ip2(n12126), .ip3(n6745), .op(n5235) );
  xnor2_1 U5779 ( .ip1(n5236), .ip2(n5235), .op(n5241) );
  nand2_1 U5780 ( .ip1(n5239), .ip2(n5241), .op(n5244) );
  nor2_1 U5781 ( .ip1(n13801), .ip2(n11858), .op(n11322) );
  nor2_1 U5782 ( .ip1(n5237), .ip2(n11322), .op(n5238) );
  nor2_1 U5783 ( .ip1(n5247), .ip2(n5238), .op(n5240) );
  nand2_1 U5784 ( .ip1(n5239), .ip2(n5240), .op(n5243) );
  nand2_1 U5785 ( .ip1(n5241), .ip2(n5240), .op(n5242) );
  nand3_1 U5786 ( .ip1(n5244), .ip2(n5243), .ip3(n5242), .op(n5250) );
  nand2_1 U5787 ( .ip1(n5248), .ip2(n5250), .op(n5253) );
  fulladder U5788 ( .a(n5247), .b(n5246), .ci(n5245), .co(n5254), .s(n5249) );
  nand2_1 U5789 ( .ip1(n5248), .ip2(n5249), .op(n5252) );
  nand2_1 U5790 ( .ip1(n5250), .ip2(n5249), .op(n5251) );
  nand3_1 U5791 ( .ip1(n5253), .ip2(n5252), .ip3(n5251), .op(n5255) );
  nand2_1 U5792 ( .ip1(n5254), .ip2(n5255), .op(n5258) );
  nand2_1 U5793 ( .ip1(n5256), .ip2(n5255), .op(n5257) );
  nand3_1 U5794 ( .ip1(n5259), .ip2(n5258), .ip3(n5257), .op(n5262) );
  nand2_1 U5795 ( .ip1(n5263), .ip2(n5262), .op(n5266) );
  nor2_1 U5796 ( .ip1(n5261), .ip2(n5260), .op(n5265) );
  nor2_1 U5797 ( .ip1(n5263), .ip2(n5262), .op(n5264) );
  ab_or_c_or_d U5798 ( .ip1(n5267), .ip2(n5266), .ip3(n5265), .ip4(n5264), 
        .op(n5268) );
  nand2_1 U5799 ( .ip1(n5269), .ip2(n5268), .op(n6765) );
  fulladder U5800 ( .a(n5272), .b(n5271), .ci(n5270), .co(n6764), .s(n5261) );
  inv_1 U5801 ( .ip(m1Inputs[21]), .op(n10866) );
  nor2_1 U5802 ( .ip1(n10476), .ip2(n10866), .op(n5340) );
  inv_1 U5803 ( .ip(m1Inputs[18]), .op(n10585) );
  nor2_1 U5804 ( .ip1(n10585), .ip2(n13801), .op(n5346) );
  inv_1 U5805 ( .ip(m1Inputs[16]), .op(n9995) );
  nor2_1 U5806 ( .ip1(n9995), .ip2(n12746), .op(n9768) );
  nand2_1 U5807 ( .ip1(n5056), .ip2(m1Inputs[20]), .op(n5273) );
  inv_1 U5808 ( .ip(m1Inputs[20]), .op(n10493) );
  nor4_1 U5809 ( .ip1(n6745), .ip2(n9047), .ip3(n10493), .ip4(n10866), .op(
        n5327) );
  or2_1 U5810 ( .ip1(n5273), .ip2(n5327), .op(n5276) );
  nand2_1 U5811 ( .ip1(n13707), .ip2(m1Inputs[21]), .op(n5274) );
  or2_1 U5812 ( .ip1(n5274), .ip2(n5327), .op(n5275) );
  nand2_1 U5813 ( .ip1(n5276), .ip2(n5275), .op(n5336) );
  inv_1 U5814 ( .ip(m1Inputs[17]), .op(n10472) );
  nor2_1 U5815 ( .ip1(n10472), .ip2(n4624), .op(n5298) );
  inv_1 U5816 ( .ip(m1Inputs[22]), .op(n10867) );
  nor2_1 U5817 ( .ip1(n13646), .ip2(n10867), .op(n5907) );
  nor2_1 U5818 ( .ip1(n9995), .ip2(n14289), .op(n9783) );
  and3_1 U5819 ( .ip1(n13707), .ip2(m1Inputs[22]), .ip3(n5323), .op(n5936) );
  buf_1 U5820 ( .ip(n13637), .op(n11974) );
  nand2_1 U5821 ( .ip1(m1Inputs[19]), .ip2(n11974), .op(n5299) );
  inv_1 U5822 ( .ip(m1Inputs[19]), .op(n10461) );
  nand2_1 U5823 ( .ip1(m1Inputs[18]), .ip2(n11974), .op(n5339) );
  nor3_1 U5824 ( .ip1(n10461), .ip2(n5339), .ip3(n13835), .op(n5280) );
  or2_1 U5825 ( .ip1(n5299), .ip2(n5280), .op(n5279) );
  nand2_1 U5826 ( .ip1(m1Inputs[18]), .ip2(n12699), .op(n5277) );
  or2_1 U5827 ( .ip1(n5277), .ip2(n5280), .op(n5278) );
  nand2_1 U5828 ( .ip1(n5279), .ip2(n5278), .op(n5288) );
  or2_1 U5829 ( .ip1(n5288), .ip2(n5280), .op(n5282) );
  nor2_1 U5830 ( .ip1(n9995), .ip2(n14384), .op(n10388) );
  or2_1 U5831 ( .ip1(n10388), .ip2(n5280), .op(n5281) );
  nand2_1 U5832 ( .ip1(n5282), .ip2(n5281), .op(n5914) );
  nand2_1 U5833 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[23]), .op(n6583)
         );
  nor3_1 U5834 ( .ip1(n10476), .ip2(n10493), .ip3(n6583), .op(n5294) );
  inv_1 U5835 ( .ip(m1Inputs[23]), .op(n10734) );
  nor2_1 U5836 ( .ip1(n10476), .ip2(n10734), .op(n5283) );
  or2_1 U5837 ( .ip1(m1Inputs[20]), .ip2(n5283), .op(n5285) );
  or2_1 U5838 ( .ip1(n9733), .ip2(n5283), .op(n5284) );
  nand2_1 U5839 ( .ip1(n5285), .ip2(n5284), .op(n5293) );
  nand2_1 U5840 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[21]), .op(n5295)
         );
  nor2_1 U5841 ( .ip1(n5293), .ip2(n5295), .op(n5286) );
  nor2_1 U5842 ( .ip1(n5294), .ip2(n5286), .op(n5913) );
  nand2_1 U5843 ( .ip1(m1Inputs[18]), .ip2(\STAGE_1/weightReg [6]), .op(n5912)
         );
  inv_1 U5844 ( .ip(n5287), .op(n5933) );
  inv_1 U5845 ( .ip(n10388), .op(n5289) );
  mux2_1 U5846 ( .ip1(n5289), .ip2(n10388), .s(n5288), .op(n5321) );
  nand4_1 U5847 ( .ip1(n4619), .ip2(n10507), .ip3(m1Inputs[19]), .ip4(
        m1Inputs[20]), .op(n5329) );
  nor2_1 U5848 ( .ip1(n13801), .ip2(n5329), .op(n5292) );
  nand2_1 U5849 ( .ip1(n5329), .ip2(m1Inputs[19]), .op(n5290) );
  mux2_1 U5850 ( .ip1(n5329), .ip2(n5290), .s(n9733), .op(n5338) );
  nor2_1 U5851 ( .ip1(n5339), .ip2(n5338), .op(n5291) );
  nor2_1 U5852 ( .ip1(n5292), .ip2(n5291), .op(n5320) );
  nor2_1 U5853 ( .ip1(n5294), .ip2(n5293), .op(n5296) );
  xor2_1 U5854 ( .ip1(n5296), .ip2(n5295), .op(n5319) );
  inv_1 U5855 ( .ip(n5297), .op(n5932) );
  nor2_1 U5856 ( .ip1(n10472), .ip2(n14836), .op(n5328) );
  fulladder U5857 ( .a(n5298), .b(n5907), .ci(n9783), .co(n5326), .s(n5335) );
  nor3_1 U5858 ( .ip1(n10493), .ip2(n13835), .ip3(n5299), .op(n5926) );
  inv_1 U5859 ( .ip(n5926), .op(n5302) );
  nand2_1 U5860 ( .ip1(m1Inputs[19]), .ip2(n12699), .op(n5300) );
  nand2_1 U5861 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[20]), .op(n5903)
         );
  nand2_1 U5862 ( .ip1(n5300), .ip2(n5903), .op(n5301) );
  nand2_1 U5863 ( .ip1(n5302), .ip2(n5301), .op(n5303) );
  nor3_1 U5864 ( .ip1(n10472), .ip2(n14384), .ip3(n5303), .op(n5925) );
  or2_1 U5865 ( .ip1(n5303), .ip2(n5925), .op(n5306) );
  nand2_1 U5866 ( .ip1(m1Inputs[17]), .ip2(n14835), .op(n5304) );
  or2_1 U5867 ( .ip1(n5304), .ip2(n5925), .op(n5305) );
  nand2_1 U5868 ( .ip1(n5306), .ip2(n5305), .op(n5930) );
  nand2_1 U5869 ( .ip1(m1Inputs[16]), .ip2(n14975), .op(n10417) );
  nand2_1 U5870 ( .ip1(m1Inputs[21]), .ip2(n12578), .op(n5307) );
  nand2_1 U5871 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[24]), .op(n6546)
         );
  nand2_1 U5872 ( .ip1(n5307), .ip2(n6546), .op(n5308) );
  nand3_1 U5873 ( .ip1(n12578), .ip2(m1Inputs[24]), .ip3(n5340), .op(n5922) );
  nand2_1 U5874 ( .ip1(n5308), .ip2(n5922), .op(n5309) );
  nor2_1 U5875 ( .ip1(n10417), .ip2(n5309), .op(n5923) );
  or2_1 U5876 ( .ip1(n10417), .ip2(n5923), .op(n5311) );
  or2_1 U5877 ( .ip1(n5309), .ip2(n5923), .op(n5310) );
  nand2_1 U5878 ( .ip1(n5311), .ip2(n5310), .op(n5929) );
  nand2_1 U5879 ( .ip1(n12809), .ip2(m1Inputs[23]), .op(n5312) );
  nand4_1 U5880 ( .ip1(n4619), .ip2(n10507), .ip3(m1Inputs[23]), .ip4(
        m1Inputs[22]), .op(n5918) );
  inv_1 U5881 ( .ip(n5918), .op(n5313) );
  or2_1 U5882 ( .ip1(n5312), .ip2(n5313), .op(n5316) );
  nand2_1 U5883 ( .ip1(n5056), .ip2(m1Inputs[22]), .op(n5314) );
  or2_1 U5884 ( .ip1(n5314), .ip2(n5313), .op(n5315) );
  nand2_1 U5885 ( .ip1(n5316), .ip2(n5315), .op(n5916) );
  inv_1 U5886 ( .ip(n5916), .op(n5318) );
  buf_1 U5887 ( .ip(n14768), .op(n13859) );
  nand2_1 U5888 ( .ip1(column[16]), .ip2(n13859), .op(n5317) );
  mux2_1 U5889 ( .ip1(n5318), .ip2(n5916), .s(n5317), .op(n5928) );
  fulladder U5890 ( .a(n5321), .b(n5320), .ci(n5319), .co(n5297), .s(n5322) );
  inv_1 U5891 ( .ip(n5322), .op(n5399) );
  nor2_1 U5892 ( .ip1(n13570), .ip2(n10867), .op(n5324) );
  nor2_1 U5893 ( .ip1(n5324), .ip2(n5323), .op(n5325) );
  nor2_1 U5894 ( .ip1(n5936), .ip2(n5325), .op(n5398) );
  fulladder U5895 ( .a(n5328), .b(n5327), .ci(n5326), .co(n5931), .s(n5397) );
  nor2_1 U5896 ( .ip1(n10585), .ip2(n9047), .op(n5361) );
  and3_1 U5897 ( .ip1(n4672), .ip2(n5361), .ip3(m1Inputs[19]), .op(n5351) );
  inv_1 U5898 ( .ip(n5329), .op(n5334) );
  nor2_1 U5899 ( .ip1(n6745), .ip2(n10461), .op(n5330) );
  or2_1 U5900 ( .ip1(m1Inputs[20]), .ip2(n5330), .op(n5332) );
  or2_1 U5901 ( .ip1(n13707), .ip2(n5330), .op(n5331) );
  nand2_1 U5902 ( .ip1(n5332), .ip2(n5331), .op(n5333) );
  nor2_1 U5903 ( .ip1(n5334), .ip2(n5333), .op(n5342) );
  nor2_1 U5904 ( .ip1(n10472), .ip2(n14783), .op(n5341) );
  fulladder U5905 ( .a(n5337), .b(n5336), .ci(n5335), .co(n5323), .s(n5344) );
  xor2_1 U5906 ( .ip1(n5339), .ip2(n5338), .op(n5343) );
  and2_1 U5907 ( .ip1(n5394), .ip2(n5393), .op(n5388) );
  fulladder U5908 ( .a(n5340), .b(n5346), .ci(n9768), .co(n5337), .s(n5380) );
  fulladder U5909 ( .a(n5351), .b(n5342), .ci(n5341), .co(n5345), .s(n5379) );
  nor2_1 U5910 ( .ip1(n10476), .ip2(n10493), .op(n5353) );
  nor2_1 U5911 ( .ip1(n9995), .ip2(n14783), .op(n9851) );
  nor2_1 U5912 ( .ip1(n10472), .ip2(n13801), .op(n5352) );
  fulladder U5913 ( .a(n5345), .b(n5344), .ci(n5343), .co(n5393), .s(n5390) );
  nor3_1 U5914 ( .ip1(n5388), .ip2(n5389), .ip3(n5390), .op(n5392) );
  nor2_1 U5915 ( .ip1(n9995), .ip2(n13570), .op(n10032) );
  and2_1 U5916 ( .ip1(n10032), .ip2(n5346), .op(n5363) );
  nor2_1 U5917 ( .ip1(n13570), .ip2(n10461), .op(n5347) );
  or2_1 U5918 ( .ip1(n4619), .ip2(n5347), .op(n5349) );
  or2_1 U5919 ( .ip1(m1Inputs[18]), .ip2(n5347), .op(n5348) );
  nand2_1 U5920 ( .ip1(n5349), .ip2(n5348), .op(n5350) );
  nor2_1 U5921 ( .ip1(n5351), .ip2(n5350), .op(n5355) );
  fulladder U5922 ( .a(n5353), .b(n9851), .ci(n5352), .co(n5378), .s(n5354) );
  fulladder U5923 ( .a(n5363), .b(n5355), .ci(n5354), .co(n5381), .s(n5374) );
  nand2_1 U5924 ( .ip1(n13707), .ip2(m1Inputs[17]), .op(n5359) );
  nor2_1 U5925 ( .ip1(n6745), .ip2(n9995), .op(n9964) );
  inv_1 U5926 ( .ip(n9964), .op(n5371) );
  or2_1 U5927 ( .ip1(n10032), .ip2(m1Inputs[18]), .op(n5357) );
  or2_1 U5928 ( .ip1(n13854), .ip2(m1Inputs[18]), .op(n5356) );
  nand2_1 U5929 ( .ip1(n5357), .ip2(n5356), .op(n5358) );
  not_ab_or_c_or_d U5930 ( .ip1(n5359), .ip2(n5371), .ip3(n5358), .ip4(n13646), 
        .op(n5364) );
  nor3_1 U5931 ( .ip1(n10032), .ip2(n6745), .ip3(n10472), .op(n5370) );
  nor2_1 U5932 ( .ip1(n13646), .ip2(n10461), .op(n5360) );
  xor2_1 U5933 ( .ip1(n5370), .ip2(n5360), .op(n5366) );
  nand2_1 U5934 ( .ip1(n5364), .ip2(n5366), .op(n5369) );
  nor2_1 U5935 ( .ip1(n9995), .ip2(n13801), .op(n9914) );
  nor2_1 U5936 ( .ip1(n5361), .ip2(n9914), .op(n5362) );
  nor2_1 U5937 ( .ip1(n5363), .ip2(n5362), .op(n5365) );
  nand2_1 U5938 ( .ip1(n5364), .ip2(n5365), .op(n5368) );
  nand2_1 U5939 ( .ip1(n5366), .ip2(n5365), .op(n5367) );
  nand3_1 U5940 ( .ip1(n5369), .ip2(n5368), .ip3(n5367), .op(n5375) );
  nor2_1 U5941 ( .ip1(n5374), .ip2(n5375), .op(n5377) );
  and3_1 U5942 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n5370), .ip3(m1Inputs[19]), 
        .op(n5373) );
  nor3_1 U5943 ( .ip1(n9047), .ip2(n10472), .ip3(n5371), .op(n5372) );
  not_ab_or_c_or_d U5944 ( .ip1(n5375), .ip2(n5374), .ip3(n5373), .ip4(n5372), 
        .op(n5376) );
  nor2_1 U5945 ( .ip1(n5377), .ip2(n5376), .op(n5383) );
  nand2_1 U5946 ( .ip1(n5381), .ip2(n5383), .op(n5386) );
  fulladder U5947 ( .a(n5380), .b(n5379), .ci(n5378), .co(n5389), .s(n5382) );
  nand2_1 U5948 ( .ip1(n5381), .ip2(n5382), .op(n5385) );
  nand2_1 U5949 ( .ip1(n5383), .ip2(n5382), .op(n5384) );
  nand3_1 U5950 ( .ip1(n5386), .ip2(n5385), .ip3(n5384), .op(n5387) );
  not_ab_or_c_or_d U5951 ( .ip1(n5390), .ip2(n5389), .ip3(n5388), .ip4(n5387), 
        .op(n5391) );
  or2_1 U5952 ( .ip1(n5392), .ip2(n5391), .op(n5396) );
  nor2_1 U5953 ( .ip1(n5394), .ip2(n5393), .op(n5395) );
  nor2_1 U5954 ( .ip1(n5396), .ip2(n5395), .op(n5938) );
  fulladder U5955 ( .a(n5399), .b(n5398), .ci(n5397), .co(n5937), .s(n5394) );
  inv_1 U5956 ( .ip(m1Inputs[85]), .op(n13847) );
  nor2_1 U5957 ( .ip1(n10476), .ip2(n13847), .op(n5461) );
  inv_1 U5958 ( .ip(m1Inputs[82]), .op(n13830) );
  nor2_1 U5959 ( .ip1(n13801), .ip2(n13830), .op(n5460) );
  inv_1 U5960 ( .ip(m1Inputs[80]), .op(n13807) );
  nor2_1 U5961 ( .ip1(n13807), .ip2(n13835), .op(n5459) );
  nand2_1 U5962 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[84]), .op(n5400)
         );
  inv_1 U5963 ( .ip(m1Inputs[84]), .op(n13765) );
  nor4_1 U5964 ( .ip1(n6745), .ip2(n9047), .ip3(n13765), .ip4(n13847), .op(
        n5444) );
  or2_1 U5965 ( .ip1(n5400), .ip2(n5444), .op(n5403) );
  nand2_1 U5966 ( .ip1(n13707), .ip2(m1Inputs[85]), .op(n5401) );
  or2_1 U5967 ( .ip1(n5401), .ip2(n5444), .op(n5402) );
  nand2_1 U5968 ( .ip1(n5403), .ip2(n5402), .op(n5453) );
  inv_1 U5969 ( .ip(m1Inputs[81]), .op(n13841) );
  nor2_1 U5970 ( .ip1(n13841), .ip2(n12746), .op(n5426) );
  inv_1 U5971 ( .ip(m1Inputs[86]), .op(n13578) );
  nor2_1 U5972 ( .ip1(n10476), .ip2(n13578), .op(n6345) );
  nor2_1 U5973 ( .ip1(n13807), .ip2(n14836), .op(n5425) );
  and3_1 U5974 ( .ip1(n10507), .ip2(m1Inputs[86]), .ip3(n5440), .op(n6383) );
  nand2_1 U5975 ( .ip1(m1Inputs[83]), .ip2(n13637), .op(n5427) );
  inv_1 U5976 ( .ip(m1Inputs[83]), .op(n13654) );
  nand2_1 U5977 ( .ip1(m1Inputs[82]), .ip2(n13637), .op(n5456) );
  nor3_1 U5978 ( .ip1(n13654), .ip2(n5456), .ip3(n13835), .op(n5407) );
  or2_1 U5979 ( .ip1(n5427), .ip2(n5407), .op(n5406) );
  nand2_1 U5980 ( .ip1(m1Inputs[82]), .ip2(\STAGE_1/weightReg [5]), .op(n5404)
         );
  or2_1 U5981 ( .ip1(n5404), .ip2(n5407), .op(n5405) );
  nand2_1 U5982 ( .ip1(n5406), .ip2(n5405), .op(n5418) );
  or2_1 U5983 ( .ip1(n5418), .ip2(n5407), .op(n5409) );
  nor2_1 U5984 ( .ip1(n13807), .ip2(n14384), .op(n5417) );
  or2_1 U5985 ( .ip1(n5417), .ip2(n5407), .op(n5408) );
  nand2_1 U5986 ( .ip1(n5409), .ip2(n5408), .op(n6352) );
  nand2_1 U5987 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[87]), .op(n6395)
         );
  nor2_1 U5988 ( .ip1(n10476), .ip2(n13765), .op(n5472) );
  and3_1 U5989 ( .ip1(n12578), .ip2(m1Inputs[87]), .ip3(n5472), .op(n5413) );
  or2_1 U5990 ( .ip1(n6395), .ip2(n5413), .op(n5412) );
  nand2_1 U5991 ( .ip1(n13614), .ip2(m1Inputs[84]), .op(n5410) );
  or2_1 U5992 ( .ip1(n5410), .ip2(n5413), .op(n5411) );
  nand2_1 U5993 ( .ip1(n5412), .ip2(n5411), .op(n5423) );
  or2_1 U5994 ( .ip1(n5423), .ip2(n5413), .op(n5415) );
  nor2_1 U5995 ( .ip1(n13854), .ip2(n13847), .op(n5422) );
  or2_1 U5996 ( .ip1(n5422), .ip2(n5413), .op(n5414) );
  nand2_1 U5997 ( .ip1(n5415), .ip2(n5414), .op(n6351) );
  nand2_1 U5998 ( .ip1(m1Inputs[82]), .ip2(n12981), .op(n6350) );
  inv_1 U5999 ( .ip(n5416), .op(n6380) );
  xnor2_1 U6000 ( .ip1(n5418), .ip2(n5417), .op(n5438) );
  nand4_1 U6001 ( .ip1(n4672), .ip2(\STAGE_1/weightReg [1]), .ip3(m1Inputs[83]), .ip4(m1Inputs[84]), .op(n5446) );
  nor2_1 U6002 ( .ip1(n13801), .ip2(n5446), .op(n5421) );
  nand2_1 U6003 ( .ip1(n5446), .ip2(m1Inputs[83]), .op(n5419) );
  mux2_1 U6004 ( .ip1(n5446), .ip2(n5419), .s(n13614), .op(n5455) );
  nor2_1 U6005 ( .ip1(n5456), .ip2(n5455), .op(n5420) );
  nor2_1 U6006 ( .ip1(n5421), .ip2(n5420), .op(n5437) );
  xnor2_1 U6007 ( .ip1(n5423), .ip2(n5422), .op(n5436) );
  inv_1 U6008 ( .ip(n5424), .op(n6379) );
  nor2_1 U6009 ( .ip1(n13841), .ip2(n14836), .op(n5445) );
  fulladder U6010 ( .a(n5426), .b(n6345), .ci(n5425), .co(n5443), .s(n5452) );
  nand2_1 U6011 ( .ip1(m1Inputs[83]), .ip2(n14369), .op(n5428) );
  nor3_1 U6012 ( .ip1(n13765), .ip2(n12746), .ip3(n5427), .op(n6366) );
  or2_1 U6013 ( .ip1(n5428), .ip2(n6366), .op(n5430) );
  nand2_1 U6014 ( .ip1(n13637), .ip2(m1Inputs[84]), .op(n6341) );
  or2_1 U6015 ( .ip1(n6341), .ip2(n6366), .op(n5429) );
  nand2_1 U6016 ( .ip1(n5430), .ip2(n5429), .op(n6365) );
  nor2_1 U6017 ( .ip1(n13841), .ip2(n14368), .op(n6367) );
  xor2_1 U6018 ( .ip1(n6365), .ip2(n6367), .op(n6377) );
  and3_1 U6019 ( .ip1(n12578), .ip2(m1Inputs[88]), .ip3(n5461), .op(n6361) );
  inv_1 U6020 ( .ip(m1Inputs[88]), .op(n13748) );
  nor2_1 U6021 ( .ip1(n13646), .ip2(n13748), .op(n6447) );
  or2_1 U6022 ( .ip1(m1Inputs[85]), .ip2(n6447), .op(n5432) );
  or2_1 U6023 ( .ip1(n9733), .ip2(n6447), .op(n5431) );
  nand2_1 U6024 ( .ip1(n5432), .ip2(n5431), .op(n5433) );
  nor2_1 U6025 ( .ip1(n6361), .ip2(n5433), .op(n6360) );
  nor2_1 U6026 ( .ip1(n13807), .ip2(n6504), .op(n6362) );
  xor2_1 U6027 ( .ip1(n6360), .ip2(n6362), .op(n6376) );
  nand2_1 U6028 ( .ip1(m1Inputs[86]), .ip2(n4672), .op(n5434) );
  nand2_1 U6029 ( .ip1(n13707), .ip2(m1Inputs[87]), .op(n6370) );
  nand2_1 U6030 ( .ip1(n5434), .ip2(n6370), .op(n5435) );
  nand4_1 U6031 ( .ip1(n4672), .ip2(n10507), .ip3(m1Inputs[87]), .ip4(
        m1Inputs[86]), .op(n6354) );
  nand2_1 U6032 ( .ip1(n5435), .ip2(n6354), .op(n6356) );
  nand2_1 U6033 ( .ip1(column[80]), .ip2(n13859), .op(n6355) );
  xor2_1 U6034 ( .ip1(n6356), .ip2(n6355), .op(n6375) );
  fulladder U6035 ( .a(n5438), .b(n5437), .ci(n5436), .co(n5424), .s(n5439) );
  inv_1 U6036 ( .ip(n5439), .op(n5520) );
  nor2_1 U6037 ( .ip1(n13570), .ip2(n13578), .op(n5441) );
  nor2_1 U6038 ( .ip1(n5441), .ip2(n5440), .op(n5442) );
  nor2_1 U6039 ( .ip1(n6383), .ip2(n5442), .op(n5519) );
  fulladder U6040 ( .a(n5445), .b(n5444), .ci(n5443), .co(n6378), .s(n5518) );
  nand2_1 U6041 ( .ip1(n13707), .ip2(m1Inputs[82]), .op(n5478) );
  nor3_1 U6042 ( .ip1(n13709), .ip2(n13654), .ip3(n5478), .op(n5469) );
  inv_1 U6043 ( .ip(n5446), .op(n5451) );
  nor2_1 U6044 ( .ip1(n13854), .ip2(n13654), .op(n5447) );
  or2_1 U6045 ( .ip1(m1Inputs[84]), .ip2(n5447), .op(n5449) );
  or2_1 U6046 ( .ip1(n10507), .ip2(n5447), .op(n5448) );
  nand2_1 U6047 ( .ip1(n5449), .ip2(n5448), .op(n5450) );
  nor2_1 U6048 ( .ip1(n5451), .ip2(n5450), .op(n5458) );
  nor2_1 U6049 ( .ip1(n13841), .ip2(n14783), .op(n5457) );
  fulladder U6050 ( .a(n5454), .b(n5453), .ci(n5452), .co(n5440), .s(n5463) );
  xor2_1 U6051 ( .ip1(n5456), .ip2(n5455), .op(n5462) );
  nand2_1 U6052 ( .ip1(n5512), .ip2(n5511), .op(n5517) );
  fulladder U6053 ( .a(n5469), .b(n5458), .ci(n5457), .co(n5464), .s(n5501) );
  nor2_1 U6054 ( .ip1(n13801), .ip2(n13841), .op(n5471) );
  nor2_1 U6055 ( .ip1(n13807), .ip2(n14783), .op(n5470) );
  fulladder U6056 ( .a(n5461), .b(n5460), .ci(n5459), .co(n5454), .s(n5499) );
  fulladder U6057 ( .a(n5464), .b(n5463), .ci(n5462), .co(n5511), .s(n5509) );
  nand2_1 U6058 ( .ip1(n5510), .ip2(n5509), .op(n5508) );
  nor4_1 U6059 ( .ip1(n13570), .ip2(n13801), .ip3(n13807), .ip4(n13830), .op(
        n5498) );
  nor2_1 U6060 ( .ip1(n13570), .ip2(n13654), .op(n5465) );
  or2_1 U6061 ( .ip1(m1Inputs[82]), .ip2(n5465), .op(n5467) );
  or2_1 U6062 ( .ip1(n4672), .ip2(n5465), .op(n5466) );
  nand2_1 U6063 ( .ip1(n5467), .ip2(n5466), .op(n5468) );
  nor2_1 U6064 ( .ip1(n5469), .ip2(n5468), .op(n5497) );
  fulladder U6065 ( .a(n5472), .b(n5471), .ci(n5470), .co(n5500), .s(n5496) );
  nand2_1 U6066 ( .ip1(n13707), .ip2(m1Inputs[81]), .op(n5477) );
  nand2_1 U6067 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[80]), .op(n5476)
         );
  or2_1 U6068 ( .ip1(m1Inputs[80]), .ip2(m1Inputs[82]), .op(n5474) );
  or2_1 U6069 ( .ip1(n13854), .ip2(m1Inputs[82]), .op(n5473) );
  nand2_1 U6070 ( .ip1(n5474), .ip2(n5473), .op(n5475) );
  not_ab_or_c_or_d U6071 ( .ip1(n5477), .ip2(n5476), .ip3(n5475), .ip4(n10476), 
        .op(n5483) );
  or2_1 U6072 ( .ip1(n5478), .ip2(n5498), .op(n5481) );
  nand2_1 U6073 ( .ip1(n13614), .ip2(m1Inputs[80]), .op(n5479) );
  or2_1 U6074 ( .ip1(n5479), .ip2(n5498), .op(n5480) );
  nand2_1 U6075 ( .ip1(n5481), .ip2(n5480), .op(n5485) );
  nand2_1 U6076 ( .ip1(n5483), .ip2(n5485), .op(n5488) );
  not_ab_or_c_or_d U6077 ( .ip1(n10507), .ip2(m1Inputs[80]), .ip3(n10555), 
        .ip4(n13841), .op(n5489) );
  nor2_1 U6078 ( .ip1(n13646), .ip2(n13654), .op(n5482) );
  xor2_1 U6079 ( .ip1(n5489), .ip2(n5482), .op(n5484) );
  nand2_1 U6080 ( .ip1(n5483), .ip2(n5484), .op(n5487) );
  nand2_1 U6081 ( .ip1(n5485), .ip2(n5484), .op(n5486) );
  nand3_1 U6082 ( .ip1(n5488), .ip2(n5487), .ip3(n5486), .op(n5493) );
  nor2_1 U6083 ( .ip1(n5492), .ip2(n5493), .op(n5495) );
  nor4_1 U6084 ( .ip1(n6745), .ip2(n9047), .ip3(n13841), .ip4(n13807), .op(
        n5491) );
  and3_1 U6085 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n5489), .ip3(m1Inputs[83]), 
        .op(n5490) );
  not_ab_or_c_or_d U6086 ( .ip1(n5493), .ip2(n5492), .ip3(n5491), .ip4(n5490), 
        .op(n5494) );
  or2_1 U6087 ( .ip1(n5495), .ip2(n5494), .op(n5503) );
  fulladder U6088 ( .a(n5498), .b(n5497), .ci(n5496), .co(n5505), .s(n5492) );
  fulladder U6089 ( .a(n5501), .b(n5500), .ci(n5499), .co(n5510), .s(n5504) );
  nor2_1 U6090 ( .ip1(n5505), .ip2(n5504), .op(n5502) );
  or2_1 U6091 ( .ip1(n5503), .ip2(n5502), .op(n5507) );
  nand2_1 U6092 ( .ip1(n5505), .ip2(n5504), .op(n5506) );
  nand3_1 U6093 ( .ip1(n5508), .ip2(n5507), .ip3(n5506), .op(n5515) );
  or2_1 U6094 ( .ip1(n5510), .ip2(n5509), .op(n5514) );
  or2_1 U6095 ( .ip1(n5512), .ip2(n5511), .op(n5513) );
  nand3_1 U6096 ( .ip1(n5515), .ip2(n5514), .ip3(n5513), .op(n5516) );
  nand2_1 U6097 ( .ip1(n5517), .ip2(n5516), .op(n6385) );
  fulladder U6098 ( .a(n5520), .b(n5519), .ci(n5518), .co(n6384), .s(n5512) );
  inv_1 U6099 ( .ip(m1Inputs[34]), .op(n11539) );
  inv_1 U6100 ( .ip(m1Inputs[37]), .op(n11555) );
  nor4_1 U6101 ( .ip1(n10476), .ip2(n13487), .ip3(n11539), .ip4(n11555), .op(
        n5521) );
  inv_1 U6102 ( .ip(n5521), .op(n5526) );
  nand2_1 U6103 ( .ip1(n13803), .ip2(m1Inputs[37]), .op(n5558) );
  or2_1 U6104 ( .ip1(n5558), .ip2(n5521), .op(n5524) );
  nand2_1 U6105 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[34]), .op(n5522)
         );
  or2_1 U6106 ( .ip1(n5522), .ip2(n5521), .op(n5523) );
  nand2_1 U6107 ( .ip1(n5524), .ip2(n5523), .op(n5588) );
  inv_1 U6108 ( .ip(m1Inputs[32]), .op(n11516) );
  nor2_1 U6109 ( .ip1(n11516), .ip2(n12746), .op(n5587) );
  nand2_1 U6110 ( .ip1(n5588), .ip2(n5587), .op(n5525) );
  nand2_1 U6111 ( .ip1(n5526), .ip2(n5525), .op(n5582) );
  nand2_1 U6112 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[36]), .op(n5527)
         );
  inv_1 U6113 ( .ip(m1Inputs[36]), .op(n11477) );
  nor4_1 U6114 ( .ip1(n6745), .ip2(n9047), .ip3(n11477), .ip4(n11555), .op(
        n5572) );
  or2_1 U6115 ( .ip1(n5527), .ip2(n5572), .op(n5530) );
  nand2_1 U6116 ( .ip1(n12809), .ip2(m1Inputs[37]), .op(n5528) );
  or2_1 U6117 ( .ip1(n5528), .ip2(n5572), .op(n5529) );
  nand2_1 U6118 ( .ip1(n5530), .ip2(n5529), .op(n5581) );
  inv_1 U6119 ( .ip(m1Inputs[33]), .op(n11549) );
  nor2_1 U6120 ( .ip1(n11549), .ip2(n12746), .op(n5553) );
  inv_1 U6121 ( .ip(m1Inputs[38]), .op(n11283) );
  nor2_1 U6122 ( .ip1(n13646), .ip2(n11283), .op(n6193) );
  nor2_1 U6123 ( .ip1(n11516), .ip2(n14289), .op(n5552) );
  and3_1 U6124 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[38]), .ip3(n5568), 
        .op(n6231) );
  nand2_1 U6125 ( .ip1(m1Inputs[35]), .ip2(n11974), .op(n5554) );
  inv_1 U6126 ( .ip(m1Inputs[35]), .op(n11370) );
  nand2_1 U6127 ( .ip1(m1Inputs[34]), .ip2(n11974), .op(n5584) );
  nor3_1 U6128 ( .ip1(n11370), .ip2(n5584), .ip3(n8942), .op(n5534) );
  or2_1 U6129 ( .ip1(n5554), .ip2(n5534), .op(n5533) );
  nand2_1 U6130 ( .ip1(m1Inputs[34]), .ip2(n12699), .op(n5531) );
  or2_1 U6131 ( .ip1(n5531), .ip2(n5534), .op(n5532) );
  nand2_1 U6132 ( .ip1(n5533), .ip2(n5532), .op(n5545) );
  or2_1 U6133 ( .ip1(n5545), .ip2(n5534), .op(n5536) );
  nor2_1 U6134 ( .ip1(n11516), .ip2(n12156), .op(n5544) );
  or2_1 U6135 ( .ip1(n5544), .ip2(n5534), .op(n5535) );
  nand2_1 U6136 ( .ip1(n5536), .ip2(n5535), .op(n6200) );
  nand2_1 U6137 ( .ip1(n13803), .ip2(m1Inputs[39]), .op(n6243) );
  nor2_1 U6138 ( .ip1(n13646), .ip2(n11477), .op(n5600) );
  and3_1 U6139 ( .ip1(n12578), .ip2(m1Inputs[39]), .ip3(n5600), .op(n5540) );
  or2_1 U6140 ( .ip1(n6243), .ip2(n5540), .op(n5539) );
  nand2_1 U6141 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[36]), .op(n5537)
         );
  or2_1 U6142 ( .ip1(n5537), .ip2(n5540), .op(n5538) );
  nand2_1 U6143 ( .ip1(n5539), .ip2(n5538), .op(n5550) );
  or2_1 U6144 ( .ip1(n5550), .ip2(n5540), .op(n5542) );
  nor2_1 U6145 ( .ip1(n13854), .ip2(n11555), .op(n5549) );
  or2_1 U6146 ( .ip1(n5549), .ip2(n5540), .op(n5541) );
  nand2_1 U6147 ( .ip1(n5542), .ip2(n5541), .op(n6199) );
  nand2_1 U6148 ( .ip1(m1Inputs[34]), .ip2(n12981), .op(n6198) );
  inv_1 U6149 ( .ip(n5543), .op(n6228) );
  xnor2_1 U6150 ( .ip1(n5545), .ip2(n5544), .op(n5566) );
  nand4_1 U6151 ( .ip1(n4672), .ip2(n10507), .ip3(m1Inputs[35]), .ip4(
        m1Inputs[36]), .op(n5574) );
  nor2_1 U6152 ( .ip1(n13801), .ip2(n5574), .op(n5548) );
  nand2_1 U6153 ( .ip1(n5574), .ip2(m1Inputs[35]), .op(n5546) );
  mux2_1 U6154 ( .ip1(n5574), .ip2(n5546), .s(n9733), .op(n5583) );
  nor2_1 U6155 ( .ip1(n5584), .ip2(n5583), .op(n5547) );
  nor2_1 U6156 ( .ip1(n5548), .ip2(n5547), .op(n5565) );
  xnor2_1 U6157 ( .ip1(n5550), .ip2(n5549), .op(n5564) );
  inv_1 U6158 ( .ip(n5551), .op(n6227) );
  nor2_1 U6159 ( .ip1(n11549), .ip2(n14289), .op(n5573) );
  fulladder U6160 ( .a(n5553), .b(n6193), .ci(n5552), .co(n5571), .s(n5580) );
  nand2_1 U6161 ( .ip1(m1Inputs[35]), .ip2(n12699), .op(n5555) );
  nor3_1 U6162 ( .ip1(n11477), .ip2(n13835), .ip3(n5554), .op(n6214) );
  or2_1 U6163 ( .ip1(n5555), .ip2(n6214), .op(n5557) );
  nand2_1 U6164 ( .ip1(n11974), .ip2(m1Inputs[36]), .op(n6189) );
  or2_1 U6165 ( .ip1(n6189), .ip2(n6214), .op(n5556) );
  nand2_1 U6166 ( .ip1(n5557), .ip2(n5556), .op(n6213) );
  nor2_1 U6167 ( .ip1(n11549), .ip2(n12156), .op(n6215) );
  xor2_1 U6168 ( .ip1(n6213), .ip2(n6215), .op(n6225) );
  nand2_1 U6169 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[37]), .op(n5559)
         );
  inv_1 U6170 ( .ip(m1Inputs[40]), .op(n11461) );
  nor3_1 U6171 ( .ip1(n13082), .ip2(n11461), .ip3(n5558), .op(n6209) );
  or2_1 U6172 ( .ip1(n5559), .ip2(n6209), .op(n5561) );
  nand2_1 U6173 ( .ip1(n13803), .ip2(m1Inputs[40]), .op(n6295) );
  or2_1 U6174 ( .ip1(n6295), .ip2(n6209), .op(n5560) );
  nand2_1 U6175 ( .ip1(n5561), .ip2(n5560), .op(n6208) );
  nor2_1 U6176 ( .ip1(n11516), .ip2(n6503), .op(n6210) );
  xor2_1 U6177 ( .ip1(n6208), .ip2(n6210), .op(n6224) );
  nand2_1 U6178 ( .ip1(m1Inputs[38]), .ip2(n4619), .op(n5562) );
  nand2_1 U6179 ( .ip1(n12809), .ip2(m1Inputs[39]), .op(n6218) );
  nand2_1 U6180 ( .ip1(n5562), .ip2(n6218), .op(n5563) );
  nand4_1 U6181 ( .ip1(n4672), .ip2(\STAGE_1/weightReg [1]), .ip3(m1Inputs[39]), .ip4(m1Inputs[38]), .op(n6202) );
  nand2_1 U6182 ( .ip1(n5563), .ip2(n6202), .op(n6204) );
  buf_1 U6183 ( .ip(n14768), .op(n13039) );
  nand2_1 U6184 ( .ip1(column[32]), .ip2(n13039), .op(n6203) );
  xor2_1 U6185 ( .ip1(n6204), .ip2(n6203), .op(n6223) );
  fulladder U6186 ( .a(n5566), .b(n5565), .ci(n5564), .co(n5551), .s(n5567) );
  inv_1 U6187 ( .ip(n5567), .op(n5648) );
  nor2_1 U6188 ( .ip1(n13570), .ip2(n11283), .op(n5569) );
  nor2_1 U6189 ( .ip1(n5569), .ip2(n5568), .op(n5570) );
  nor2_1 U6190 ( .ip1(n6231), .ip2(n5570), .op(n5647) );
  fulladder U6191 ( .a(n5573), .b(n5572), .ci(n5571), .co(n6226), .s(n5646) );
  nand2_1 U6192 ( .ip1(n12809), .ip2(m1Inputs[34]), .op(n5612) );
  nor3_1 U6193 ( .ip1(n13709), .ip2(n11370), .ip3(n5612), .op(n5597) );
  inv_1 U6194 ( .ip(n5574), .op(n5579) );
  nor2_1 U6195 ( .ip1(n13854), .ip2(n11370), .op(n5575) );
  or2_1 U6196 ( .ip1(m1Inputs[36]), .ip2(n5575), .op(n5577) );
  or2_1 U6197 ( .ip1(n10507), .ip2(n5575), .op(n5576) );
  nand2_1 U6198 ( .ip1(n5577), .ip2(n5576), .op(n5578) );
  nor2_1 U6199 ( .ip1(n5579), .ip2(n5578), .op(n5586) );
  nor2_1 U6200 ( .ip1(n11549), .ip2(n14783), .op(n5585) );
  fulladder U6201 ( .a(n5582), .b(n5581), .ci(n5580), .co(n5568), .s(n5591) );
  xor2_1 U6202 ( .ip1(n5584), .ip2(n5583), .op(n5590) );
  nand2_1 U6203 ( .ip1(n5637), .ip2(n5636), .op(n5645) );
  fulladder U6204 ( .a(n5597), .b(n5586), .ci(n5585), .co(n5592), .s(n5629) );
  nor2_1 U6205 ( .ip1(n13801), .ip2(n11549), .op(n5599) );
  nor2_1 U6206 ( .ip1(n11516), .ip2(n14783), .op(n5598) );
  xor2_1 U6207 ( .ip1(n5588), .ip2(n5587), .op(n5627) );
  inv_1 U6208 ( .ip(n5589), .op(n5643) );
  fulladder U6209 ( .a(n5592), .b(n5591), .ci(n5590), .co(n5636), .s(n5639) );
  nor4_1 U6210 ( .ip1(n13570), .ip2(n13082), .ip3(n11516), .ip4(n11539), .op(
        n5613) );
  nor2_1 U6211 ( .ip1(n13570), .ip2(n11370), .op(n5593) );
  or2_1 U6212 ( .ip1(m1Inputs[34]), .ip2(n5593), .op(n5595) );
  or2_1 U6213 ( .ip1(n4619), .ip2(n5593), .op(n5594) );
  nand2_1 U6214 ( .ip1(n5595), .ip2(n5594), .op(n5596) );
  nor2_1 U6215 ( .ip1(n5597), .ip2(n5596), .op(n5602) );
  fulladder U6216 ( .a(n5600), .b(n5599), .ci(n5598), .co(n5628), .s(n5601) );
  fulladder U6217 ( .a(n5613), .b(n5602), .ci(n5601), .co(n5630), .s(n5620) );
  nand2_1 U6218 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[35]), .op(n5605)
         );
  nand4_1 U6219 ( .ip1(n4619), .ip2(\STAGE_1/weightReg [1]), .ip3(m1Inputs[33]), .ip4(m1Inputs[32]), .op(n5604) );
  and2_1 U6220 ( .ip1(n5605), .ip2(n5604), .op(n5603) );
  nor3_1 U6221 ( .ip1(n5603), .ip2(n11549), .ip3(n6745), .op(n5619) );
  nand2_1 U6222 ( .ip1(n5620), .ip2(n5619), .op(n5626) );
  xor2_1 U6223 ( .ip1(n5605), .ip2(n5604), .op(n5607) );
  nand2_1 U6224 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[33]), .op(n5606)
         );
  xor2_1 U6225 ( .ip1(n5607), .ip2(n5606), .op(n5624) );
  nand2_1 U6226 ( .ip1(n12809), .ip2(m1Inputs[33]), .op(n5609) );
  nand2_1 U6227 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[32]), .op(n5608)
         );
  not_ab_or_c_or_d U6228 ( .ip1(n5609), .ip2(n5608), .ip3(n13646), .ip4(n11539), .op(n5611) );
  nor4_1 U6229 ( .ip1(n9047), .ip2(n11549), .ip3(n11516), .ip4(n5739), .op(
        n5610) );
  nor2_1 U6230 ( .ip1(n5611), .ip2(n5610), .op(n5623) );
  or2_1 U6231 ( .ip1(n5612), .ip2(n5613), .op(n5616) );
  nand2_1 U6232 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[32]), .op(n5614)
         );
  or2_1 U6233 ( .ip1(n5614), .ip2(n5613), .op(n5615) );
  nand2_1 U6234 ( .ip1(n5616), .ip2(n5615), .op(n5618) );
  nor2_1 U6235 ( .ip1(n5623), .ip2(n5624), .op(n5617) );
  nor2_1 U6236 ( .ip1(n5618), .ip2(n5617), .op(n5622) );
  nor2_1 U6237 ( .ip1(n5620), .ip2(n5619), .op(n5621) );
  ab_or_c_or_d U6238 ( .ip1(n5624), .ip2(n5623), .ip3(n5622), .ip4(n5621), 
        .op(n5625) );
  nand2_1 U6239 ( .ip1(n5626), .ip2(n5625), .op(n5632) );
  nand2_1 U6240 ( .ip1(n5630), .ip2(n5632), .op(n5635) );
  fulladder U6241 ( .a(n5629), .b(n5628), .ci(n5627), .co(n5589), .s(n5631) );
  nand2_1 U6242 ( .ip1(n5630), .ip2(n5631), .op(n5634) );
  nand2_1 U6243 ( .ip1(n5632), .ip2(n5631), .op(n5633) );
  nand3_1 U6244 ( .ip1(n5635), .ip2(n5634), .ip3(n5633), .op(n5638) );
  nand2_1 U6245 ( .ip1(n5639), .ip2(n5638), .op(n5642) );
  nor2_1 U6246 ( .ip1(n5637), .ip2(n5636), .op(n5641) );
  nor2_1 U6247 ( .ip1(n5639), .ip2(n5638), .op(n5640) );
  ab_or_c_or_d U6248 ( .ip1(n5643), .ip2(n5642), .ip3(n5641), .ip4(n5640), 
        .op(n5644) );
  nand2_1 U6249 ( .ip1(n5645), .ip2(n5644), .op(n6233) );
  fulladder U6250 ( .a(n5648), .b(n5647), .ci(n5646), .co(n6232), .s(n5637) );
  inv_1 U6251 ( .ip(m1Inputs[5]), .op(n10166) );
  nor2_1 U6252 ( .ip1(n13570), .ip2(n10166), .op(n5650) );
  nand2_1 U6253 ( .ip1(n4672), .ip2(m1Inputs[4]), .op(n5649) );
  xor2_1 U6254 ( .ip1(n5650), .ip2(n5649), .op(n5699) );
  nand2_1 U6255 ( .ip1(n13803), .ip2(m1Inputs[5]), .op(n5685) );
  inv_1 U6256 ( .ip(m1Inputs[2]), .op(n10150) );
  nor4_1 U6257 ( .ip1(n10476), .ip2(n13082), .ip3(n10150), .ip4(n10166), .op(
        n5654) );
  or2_1 U6258 ( .ip1(n5685), .ip2(n5654), .op(n5653) );
  nand2_1 U6259 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[2]), .op(n5651)
         );
  or2_1 U6260 ( .ip1(n5651), .ip2(n5654), .op(n5652) );
  nand2_1 U6261 ( .ip1(n5653), .ip2(n5652), .op(n5719) );
  or2_1 U6262 ( .ip1(n5719), .ip2(n5654), .op(n5656) );
  inv_1 U6263 ( .ip(m1Inputs[0]), .op(n10127) );
  nor2_1 U6264 ( .ip1(n10127), .ip2(n12746), .op(n5718) );
  or2_1 U6265 ( .ip1(n5718), .ip2(n5654), .op(n5655) );
  nand2_1 U6266 ( .ip1(n5656), .ip2(n5655), .op(n5698) );
  inv_1 U6267 ( .ip(m1Inputs[1]), .op(n10160) );
  nor2_1 U6268 ( .ip1(n10160), .ip2(n12746), .op(n5680) );
  inv_1 U6269 ( .ip(m1Inputs[6]), .op(n9908) );
  nor2_1 U6270 ( .ip1(n10476), .ip2(n9908), .op(n6040) );
  nor2_1 U6271 ( .ip1(n10127), .ip2(n14836), .op(n5679) );
  inv_1 U6272 ( .ip(n5657), .op(n5697) );
  nor3_1 U6273 ( .ip1(n5707), .ip2(n9908), .ip3(n9047), .op(n6078) );
  nand2_1 U6274 ( .ip1(m1Inputs[3]), .ip2(\STAGE_1/weightReg [4]), .op(n5681)
         );
  inv_1 U6275 ( .ip(m1Inputs[3]), .op(n10003) );
  nand2_1 U6276 ( .ip1(m1Inputs[2]), .ip2(n11974), .op(n5702) );
  nor3_1 U6277 ( .ip1(n10003), .ip2(n5702), .ip3(n4624), .op(n5661) );
  or2_1 U6278 ( .ip1(n5681), .ip2(n5661), .op(n5660) );
  nand2_1 U6279 ( .ip1(m1Inputs[2]), .ip2(n12699), .op(n5658) );
  or2_1 U6280 ( .ip1(n5658), .ip2(n5661), .op(n5659) );
  nand2_1 U6281 ( .ip1(n5660), .ip2(n5659), .op(n5672) );
  or2_1 U6282 ( .ip1(n5672), .ip2(n5661), .op(n5663) );
  nor2_1 U6283 ( .ip1(n10127), .ip2(n14384), .op(n5671) );
  or2_1 U6284 ( .ip1(n5671), .ip2(n5661), .op(n5662) );
  nand2_1 U6285 ( .ip1(n5663), .ip2(n5662), .op(n6047) );
  nand2_1 U6286 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[7]), .op(n6090)
         );
  inv_1 U6287 ( .ip(m1Inputs[4]), .op(n10088) );
  nor2_1 U6288 ( .ip1(n13646), .ip2(n10088), .op(n5729) );
  and3_1 U6289 ( .ip1(n9733), .ip2(m1Inputs[7]), .ip3(n5729), .op(n5667) );
  or2_1 U6290 ( .ip1(n6090), .ip2(n5667), .op(n5666) );
  nand2_1 U6291 ( .ip1(n9733), .ip2(m1Inputs[4]), .op(n5664) );
  or2_1 U6292 ( .ip1(n5664), .ip2(n5667), .op(n5665) );
  nand2_1 U6293 ( .ip1(n5666), .ip2(n5665), .op(n5677) );
  or2_1 U6294 ( .ip1(n5677), .ip2(n5667), .op(n5669) );
  nor2_1 U6295 ( .ip1(n6745), .ip2(n10166), .op(n5676) );
  or2_1 U6296 ( .ip1(n5676), .ip2(n5667), .op(n5668) );
  nand2_1 U6297 ( .ip1(n5669), .ip2(n5668), .op(n6046) );
  nand2_1 U6298 ( .ip1(m1Inputs[2]), .ip2(n12981), .op(n6045) );
  inv_1 U6299 ( .ip(n5670), .op(n6075) );
  xnor2_1 U6300 ( .ip1(n5672), .ip2(n5671), .op(n5705) );
  nand4_1 U6301 ( .ip1(n4619), .ip2(\STAGE_1/weightReg [1]), .ip3(m1Inputs[3]), 
        .ip4(m1Inputs[4]), .op(n5691) );
  nor2_1 U6302 ( .ip1(n13082), .ip2(n5691), .op(n5675) );
  nand2_1 U6303 ( .ip1(n5691), .ip2(m1Inputs[3]), .op(n5673) );
  mux2_1 U6304 ( .ip1(n5691), .ip2(n5673), .s(n9733), .op(n5701) );
  nor2_1 U6305 ( .ip1(n5702), .ip2(n5701), .op(n5674) );
  nor2_1 U6306 ( .ip1(n5675), .ip2(n5674), .op(n5704) );
  xnor2_1 U6307 ( .ip1(n5677), .ip2(n5676), .op(n5703) );
  inv_1 U6308 ( .ip(n5678), .op(n6074) );
  nor2_1 U6309 ( .ip1(n10160), .ip2(n14289), .op(n5713) );
  nor4_1 U6310 ( .ip1(n6745), .ip2(n9047), .ip3(n10088), .ip4(n10166), .op(
        n5712) );
  fulladder U6311 ( .a(n5680), .b(n6040), .ci(n5679), .co(n5711), .s(n5657) );
  nand2_1 U6312 ( .ip1(m1Inputs[3]), .ip2(\STAGE_1/weightReg [5]), .op(n5682)
         );
  nor3_1 U6313 ( .ip1(n10088), .ip2(n12746), .ip3(n5681), .op(n6061) );
  or2_1 U6314 ( .ip1(n5682), .ip2(n6061), .op(n5684) );
  nand2_1 U6315 ( .ip1(n13637), .ip2(m1Inputs[4]), .op(n6036) );
  or2_1 U6316 ( .ip1(n6036), .ip2(n6061), .op(n5683) );
  nand2_1 U6317 ( .ip1(n5684), .ip2(n5683), .op(n6060) );
  nor2_1 U6318 ( .ip1(n10160), .ip2(n14384), .op(n6062) );
  xor2_1 U6319 ( .ip1(n6060), .ip2(n6062), .op(n6072) );
  nand2_1 U6320 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[5]), .op(n5686)
         );
  inv_1 U6321 ( .ip(m1Inputs[8]), .op(n10072) );
  nor3_1 U6322 ( .ip1(n13082), .ip2(n10072), .ip3(n5685), .op(n6056) );
  or2_1 U6323 ( .ip1(n5686), .ip2(n6056), .op(n5688) );
  nand2_1 U6324 ( .ip1(n13803), .ip2(m1Inputs[8]), .op(n6143) );
  or2_1 U6325 ( .ip1(n6143), .ip2(n6056), .op(n5687) );
  nand2_1 U6326 ( .ip1(n5688), .ip2(n5687), .op(n6055) );
  nor2_1 U6327 ( .ip1(n10127), .ip2(n6503), .op(n6057) );
  xor2_1 U6328 ( .ip1(n6055), .ip2(n6057), .op(n6071) );
  nand2_1 U6329 ( .ip1(m1Inputs[6]), .ip2(n4619), .op(n5689) );
  nand2_1 U6330 ( .ip1(n10507), .ip2(m1Inputs[7]), .op(n6065) );
  nand2_1 U6331 ( .ip1(n5689), .ip2(n6065), .op(n5690) );
  nand4_1 U6332 ( .ip1(n4619), .ip2(\STAGE_1/weightReg [1]), .ip3(m1Inputs[7]), 
        .ip4(m1Inputs[6]), .op(n6049) );
  nand2_1 U6333 ( .ip1(n5690), .ip2(n6049), .op(n6051) );
  nand2_1 U6334 ( .ip1(column[0]), .ip2(n13859), .op(n6050) );
  xor2_1 U6335 ( .ip1(n6051), .ip2(n6050), .op(n6070) );
  nand2_1 U6336 ( .ip1(n10507), .ip2(m1Inputs[2]), .op(n5742) );
  nor3_1 U6337 ( .ip1(n10555), .ip2(n10003), .ip3(n5742), .op(n5726) );
  inv_1 U6338 ( .ip(n5691), .op(n5696) );
  nor2_1 U6339 ( .ip1(n6745), .ip2(n10003), .op(n5692) );
  or2_1 U6340 ( .ip1(m1Inputs[4]), .ip2(n5692), .op(n5694) );
  or2_1 U6341 ( .ip1(n10507), .ip2(n5692), .op(n5693) );
  nand2_1 U6342 ( .ip1(n5694), .ip2(n5693), .op(n5695) );
  nor2_1 U6343 ( .ip1(n5696), .ip2(n5695), .op(n5721) );
  nor2_1 U6344 ( .ip1(n10160), .ip2(n14783), .op(n5720) );
  fulladder U6345 ( .a(n5699), .b(n5698), .ci(n5697), .co(n5707), .s(n5700) );
  inv_1 U6346 ( .ip(n5700), .op(n5715) );
  xor2_1 U6347 ( .ip1(n5702), .ip2(n5701), .op(n5714) );
  fulladder U6348 ( .a(n5705), .b(n5704), .ci(n5703), .co(n5678), .s(n5706) );
  inv_1 U6349 ( .ip(n5706), .op(n5778) );
  or2_1 U6350 ( .ip1(n5707), .ip2(n6078), .op(n5710) );
  nand2_1 U6351 ( .ip1(n13707), .ip2(m1Inputs[6]), .op(n5708) );
  or2_1 U6352 ( .ip1(n5708), .ip2(n6078), .op(n5709) );
  nand2_1 U6353 ( .ip1(n5710), .ip2(n5709), .op(n5777) );
  fulladder U6354 ( .a(n5713), .b(n5712), .ci(n5711), .co(n6073), .s(n5776) );
  nand2_1 U6355 ( .ip1(n5767), .ip2(n5766), .op(n5775) );
  fulladder U6356 ( .a(n5716), .b(n5715), .ci(n5714), .co(n5767), .s(n5717) );
  inv_1 U6357 ( .ip(n5717), .op(n5773) );
  xor2_1 U6358 ( .ip1(n5719), .ip2(n5718), .op(n5759) );
  fulladder U6359 ( .a(n5726), .b(n5721), .ci(n5720), .co(n5716), .s(n5758) );
  nor2_1 U6360 ( .ip1(n10127), .ip2(n14783), .op(n5728) );
  nor2_1 U6361 ( .ip1(n13801), .ip2(n10160), .op(n5727) );
  nor4_1 U6362 ( .ip1(n9047), .ip2(n13801), .ip3(n10127), .ip4(n10150), .op(
        n5743) );
  nor2_1 U6363 ( .ip1(n13570), .ip2(n10003), .op(n5722) );
  or2_1 U6364 ( .ip1(m1Inputs[2]), .ip2(n5722), .op(n5724) );
  or2_1 U6365 ( .ip1(n4619), .ip2(n5722), .op(n5723) );
  nand2_1 U6366 ( .ip1(n5724), .ip2(n5723), .op(n5725) );
  nor2_1 U6367 ( .ip1(n5726), .ip2(n5725), .op(n5731) );
  fulladder U6368 ( .a(n5729), .b(n5728), .ci(n5727), .co(n5757), .s(n5730) );
  fulladder U6369 ( .a(n5743), .b(n5731), .ci(n5730), .co(n5760), .s(n5750) );
  nand4_1 U6370 ( .ip1(n4619), .ip2(\STAGE_1/weightReg [1]), .ip3(m1Inputs[0]), 
        .ip4(m1Inputs[1]), .op(n5734) );
  nand2_1 U6371 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[3]), .op(n5733)
         );
  and2_1 U6372 ( .ip1(n5734), .ip2(n5733), .op(n5732) );
  nor3_1 U6373 ( .ip1(n5732), .ip2(n10160), .ip3(n6745), .op(n5749) );
  nand2_1 U6374 ( .ip1(n5750), .ip2(n5749), .op(n5756) );
  xor2_1 U6375 ( .ip1(n5734), .ip2(n5733), .op(n5736) );
  nand2_1 U6376 ( .ip1(n4672), .ip2(m1Inputs[1]), .op(n5735) );
  xor2_1 U6377 ( .ip1(n5736), .ip2(n5735), .op(n5754) );
  nand2_1 U6378 ( .ip1(n4619), .ip2(m1Inputs[0]), .op(n5738) );
  nand2_1 U6379 ( .ip1(n13707), .ip2(m1Inputs[1]), .op(n5737) );
  not_ab_or_c_or_d U6380 ( .ip1(n5738), .ip2(n5737), .ip3(n13646), .ip4(n10150), .op(n5741) );
  nor4_1 U6381 ( .ip1(n13570), .ip2(n5739), .ip3(n10127), .ip4(n10160), .op(
        n5740) );
  nor2_1 U6382 ( .ip1(n5741), .ip2(n5740), .op(n5753) );
  or2_1 U6383 ( .ip1(n5742), .ip2(n5743), .op(n5746) );
  nand2_1 U6384 ( .ip1(n9733), .ip2(m1Inputs[0]), .op(n5744) );
  or2_1 U6385 ( .ip1(n5744), .ip2(n5743), .op(n5745) );
  nand2_1 U6386 ( .ip1(n5746), .ip2(n5745), .op(n5748) );
  nor2_1 U6387 ( .ip1(n5753), .ip2(n5754), .op(n5747) );
  nor2_1 U6388 ( .ip1(n5748), .ip2(n5747), .op(n5752) );
  nor2_1 U6389 ( .ip1(n5750), .ip2(n5749), .op(n5751) );
  ab_or_c_or_d U6390 ( .ip1(n5754), .ip2(n5753), .ip3(n5752), .ip4(n5751), 
        .op(n5755) );
  nand2_1 U6391 ( .ip1(n5756), .ip2(n5755), .op(n5762) );
  nand2_1 U6392 ( .ip1(n5760), .ip2(n5762), .op(n5765) );
  fulladder U6393 ( .a(n5759), .b(n5758), .ci(n5757), .co(n5769), .s(n5761) );
  nand2_1 U6394 ( .ip1(n5760), .ip2(n5761), .op(n5764) );
  nand2_1 U6395 ( .ip1(n5762), .ip2(n5761), .op(n5763) );
  nand3_1 U6396 ( .ip1(n5765), .ip2(n5764), .ip3(n5763), .op(n5768) );
  nand2_1 U6397 ( .ip1(n5769), .ip2(n5768), .op(n5772) );
  nor2_1 U6398 ( .ip1(n5767), .ip2(n5766), .op(n5771) );
  nor2_1 U6399 ( .ip1(n5769), .ip2(n5768), .op(n5770) );
  ab_or_c_or_d U6400 ( .ip1(n5773), .ip2(n5772), .ip3(n5771), .ip4(n5770), 
        .op(n5774) );
  nand2_1 U6401 ( .ip1(n5775), .ip2(n5774), .op(n6080) );
  fulladder U6402 ( .a(n5778), .b(n5777), .ci(n5776), .co(n6079), .s(n5766) );
  inv_1 U6403 ( .ip(m1Inputs[69]), .op(n12999) );
  nor2_1 U6404 ( .ip1(n13646), .ip2(n12999), .op(n5838) );
  inv_1 U6405 ( .ip(m1Inputs[66]), .op(n13050) );
  nor2_1 U6406 ( .ip1(n13801), .ip2(n13050), .op(n5837) );
  inv_1 U6407 ( .ip(m1Inputs[64]), .op(n12964) );
  nor2_1 U6408 ( .ip1(n12964), .ip2(n12746), .op(n5836) );
  nand2_1 U6409 ( .ip1(n4672), .ip2(m1Inputs[68]), .op(n5779) );
  inv_1 U6410 ( .ip(m1Inputs[68]), .op(n12925) );
  nor4_1 U6411 ( .ip1(n6745), .ip2(n9047), .ip3(n12925), .ip4(n12999), .op(
        n5823) );
  or2_1 U6412 ( .ip1(n5779), .ip2(n5823), .op(n5782) );
  nand2_1 U6413 ( .ip1(n13707), .ip2(m1Inputs[69]), .op(n5780) );
  or2_1 U6414 ( .ip1(n5780), .ip2(n5823), .op(n5781) );
  nand2_1 U6415 ( .ip1(n5782), .ip2(n5781), .op(n5832) );
  inv_1 U6416 ( .ip(m1Inputs[65]), .op(n13076) );
  nor2_1 U6417 ( .ip1(n13076), .ip2(n13835), .op(n5805) );
  inv_1 U6418 ( .ip(m1Inputs[70]), .op(n13045) );
  nor2_1 U6419 ( .ip1(n13646), .ip2(n13045), .op(n5944) );
  nor2_1 U6420 ( .ip1(n12964), .ip2(n14289), .op(n5804) );
  and3_1 U6421 ( .ip1(n10507), .ip2(m1Inputs[70]), .ip3(n5819), .op(n5982) );
  nand2_1 U6422 ( .ip1(m1Inputs[67]), .ip2(n13637), .op(n5806) );
  inv_1 U6423 ( .ip(m1Inputs[67]), .op(n12845) );
  nand2_1 U6424 ( .ip1(m1Inputs[66]), .ip2(n13637), .op(n5835) );
  nor3_1 U6425 ( .ip1(n12845), .ip2(n5835), .ip3(n4624), .op(n5786) );
  or2_1 U6426 ( .ip1(n5806), .ip2(n5786), .op(n5785) );
  nand2_1 U6427 ( .ip1(m1Inputs[66]), .ip2(n14369), .op(n5783) );
  or2_1 U6428 ( .ip1(n5783), .ip2(n5786), .op(n5784) );
  nand2_1 U6429 ( .ip1(n5785), .ip2(n5784), .op(n5797) );
  or2_1 U6430 ( .ip1(n5797), .ip2(n5786), .op(n5788) );
  nor2_1 U6431 ( .ip1(n12964), .ip2(n14384), .op(n5796) );
  or2_1 U6432 ( .ip1(n5796), .ip2(n5786), .op(n5787) );
  nand2_1 U6433 ( .ip1(n5788), .ip2(n5787), .op(n5951) );
  nand2_1 U6434 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[71]), .op(n5986)
         );
  nor2_1 U6435 ( .ip1(n13646), .ip2(n12925), .op(n5852) );
  and3_1 U6436 ( .ip1(n12578), .ip2(m1Inputs[71]), .ip3(n5852), .op(n5792) );
  or2_1 U6437 ( .ip1(n5986), .ip2(n5792), .op(n5791) );
  nand2_1 U6438 ( .ip1(n13614), .ip2(m1Inputs[68]), .op(n5789) );
  or2_1 U6439 ( .ip1(n5789), .ip2(n5792), .op(n5790) );
  nand2_1 U6440 ( .ip1(n5791), .ip2(n5790), .op(n5802) );
  or2_1 U6441 ( .ip1(n5802), .ip2(n5792), .op(n5794) );
  nor2_1 U6442 ( .ip1(n13854), .ip2(n12999), .op(n5801) );
  or2_1 U6443 ( .ip1(n5801), .ip2(n5792), .op(n5793) );
  nand2_1 U6444 ( .ip1(n5794), .ip2(n5793), .op(n5950) );
  nand2_1 U6445 ( .ip1(m1Inputs[66]), .ip2(n12981), .op(n5949) );
  inv_1 U6446 ( .ip(n5795), .op(n5979) );
  xnor2_1 U6447 ( .ip1(n5797), .ip2(n5796), .op(n5817) );
  nand4_1 U6448 ( .ip1(n4672), .ip2(n10507), .ip3(m1Inputs[67]), .ip4(
        m1Inputs[68]), .op(n5825) );
  nor2_1 U6449 ( .ip1(n13801), .ip2(n5825), .op(n5800) );
  nand2_1 U6450 ( .ip1(n5825), .ip2(m1Inputs[67]), .op(n5798) );
  mux2_1 U6451 ( .ip1(n5825), .ip2(n5798), .s(n9733), .op(n5834) );
  nor2_1 U6452 ( .ip1(n5835), .ip2(n5834), .op(n5799) );
  nor2_1 U6453 ( .ip1(n5800), .ip2(n5799), .op(n5816) );
  xnor2_1 U6454 ( .ip1(n5802), .ip2(n5801), .op(n5815) );
  inv_1 U6455 ( .ip(n5803), .op(n5978) );
  nor2_1 U6456 ( .ip1(n13076), .ip2(n14289), .op(n5824) );
  fulladder U6457 ( .a(n5805), .b(n5944), .ci(n5804), .co(n5822), .s(n5831) );
  nand2_1 U6458 ( .ip1(m1Inputs[67]), .ip2(n14369), .op(n5807) );
  nor3_1 U6459 ( .ip1(n12925), .ip2(n13835), .ip3(n5806), .op(n5965) );
  or2_1 U6460 ( .ip1(n5807), .ip2(n5965), .op(n5809) );
  nand2_1 U6461 ( .ip1(n13637), .ip2(m1Inputs[68]), .op(n5940) );
  or2_1 U6462 ( .ip1(n5940), .ip2(n5965), .op(n5808) );
  nand2_1 U6463 ( .ip1(n5809), .ip2(n5808), .op(n5964) );
  nor2_1 U6464 ( .ip1(n13076), .ip2(n14368), .op(n5966) );
  xor2_1 U6465 ( .ip1(n5964), .ip2(n5966), .op(n5976) );
  and3_1 U6466 ( .ip1(n12578), .ip2(m1Inputs[72]), .ip3(n5838), .op(n5960) );
  inv_1 U6467 ( .ip(m1Inputs[72]), .op(n13071) );
  nor2_1 U6468 ( .ip1(n13646), .ip2(n13071), .op(n12577) );
  or2_1 U6469 ( .ip1(m1Inputs[69]), .ip2(n12577), .op(n5811) );
  or2_1 U6470 ( .ip1(n9733), .ip2(n12577), .op(n5810) );
  nand2_1 U6471 ( .ip1(n5811), .ip2(n5810), .op(n5812) );
  nor2_1 U6472 ( .ip1(n5960), .ip2(n5812), .op(n5959) );
  nor2_1 U6473 ( .ip1(n12964), .ip2(n6504), .op(n5961) );
  xor2_1 U6474 ( .ip1(n5959), .ip2(n5961), .op(n5975) );
  nand2_1 U6475 ( .ip1(m1Inputs[70]), .ip2(n4672), .op(n5813) );
  nand2_1 U6476 ( .ip1(n13707), .ip2(m1Inputs[71]), .op(n5969) );
  nand2_1 U6477 ( .ip1(n5813), .ip2(n5969), .op(n5814) );
  nand4_1 U6478 ( .ip1(n4619), .ip2(n10507), .ip3(m1Inputs[71]), .ip4(
        m1Inputs[70]), .op(n5953) );
  nand2_1 U6479 ( .ip1(n5814), .ip2(n5953), .op(n5955) );
  nand2_1 U6480 ( .ip1(column[64]), .ip2(n13039), .op(n5954) );
  xor2_1 U6481 ( .ip1(n5955), .ip2(n5954), .op(n5974) );
  fulladder U6482 ( .a(n5817), .b(n5816), .ci(n5815), .co(n5803), .s(n5818) );
  inv_1 U6483 ( .ip(n5818), .op(n5902) );
  nor2_1 U6484 ( .ip1(n9047), .ip2(n13045), .op(n5820) );
  nor2_1 U6485 ( .ip1(n5820), .ip2(n5819), .op(n5821) );
  nor2_1 U6486 ( .ip1(n5982), .ip2(n5821), .op(n5901) );
  fulladder U6487 ( .a(n5824), .b(n5823), .ci(n5822), .co(n5977), .s(n5900) );
  nand2_1 U6488 ( .ip1(n13707), .ip2(m1Inputs[66]), .op(n5855) );
  nor3_1 U6489 ( .ip1(n13854), .ip2(n12845), .ip3(n5855), .op(n5849) );
  inv_1 U6490 ( .ip(n5825), .op(n5830) );
  nor2_1 U6491 ( .ip1(n13854), .ip2(n12845), .op(n5826) );
  or2_1 U6492 ( .ip1(m1Inputs[68]), .ip2(n5826), .op(n5828) );
  or2_1 U6493 ( .ip1(n10507), .ip2(n5826), .op(n5827) );
  nand2_1 U6494 ( .ip1(n5828), .ip2(n5827), .op(n5829) );
  nor2_1 U6495 ( .ip1(n5830), .ip2(n5829), .op(n5840) );
  nor2_1 U6496 ( .ip1(n13076), .ip2(n14783), .op(n5839) );
  fulladder U6497 ( .a(n5833), .b(n5832), .ci(n5831), .co(n5819), .s(n5843) );
  xor2_1 U6498 ( .ip1(n5835), .ip2(n5834), .op(n5842) );
  nand2_1 U6499 ( .ip1(n5891), .ip2(n5890), .op(n5899) );
  fulladder U6500 ( .a(n5838), .b(n5837), .ci(n5836), .co(n5833), .s(n5880) );
  fulladder U6501 ( .a(n5849), .b(n5840), .ci(n5839), .co(n5844), .s(n5879) );
  nor2_1 U6502 ( .ip1(n12964), .ip2(n14783), .op(n5851) );
  nor2_1 U6503 ( .ip1(n13801), .ip2(n13076), .op(n5850) );
  inv_1 U6504 ( .ip(n5841), .op(n5897) );
  fulladder U6505 ( .a(n5844), .b(n5843), .ci(n5842), .co(n5890), .s(n5893) );
  nor4_1 U6506 ( .ip1(n13570), .ip2(n13082), .ip3(n12964), .ip4(n13050), .op(
        n5883) );
  nor2_1 U6507 ( .ip1(n9047), .ip2(n12845), .op(n5845) );
  or2_1 U6508 ( .ip1(m1Inputs[66]), .ip2(n5845), .op(n5847) );
  or2_1 U6509 ( .ip1(n4672), .ip2(n5845), .op(n5846) );
  nand2_1 U6510 ( .ip1(n5847), .ip2(n5846), .op(n5848) );
  nor2_1 U6511 ( .ip1(n5849), .ip2(n5848), .op(n5882) );
  fulladder U6512 ( .a(n5852), .b(n5851), .ci(n5850), .co(n5878), .s(n5881) );
  nand4_1 U6513 ( .ip1(n4672), .ip2(n10507), .ip3(m1Inputs[65]), .ip4(
        m1Inputs[64]), .op(n5854) );
  not_ab_or_c_or_d U6514 ( .ip1(n13707), .ip2(m1Inputs[64]), .ip3(n10555), 
        .ip4(n13076), .op(n5865) );
  nand3_1 U6515 ( .ip1(\STAGE_1/weightReg [0]), .ip2(n5865), .ip3(m1Inputs[67]), .op(n5853) );
  nand2_1 U6516 ( .ip1(n5854), .ip2(n5853), .op(n5874) );
  nand2_1 U6517 ( .ip1(n5872), .ip2(n5874), .op(n5877) );
  or2_1 U6518 ( .ip1(n5855), .ip2(n5883), .op(n5858) );
  nand2_1 U6519 ( .ip1(n13614), .ip2(m1Inputs[64]), .op(n5856) );
  or2_1 U6520 ( .ip1(n5856), .ip2(n5883), .op(n5857) );
  nand2_1 U6521 ( .ip1(n5858), .ip2(n5857), .op(n5866) );
  nand2_1 U6522 ( .ip1(n13707), .ip2(m1Inputs[65]), .op(n5863) );
  nand2_1 U6523 ( .ip1(n5056), .ip2(m1Inputs[64]), .op(n5862) );
  or2_1 U6524 ( .ip1(m1Inputs[64]), .ip2(m1Inputs[66]), .op(n5860) );
  or2_1 U6525 ( .ip1(n13854), .ip2(m1Inputs[66]), .op(n5859) );
  nand2_1 U6526 ( .ip1(n5860), .ip2(n5859), .op(n5861) );
  not_ab_or_c_or_d U6527 ( .ip1(n5863), .ip2(n5862), .ip3(n5861), .ip4(n10476), 
        .op(n5868) );
  nand2_1 U6528 ( .ip1(n5866), .ip2(n5868), .op(n5871) );
  nor2_1 U6529 ( .ip1(n13646), .ip2(n12845), .op(n5864) );
  xor2_1 U6530 ( .ip1(n5865), .ip2(n5864), .op(n5867) );
  nand2_1 U6531 ( .ip1(n5866), .ip2(n5867), .op(n5870) );
  nand2_1 U6532 ( .ip1(n5868), .ip2(n5867), .op(n5869) );
  nand3_1 U6533 ( .ip1(n5871), .ip2(n5870), .ip3(n5869), .op(n5873) );
  nand2_1 U6534 ( .ip1(n5872), .ip2(n5873), .op(n5876) );
  nand2_1 U6535 ( .ip1(n5874), .ip2(n5873), .op(n5875) );
  nand3_1 U6536 ( .ip1(n5877), .ip2(n5876), .ip3(n5875), .op(n5884) );
  fulladder U6537 ( .a(n5880), .b(n5879), .ci(n5878), .co(n5841), .s(n5886) );
  nand2_1 U6538 ( .ip1(n5884), .ip2(n5886), .op(n5889) );
  fulladder U6539 ( .a(n5883), .b(n5882), .ci(n5881), .co(n5885), .s(n5872) );
  nand2_1 U6540 ( .ip1(n5884), .ip2(n5885), .op(n5888) );
  nand2_1 U6541 ( .ip1(n5886), .ip2(n5885), .op(n5887) );
  nand3_1 U6542 ( .ip1(n5889), .ip2(n5888), .ip3(n5887), .op(n5892) );
  nand2_1 U6543 ( .ip1(n5893), .ip2(n5892), .op(n5896) );
  nor2_1 U6544 ( .ip1(n5891), .ip2(n5890), .op(n5895) );
  nor2_1 U6545 ( .ip1(n5893), .ip2(n5892), .op(n5894) );
  ab_or_c_or_d U6546 ( .ip1(n5897), .ip2(n5896), .ip3(n5895), .ip4(n5894), 
        .op(n5898) );
  nand2_1 U6547 ( .ip1(n5899), .ip2(n5898), .op(n5984) );
  fulladder U6548 ( .a(n5902), .b(n5901), .ci(n5900), .co(n5983), .s(n5891) );
  nand2_1 U6549 ( .ip1(m1Inputs[20]), .ip2(n12699), .op(n5904) );
  nor3_1 U6550 ( .ip1(n13835), .ip2(n10866), .ip3(n5903), .op(n6640) );
  or2_1 U6551 ( .ip1(n5904), .ip2(n6640), .op(n5906) );
  nand2_1 U6552 ( .ip1(n13637), .ip2(m1Inputs[21]), .op(n6610) );
  or2_1 U6553 ( .ip1(n6610), .ip2(n6640), .op(n5905) );
  nand2_1 U6554 ( .ip1(n5906), .ip2(n5905), .op(n6639) );
  nor2_1 U6555 ( .ip1(n10472), .ip2(n6503), .op(n6641) );
  xnor2_1 U6556 ( .ip1(n6639), .ip2(n6641), .op(n6695) );
  and3_1 U6557 ( .ip1(n12578), .ip2(m1Inputs[25]), .ip3(n5907), .op(n6636) );
  inv_1 U6558 ( .ip(m1Inputs[25]), .op(n10753) );
  nor2_1 U6559 ( .ip1(n13646), .ip2(n10753), .op(n5908) );
  or2_1 U6560 ( .ip1(m1Inputs[22]), .ip2(n5908), .op(n5910) );
  or2_1 U6561 ( .ip1(n9733), .ip2(n5908), .op(n5909) );
  nand2_1 U6562 ( .ip1(n5910), .ip2(n5909), .op(n6634) );
  nor2_1 U6563 ( .ip1(n6636), .ip2(n6634), .op(n5911) );
  inv_1 U6564 ( .ip(n13766), .op(n14994) );
  nand2_1 U6565 ( .ip1(m1Inputs[16]), .ip2(n14994), .op(n6633) );
  xor2_1 U6566 ( .ip1(n5911), .ip2(n6633), .op(n6694) );
  fulladder U6567 ( .a(n5914), .b(n5913), .ci(n5912), .co(n6693), .s(n5287) );
  inv_1 U6568 ( .ip(n5915), .op(n6719) );
  nor2_1 U6569 ( .ip1(n10585), .ip2(n12156), .op(n6676) );
  nor2_1 U6570 ( .ip1(n10461), .ip2(n14289), .op(n6675) );
  buf_1 U6571 ( .ip(n14768), .op(n15042) );
  nand3_1 U6572 ( .ip1(column[16]), .ip2(n15042), .ip3(n5916), .op(n5917) );
  nand2_1 U6573 ( .ip1(n5918), .ip2(n5917), .op(n6674) );
  nand2_1 U6574 ( .ip1(n10507), .ip2(m1Inputs[24]), .op(n6573) );
  inv_1 U6575 ( .ip(m1Inputs[24]), .op(n10812) );
  nor4_1 U6576 ( .ip1(n6745), .ip2(n13570), .ip3(n10812), .ip4(n10734), .op(
        n6646) );
  or2_1 U6577 ( .ip1(n6573), .ip2(n6646), .op(n5921) );
  nand2_1 U6578 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[23]), .op(n5919)
         );
  or2_1 U6579 ( .ip1(n5919), .ip2(n6646), .op(n5920) );
  nand2_1 U6580 ( .ip1(n5921), .ip2(n5920), .op(n6644) );
  nand2_1 U6581 ( .ip1(column[17]), .ip2(n13859), .op(n6645) );
  xor2_1 U6582 ( .ip1(n6644), .ip2(n6645), .op(n6672) );
  inv_1 U6583 ( .ip(n5922), .op(n5924) );
  nor2_1 U6584 ( .ip1(n5924), .ip2(n5923), .op(n6671) );
  nor2_1 U6585 ( .ip1(n5926), .ip2(n5925), .op(n6670) );
  inv_1 U6586 ( .ip(n5927), .op(n6709) );
  fulladder U6587 ( .a(n5930), .b(n5929), .ci(n5928), .co(n6708), .s(n5934) );
  fulladder U6588 ( .a(n5933), .b(n5932), .ci(n5931), .co(n6717), .s(n5935) );
  fulladder U6589 ( .a(n5936), .b(n5935), .ci(n5934), .co(n6715), .s(n5939) );
  fulladder U6590 ( .a(n5939), .b(n5938), .ci(n5937), .co(n6714), .s(
        \STAGE_1/M2/sum [0]) );
  nand2_1 U6591 ( .ip1(m1Inputs[68]), .ip2(n14369), .op(n5941) );
  nor3_1 U6592 ( .ip1(n4624), .ip2(n12999), .ip3(n5940), .op(n5997) );
  or2_1 U6593 ( .ip1(n5941), .ip2(n5997), .op(n5943) );
  nand2_1 U6594 ( .ip1(n13637), .ip2(m1Inputs[69]), .op(n6019) );
  or2_1 U6595 ( .ip1(n6019), .ip2(n5997), .op(n5942) );
  nand2_1 U6596 ( .ip1(n5943), .ip2(n5942), .op(n5996) );
  nor2_1 U6597 ( .ip1(n13076), .ip2(n6504), .op(n5998) );
  xnor2_1 U6598 ( .ip1(n5996), .ip2(n5998), .op(n6025) );
  and3_1 U6599 ( .ip1(n12578), .ip2(m1Inputs[73]), .ip3(n5944), .op(n6018) );
  inv_1 U6600 ( .ip(m1Inputs[73]), .op(n13081) );
  nor2_1 U6601 ( .ip1(n13646), .ip2(n13081), .op(n5945) );
  or2_1 U6602 ( .ip1(m1Inputs[70]), .ip2(n5945), .op(n5947) );
  or2_1 U6603 ( .ip1(n9733), .ip2(n5945), .op(n5946) );
  nand2_1 U6604 ( .ip1(n5947), .ip2(n5946), .op(n6016) );
  nor2_1 U6605 ( .ip1(n6018), .ip2(n6016), .op(n5948) );
  nand2_1 U6606 ( .ip1(m1Inputs[64]), .ip2(\STAGE_1/weightReg [9]), .op(n6015)
         );
  xor2_1 U6607 ( .ip1(n5948), .ip2(n6015), .op(n6024) );
  fulladder U6608 ( .a(n5951), .b(n5950), .ci(n5949), .co(n6023), .s(n5795) );
  inv_1 U6609 ( .ip(n5952), .op(n6035) );
  inv_1 U6610 ( .ip(n5953), .op(n5957) );
  nor2_1 U6611 ( .ip1(n5955), .ip2(n5954), .op(n5956) );
  nor2_1 U6612 ( .ip1(n5957), .ip2(n5956), .op(n5994) );
  nand2_1 U6613 ( .ip1(m1Inputs[67]), .ip2(n12981), .op(n6011) );
  nand2_1 U6614 ( .ip1(m1Inputs[66]), .ip2(n4627), .op(n5993) );
  inv_1 U6615 ( .ip(n5958), .op(n6029) );
  or2_1 U6616 ( .ip1(n5959), .ip2(n5960), .op(n5963) );
  or2_1 U6617 ( .ip1(n5961), .ip2(n5960), .op(n5962) );
  nand2_1 U6618 ( .ip1(n5963), .ip2(n5962), .op(n5992) );
  or2_1 U6619 ( .ip1(n5964), .ip2(n5965), .op(n5968) );
  or2_1 U6620 ( .ip1(n5966), .ip2(n5965), .op(n5967) );
  nand2_1 U6621 ( .ip1(n5968), .ip2(n5967), .op(n5991) );
  nand2_1 U6622 ( .ip1(n4672), .ip2(m1Inputs[71]), .op(n5970) );
  nor3_1 U6623 ( .ip1(n13854), .ip2(n13071), .ip3(n5969), .op(n6003) );
  or2_1 U6624 ( .ip1(n5970), .ip2(n6003), .op(n5972) );
  nand2_1 U6625 ( .ip1(n13707), .ip2(m1Inputs[72]), .op(n6007) );
  or2_1 U6626 ( .ip1(n6007), .ip2(n6003), .op(n5971) );
  nand2_1 U6627 ( .ip1(n5972), .ip2(n5971), .op(n6001) );
  nand2_1 U6628 ( .ip1(column[65]), .ip2(n15042), .op(n6002) );
  xor2_1 U6629 ( .ip1(n6001), .ip2(n6002), .op(n5990) );
  inv_1 U6630 ( .ip(n5973), .op(n6028) );
  fulladder U6631 ( .a(n5976), .b(n5975), .ci(n5974), .co(n6027), .s(n5980) );
  fulladder U6632 ( .a(n5979), .b(n5978), .ci(n5977), .co(n6033), .s(n5981) );
  fulladder U6633 ( .a(n5982), .b(n5981), .ci(n5980), .co(n6031), .s(n5985) );
  fulladder U6634 ( .a(n5985), .b(n5984), .ci(n5983), .co(n6030), .s(
        \STAGE_1/M5/sum [0]) );
  nand2_1 U6635 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[71]), .op(n5987)
         );
  inv_1 U6636 ( .ip(m1Inputs[74]), .op(n12959) );
  nor3_1 U6637 ( .ip1(n13082), .ip2(n12959), .ip3(n5986), .op(n12546) );
  or2_1 U6638 ( .ip1(n5987), .ip2(n12546), .op(n5989) );
  nand2_1 U6639 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[74]), .op(n12958) );
  or2_1 U6640 ( .ip1(n12958), .ip2(n12546), .op(n5988) );
  nand2_1 U6641 ( .ip1(n5989), .ip2(n5988), .op(n12545) );
  inv_1 U6642 ( .ip(\STAGE_1/weightReg [10]), .op(n13594) );
  buf_1 U6643 ( .ip(n13594), .op(n13390) );
  nor2_1 U6644 ( .ip1(n12964), .ip2(n13390), .op(n12547) );
  xnor2_1 U6645 ( .ip1(n12545), .ip2(n12547), .op(n12585) );
  fulladder U6646 ( .a(n5992), .b(n5991), .ci(n5990), .co(n12584), .s(n5973)
         );
  fulladder U6647 ( .a(n5994), .b(n6011), .ci(n5993), .co(n12583), .s(n5958)
         );
  inv_1 U6648 ( .ip(n5995), .op(n12592) );
  or2_1 U6649 ( .ip1(n5996), .ip2(n5997), .op(n6000) );
  or2_1 U6650 ( .ip1(n5998), .ip2(n5997), .op(n5999) );
  nand2_1 U6651 ( .ip1(n6000), .ip2(n5999), .op(n12555) );
  or2_1 U6652 ( .ip1(n6001), .ip2(n6003), .op(n6006) );
  inv_1 U6653 ( .ip(n6002), .op(n6004) );
  or2_1 U6654 ( .ip1(n6004), .ip2(n6003), .op(n6005) );
  nand2_1 U6655 ( .ip1(n6006), .ip2(n6005), .op(n12554) );
  nand2_1 U6656 ( .ip1(n4672), .ip2(m1Inputs[72]), .op(n6008) );
  nor3_1 U6657 ( .ip1(n13854), .ip2(n13081), .ip3(n6007), .op(n12541) );
  or2_1 U6658 ( .ip1(n6008), .ip2(n12541), .op(n6010) );
  nand2_1 U6659 ( .ip1(n13707), .ip2(m1Inputs[73]), .op(n12565) );
  or2_1 U6660 ( .ip1(n12565), .ip2(n12541), .op(n6009) );
  nand2_1 U6661 ( .ip1(n6010), .ip2(n6009), .op(n12539) );
  nand2_1 U6662 ( .ip1(column[66]), .ip2(n13039), .op(n12540) );
  xor2_1 U6663 ( .ip1(n12539), .ip2(n12540), .op(n12553) );
  nor3_1 U6664 ( .ip1(n12925), .ip2(n14384), .ip3(n6011), .op(n12559) );
  nor2_1 U6665 ( .ip1(n12925), .ip2(n14289), .op(n12569) );
  or2_1 U6666 ( .ip1(n14835), .ip2(n12569), .op(n6013) );
  or2_1 U6667 ( .ip1(m1Inputs[67]), .ip2(n12569), .op(n6012) );
  nand2_1 U6668 ( .ip1(n6013), .ip2(n6012), .op(n12557) );
  nor2_1 U6669 ( .ip1(n12559), .ip2(n12557), .op(n6014) );
  nand2_1 U6670 ( .ip1(m1Inputs[66]), .ip2(n14975), .op(n12556) );
  xor2_1 U6671 ( .ip1(n6014), .ip2(n12556), .op(n12552) );
  nor2_1 U6672 ( .ip1(n6016), .ip2(n6015), .op(n6017) );
  nor2_1 U6673 ( .ip1(n6018), .ip2(n6017), .op(n12551) );
  nand2_1 U6674 ( .ip1(n14369), .ip2(m1Inputs[69]), .op(n6020) );
  nor3_1 U6675 ( .ip1(n13045), .ip2(n13835), .ip3(n6019), .op(n12561) );
  or2_1 U6676 ( .ip1(n6020), .ip2(n12561), .op(n6022) );
  nand2_1 U6677 ( .ip1(m1Inputs[70]), .ip2(n13637), .op(n12573) );
  or2_1 U6678 ( .ip1(n12573), .ip2(n12561), .op(n6021) );
  nand2_1 U6679 ( .ip1(n6022), .ip2(n6021), .op(n12560) );
  nor2_1 U6680 ( .ip1(n13076), .ip2(n12083), .op(n12562) );
  xnor2_1 U6681 ( .ip1(n12560), .ip2(n12562), .op(n12550) );
  fulladder U6682 ( .a(n6025), .b(n6024), .ci(n6023), .co(n12586), .s(n5952)
         );
  inv_1 U6683 ( .ip(n6026), .op(n12591) );
  fulladder U6684 ( .a(n6029), .b(n6028), .ci(n6027), .co(n12590), .s(n6034)
         );
  fulladder U6685 ( .a(n6032), .b(n6031), .ci(n6030), .co(n12594), .s(
        \STAGE_1/M5/sum [1]) );
  fulladder U6686 ( .a(n6035), .b(n6034), .ci(n6033), .co(n12593), .s(n6032)
         );
  nand2_1 U6687 ( .ip1(m1Inputs[4]), .ip2(n12699), .op(n6037) );
  nor3_1 U6688 ( .ip1(n10166), .ip2(n4624), .ip3(n6036), .op(n6109) );
  or2_1 U6689 ( .ip1(n6037), .ip2(n6109), .op(n6039) );
  nand2_1 U6690 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[5]), .op(n6104)
         );
  or2_1 U6691 ( .ip1(n6104), .ip2(n6109), .op(n6038) );
  nand2_1 U6692 ( .ip1(n6039), .ip2(n6038), .op(n6108) );
  nor2_1 U6693 ( .ip1(n10160), .ip2(n6503), .op(n6110) );
  xnor2_1 U6694 ( .ip1(n6108), .ip2(n6110), .op(n6164) );
  and3_1 U6695 ( .ip1(n9733), .ip2(m1Inputs[9]), .ip3(n6040), .op(n6103) );
  inv_1 U6696 ( .ip(m1Inputs[9]), .op(n10155) );
  nor2_1 U6697 ( .ip1(n13646), .ip2(n10155), .op(n6041) );
  or2_1 U6698 ( .ip1(m1Inputs[6]), .ip2(n6041), .op(n6043) );
  or2_1 U6699 ( .ip1(n9733), .ip2(n6041), .op(n6042) );
  nand2_1 U6700 ( .ip1(n6043), .ip2(n6042), .op(n6101) );
  nor2_1 U6701 ( .ip1(n6103), .ip2(n6101), .op(n6044) );
  nand2_1 U6702 ( .ip1(m1Inputs[0]), .ip2(n14994), .op(n6100) );
  xor2_1 U6703 ( .ip1(n6044), .ip2(n6100), .op(n6163) );
  fulladder U6704 ( .a(n6047), .b(n6046), .ci(n6045), .co(n6162), .s(n5670) );
  inv_1 U6705 ( .ip(n6048), .op(n6185) );
  inv_1 U6706 ( .ip(n6049), .op(n6053) );
  nor2_1 U6707 ( .ip1(n6051), .ip2(n6050), .op(n6052) );
  nor2_1 U6708 ( .ip1(n6053), .ip2(n6052), .op(n6155) );
  nand2_1 U6709 ( .ip1(m1Inputs[3]), .ip2(n12981), .op(n6154) );
  nand2_1 U6710 ( .ip1(m1Inputs[2]), .ip2(\STAGE_1/weightReg [7]), .op(n6153)
         );
  inv_1 U6711 ( .ip(n6054), .op(n6176) );
  or2_1 U6712 ( .ip1(n6055), .ip2(n6056), .op(n6059) );
  or2_1 U6713 ( .ip1(n6057), .ip2(n6056), .op(n6058) );
  nand2_1 U6714 ( .ip1(n6059), .ip2(n6058), .op(n6152) );
  or2_1 U6715 ( .ip1(n6060), .ip2(n6061), .op(n6064) );
  or2_1 U6716 ( .ip1(n6062), .ip2(n6061), .op(n6063) );
  nand2_1 U6717 ( .ip1(n6064), .ip2(n6063), .op(n6151) );
  nand2_1 U6718 ( .ip1(n4672), .ip2(m1Inputs[7]), .op(n6066) );
  nor3_1 U6719 ( .ip1(n10555), .ip2(n10072), .ip3(n6065), .op(n6115) );
  or2_1 U6720 ( .ip1(n6066), .ip2(n6115), .op(n6068) );
  nand2_1 U6721 ( .ip1(n12809), .ip2(m1Inputs[8]), .op(n6082) );
  or2_1 U6722 ( .ip1(n6082), .ip2(n6115), .op(n6067) );
  nand2_1 U6723 ( .ip1(n6068), .ip2(n6067), .op(n6113) );
  nand2_1 U6724 ( .ip1(column[1]), .ip2(n13859), .op(n6114) );
  xor2_1 U6725 ( .ip1(n6113), .ip2(n6114), .op(n6150) );
  inv_1 U6726 ( .ip(n6069), .op(n6175) );
  fulladder U6727 ( .a(n6072), .b(n6071), .ci(n6070), .co(n6174), .s(n6076) );
  fulladder U6728 ( .a(n6075), .b(n6074), .ci(n6073), .co(n6183), .s(n6077) );
  fulladder U6729 ( .a(n6078), .b(n6077), .ci(n6076), .co(n6181), .s(n6081) );
  fulladder U6730 ( .a(n6081), .b(n6080), .ci(n6079), .co(n6180), .s(
        \STAGE_1/M1/sum [0]) );
  nand2_1 U6731 ( .ip1(n4672), .ip2(m1Inputs[8]), .op(n6083) );
  nor3_1 U6732 ( .ip1(n10555), .ip2(n10155), .ip3(n6082), .op(n6086) );
  or2_1 U6733 ( .ip1(n6083), .ip2(n6086), .op(n6085) );
  nand2_1 U6734 ( .ip1(n10507), .ip2(m1Inputs[9]), .op(n6131) );
  or2_1 U6735 ( .ip1(n6131), .ip2(n6086), .op(n6084) );
  nand2_1 U6736 ( .ip1(n6085), .ip2(n6084), .op(n6120) );
  or2_1 U6737 ( .ip1(n6120), .ip2(n6086), .op(n6089) );
  nand2_1 U6738 ( .ip1(column[2]), .ip2(n13039), .op(n6119) );
  inv_1 U6739 ( .ip(n6119), .op(n6087) );
  or2_1 U6740 ( .ip1(n6087), .ip2(n6086), .op(n6088) );
  nand2_1 U6741 ( .ip1(n6089), .ip2(n6088), .op(n9726) );
  nand2_1 U6742 ( .ip1(n9733), .ip2(m1Inputs[7]), .op(n6091) );
  inv_1 U6743 ( .ip(m1Inputs[10]), .op(n10122) );
  nor3_1 U6744 ( .ip1(n13801), .ip2(n10122), .ip3(n6090), .op(n6094) );
  or2_1 U6745 ( .ip1(n6091), .ip2(n6094), .op(n6093) );
  nand2_1 U6746 ( .ip1(n13803), .ip2(m1Inputs[10]), .op(n10121) );
  or2_1 U6747 ( .ip1(n10121), .ip2(n6094), .op(n6092) );
  nand2_1 U6748 ( .ip1(n6093), .ip2(n6092), .op(n6149) );
  or2_1 U6749 ( .ip1(n6149), .ip2(n6094), .op(n6096) );
  nor2_1 U6750 ( .ip1(n10127), .ip2(n13594), .op(n6148) );
  or2_1 U6751 ( .ip1(n6148), .ip2(n6094), .op(n6095) );
  nand2_1 U6752 ( .ip1(n6096), .ip2(n6095), .op(n9725) );
  nand2_1 U6753 ( .ip1(m1Inputs[3]), .ip2(n14975), .op(n9724) );
  inv_1 U6754 ( .ip(n14836), .op(n13749) );
  nand2_1 U6755 ( .ip1(m1Inputs[4]), .ip2(n13749), .op(n6135) );
  nor3_1 U6756 ( .ip1(n10088), .ip2(n14368), .ip3(n6154), .op(n6122) );
  or2_1 U6757 ( .ip1(n6135), .ip2(n6122), .op(n6099) );
  nand2_1 U6758 ( .ip1(m1Inputs[3]), .ip2(n14835), .op(n6097) );
  or2_1 U6759 ( .ip1(n6097), .ip2(n6122), .op(n6098) );
  nand2_1 U6760 ( .ip1(n6099), .ip2(n6098), .op(n6121) );
  nor2_1 U6761 ( .ip1(n10150), .ip2(n6504), .op(n6123) );
  xnor2_1 U6762 ( .ip1(n6121), .ip2(n6123), .op(n6161) );
  nor2_1 U6763 ( .ip1(n6101), .ip2(n6100), .op(n6102) );
  nor2_1 U6764 ( .ip1(n6103), .ip2(n6102), .op(n6160) );
  nand2_1 U6765 ( .ip1(m1Inputs[5]), .ip2(\STAGE_1/weightReg [5]), .op(n6105)
         );
  nor3_1 U6766 ( .ip1(n9908), .ip2(n4624), .ip3(n6104), .op(n6127) );
  or2_1 U6767 ( .ip1(n6105), .ip2(n6127), .op(n6107) );
  nand2_1 U6768 ( .ip1(m1Inputs[6]), .ip2(\STAGE_1/weightReg [4]), .op(n6139)
         );
  or2_1 U6769 ( .ip1(n6139), .ip2(n6127), .op(n6106) );
  nand2_1 U6770 ( .ip1(n6107), .ip2(n6106), .op(n6126) );
  nor2_1 U6771 ( .ip1(n10160), .ip2(n12083), .op(n6128) );
  xnor2_1 U6772 ( .ip1(n6126), .ip2(n6128), .op(n6159) );
  or2_1 U6773 ( .ip1(n6108), .ip2(n6109), .op(n6112) );
  or2_1 U6774 ( .ip1(n6110), .ip2(n6109), .op(n6111) );
  nand2_1 U6775 ( .ip1(n6112), .ip2(n6111), .op(n6158) );
  or2_1 U6776 ( .ip1(n6113), .ip2(n6115), .op(n6118) );
  inv_1 U6777 ( .ip(n6114), .op(n6116) );
  or2_1 U6778 ( .ip1(n6116), .ip2(n6115), .op(n6117) );
  nand2_1 U6779 ( .ip1(n6118), .ip2(n6117), .op(n6157) );
  xor2_1 U6780 ( .ip1(n6120), .ip2(n6119), .op(n6156) );
  or2_1 U6781 ( .ip1(n6121), .ip2(n6122), .op(n6125) );
  or2_1 U6782 ( .ip1(n6123), .ip2(n6122), .op(n6124) );
  nand2_1 U6783 ( .ip1(n6125), .ip2(n6124), .op(n9710) );
  or2_1 U6784 ( .ip1(n6126), .ip2(n6127), .op(n6130) );
  or2_1 U6785 ( .ip1(n6128), .ip2(n6127), .op(n6129) );
  nand2_1 U6786 ( .ip1(n6130), .ip2(n6129), .op(n9709) );
  nand2_1 U6787 ( .ip1(n4619), .ip2(m1Inputs[9]), .op(n6132) );
  nor3_1 U6788 ( .ip1(n10555), .ip2(n10122), .ip3(n6131), .op(n9729) );
  or2_1 U6789 ( .ip1(n6132), .ip2(n9729), .op(n6134) );
  nand2_1 U6790 ( .ip1(n10507), .ip2(m1Inputs[10]), .op(n9700) );
  or2_1 U6791 ( .ip1(n9700), .ip2(n9729), .op(n6133) );
  nand2_1 U6792 ( .ip1(n6134), .ip2(n6133), .op(n9727) );
  nand2_1 U6793 ( .ip1(column[3]), .ip2(n13859), .op(n9728) );
  xor2_1 U6794 ( .ip1(n9727), .ip2(n9728), .op(n9708) );
  nand2_1 U6795 ( .ip1(m1Inputs[4]), .ip2(n14835), .op(n6136) );
  nor3_1 U6796 ( .ip1(n10166), .ip2(n14384), .ip3(n6135), .op(n9696) );
  or2_1 U6797 ( .ip1(n6136), .ip2(n9696), .op(n6138) );
  nand2_1 U6798 ( .ip1(m1Inputs[5]), .ip2(n12981), .op(n9720) );
  or2_1 U6799 ( .ip1(n9720), .ip2(n9696), .op(n6137) );
  nand2_1 U6800 ( .ip1(n6138), .ip2(n6137), .op(n9695) );
  nor2_1 U6801 ( .ip1(n10150), .ip2(n13766), .op(n9697) );
  xor2_1 U6802 ( .ip1(n9695), .ip2(n9697), .op(n9706) );
  nand2_1 U6803 ( .ip1(m1Inputs[6]), .ip2(\STAGE_1/weightReg [5]), .op(n6140)
         );
  inv_1 U6804 ( .ip(m1Inputs[7]), .op(n10145) );
  nor3_1 U6805 ( .ip1(n10145), .ip2(n4624), .ip3(n6139), .op(n9712) );
  or2_1 U6806 ( .ip1(n6140), .ip2(n9712), .op(n6142) );
  nand2_1 U6807 ( .ip1(m1Inputs[7]), .ip2(n11974), .op(n9716) );
  or2_1 U6808 ( .ip1(n9716), .ip2(n9712), .op(n6141) );
  nand2_1 U6809 ( .ip1(n6142), .ip2(n6141), .op(n9711) );
  nor2_1 U6810 ( .ip1(n10160), .ip2(n13594), .op(n9713) );
  xor2_1 U6811 ( .ip1(n9711), .ip2(n9713), .op(n9705) );
  nand2_1 U6812 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[8]), .op(n6144)
         );
  inv_1 U6813 ( .ip(m1Inputs[11]), .op(n10083) );
  nor3_1 U6814 ( .ip1(n13801), .ip2(n10083), .ip3(n6143), .op(n9691) );
  or2_1 U6815 ( .ip1(n6144), .ip2(n9691), .op(n6146) );
  nand2_1 U6816 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[11]), .op(n10082) );
  or2_1 U6817 ( .ip1(n10082), .ip2(n9691), .op(n6145) );
  nand2_1 U6818 ( .ip1(n6146), .ip2(n6145), .op(n9690) );
  inv_1 U6819 ( .ip(\STAGE_1/weightReg [11]), .op(n13579) );
  nor2_1 U6820 ( .ip1(n10127), .ip2(n13579), .op(n9692) );
  xor2_1 U6821 ( .ip1(n9690), .ip2(n9692), .op(n9704) );
  inv_1 U6822 ( .ip(n6147), .op(n9742) );
  xnor2_1 U6823 ( .ip1(n6149), .ip2(n6148), .op(n6168) );
  fulladder U6824 ( .a(n6152), .b(n6151), .ci(n6150), .co(n6167), .s(n6069) );
  fulladder U6825 ( .a(n6155), .b(n6154), .ci(n6153), .co(n6166), .s(n6054) );
  fulladder U6826 ( .a(n6158), .b(n6157), .ci(n6156), .co(n9738), .s(n6172) );
  fulladder U6827 ( .a(n6161), .b(n6160), .ci(n6159), .co(n9739), .s(n6171) );
  fulladder U6828 ( .a(n6164), .b(n6163), .ci(n6162), .co(n6170), .s(n6048) );
  inv_1 U6829 ( .ip(n6165), .op(n9751) );
  fulladder U6830 ( .a(n6168), .b(n6167), .ci(n6166), .co(n9741), .s(n6169) );
  inv_1 U6831 ( .ip(n6169), .op(n6179) );
  fulladder U6832 ( .a(n6172), .b(n6171), .ci(n6170), .co(n9745), .s(n6173) );
  inv_1 U6833 ( .ip(n6173), .op(n6178) );
  fulladder U6834 ( .a(n6176), .b(n6175), .ci(n6174), .co(n6177), .s(n6184) );
  fulladder U6835 ( .a(n6179), .b(n6178), .ci(n6177), .co(n9750), .s(n6188) );
  fulladder U6836 ( .a(n6182), .b(n6181), .ci(n6180), .co(n6187), .s(
        \STAGE_1/M1/sum [1]) );
  fulladder U6837 ( .a(n6185), .b(n6184), .ci(n6183), .co(n6186), .s(n6182) );
  fulladder U6838 ( .a(n6188), .b(n6187), .ci(n6186), .co(n9749), .s(
        \STAGE_1/M1/sum [2]) );
  nand2_1 U6839 ( .ip1(m1Inputs[36]), .ip2(n12699), .op(n6190) );
  nor3_1 U6840 ( .ip1(n8942), .ip2(n11555), .ip3(n6189), .op(n6262) );
  or2_1 U6841 ( .ip1(n6190), .ip2(n6262), .op(n6192) );
  nand2_1 U6842 ( .ip1(n13637), .ip2(m1Inputs[37]), .op(n6257) );
  or2_1 U6843 ( .ip1(n6257), .ip2(n6262), .op(n6191) );
  nand2_1 U6844 ( .ip1(n6192), .ip2(n6191), .op(n6261) );
  nor2_1 U6845 ( .ip1(n11549), .ip2(n6503), .op(n6263) );
  xnor2_1 U6846 ( .ip1(n6261), .ip2(n6263), .op(n6316) );
  and3_1 U6847 ( .ip1(n9733), .ip2(m1Inputs[41]), .ip3(n6193), .op(n6256) );
  inv_1 U6848 ( .ip(m1Inputs[41]), .op(n11544) );
  nor2_1 U6849 ( .ip1(n13646), .ip2(n11544), .op(n6194) );
  or2_1 U6850 ( .ip1(m1Inputs[38]), .ip2(n6194), .op(n6196) );
  or2_1 U6851 ( .ip1(n9733), .ip2(n6194), .op(n6195) );
  nand2_1 U6852 ( .ip1(n6196), .ip2(n6195), .op(n6254) );
  nor2_1 U6853 ( .ip1(n6256), .ip2(n6254), .op(n6197) );
  nand2_1 U6854 ( .ip1(m1Inputs[32]), .ip2(n14994), .op(n6253) );
  xor2_1 U6855 ( .ip1(n6197), .ip2(n6253), .op(n6315) );
  fulladder U6856 ( .a(n6200), .b(n6199), .ci(n6198), .co(n6314), .s(n5543) );
  inv_1 U6857 ( .ip(n6201), .op(n6337) );
  inv_1 U6858 ( .ip(n6202), .op(n6206) );
  nor2_1 U6859 ( .ip1(n6204), .ip2(n6203), .op(n6205) );
  nor2_1 U6860 ( .ip1(n6206), .ip2(n6205), .op(n6307) );
  nand2_1 U6861 ( .ip1(m1Inputs[35]), .ip2(n12981), .op(n6306) );
  nand2_1 U6862 ( .ip1(m1Inputs[34]), .ip2(n14835), .op(n6305) );
  inv_1 U6863 ( .ip(n6207), .op(n6328) );
  or2_1 U6864 ( .ip1(n6208), .ip2(n6209), .op(n6212) );
  or2_1 U6865 ( .ip1(n6210), .ip2(n6209), .op(n6211) );
  nand2_1 U6866 ( .ip1(n6212), .ip2(n6211), .op(n6304) );
  or2_1 U6867 ( .ip1(n6213), .ip2(n6214), .op(n6217) );
  or2_1 U6868 ( .ip1(n6215), .ip2(n6214), .op(n6216) );
  nand2_1 U6869 ( .ip1(n6217), .ip2(n6216), .op(n6303) );
  nand2_1 U6870 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[39]), .op(n6219)
         );
  nor3_1 U6871 ( .ip1(n13709), .ip2(n11461), .ip3(n6218), .op(n6268) );
  or2_1 U6872 ( .ip1(n6219), .ip2(n6268), .op(n6221) );
  nand2_1 U6873 ( .ip1(n12809), .ip2(m1Inputs[40]), .op(n6235) );
  or2_1 U6874 ( .ip1(n6235), .ip2(n6268), .op(n6220) );
  nand2_1 U6875 ( .ip1(n6221), .ip2(n6220), .op(n6266) );
  nand2_1 U6876 ( .ip1(column[33]), .ip2(n13039), .op(n6267) );
  xor2_1 U6877 ( .ip1(n6266), .ip2(n6267), .op(n6302) );
  inv_1 U6878 ( .ip(n6222), .op(n6327) );
  fulladder U6879 ( .a(n6225), .b(n6224), .ci(n6223), .co(n6326), .s(n6229) );
  fulladder U6880 ( .a(n6228), .b(n6227), .ci(n6226), .co(n6335), .s(n6230) );
  fulladder U6881 ( .a(n6231), .b(n6230), .ci(n6229), .co(n6333), .s(n6234) );
  fulladder U6882 ( .a(n6234), .b(n6233), .ci(n6232), .co(n6332), .s(
        \STAGE_1/M3/sum [0]) );
  nand2_1 U6883 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[40]), .op(n6236)
         );
  nor3_1 U6884 ( .ip1(n13709), .ip2(n11544), .ip3(n6235), .op(n6239) );
  or2_1 U6885 ( .ip1(n6236), .ip2(n6239), .op(n6238) );
  nand2_1 U6886 ( .ip1(n12809), .ip2(m1Inputs[41]), .op(n6283) );
  or2_1 U6887 ( .ip1(n6283), .ip2(n6239), .op(n6237) );
  nand2_1 U6888 ( .ip1(n6238), .ip2(n6237), .op(n6273) );
  or2_1 U6889 ( .ip1(n6273), .ip2(n6239), .op(n6242) );
  nand2_1 U6890 ( .ip1(column[34]), .ip2(n13039), .op(n6272) );
  inv_1 U6891 ( .ip(n6272), .op(n6240) );
  or2_1 U6892 ( .ip1(n6240), .ip2(n6239), .op(n6241) );
  nand2_1 U6893 ( .ip1(n6242), .ip2(n6241), .op(n11123) );
  nand2_1 U6894 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[39]), .op(n6244)
         );
  inv_1 U6895 ( .ip(m1Inputs[42]), .op(n11511) );
  nor3_1 U6896 ( .ip1(n13082), .ip2(n11511), .ip3(n6243), .op(n6247) );
  or2_1 U6897 ( .ip1(n6244), .ip2(n6247), .op(n6246) );
  nand2_1 U6898 ( .ip1(n13803), .ip2(m1Inputs[42]), .op(n11510) );
  or2_1 U6899 ( .ip1(n11510), .ip2(n6247), .op(n6245) );
  nand2_1 U6900 ( .ip1(n6246), .ip2(n6245), .op(n6301) );
  or2_1 U6901 ( .ip1(n6301), .ip2(n6247), .op(n6249) );
  nor2_1 U6902 ( .ip1(n11516), .ip2(n13390), .op(n6300) );
  or2_1 U6903 ( .ip1(n6300), .ip2(n6247), .op(n6248) );
  nand2_1 U6904 ( .ip1(n6249), .ip2(n6248), .op(n11122) );
  nand2_1 U6905 ( .ip1(m1Inputs[35]), .ip2(n14975), .op(n11121) );
  nor3_1 U6906 ( .ip1(n11477), .ip2(n14384), .ip3(n6306), .op(n6277) );
  nor2_1 U6907 ( .ip1(n11477), .ip2(n14289), .op(n6287) );
  or2_1 U6908 ( .ip1(n14835), .ip2(n6287), .op(n6251) );
  or2_1 U6909 ( .ip1(m1Inputs[35]), .ip2(n6287), .op(n6250) );
  nand2_1 U6910 ( .ip1(n6251), .ip2(n6250), .op(n6275) );
  nor2_1 U6911 ( .ip1(n6277), .ip2(n6275), .op(n6252) );
  nand2_1 U6912 ( .ip1(m1Inputs[34]), .ip2(n14975), .op(n6274) );
  xor2_1 U6913 ( .ip1(n6252), .ip2(n6274), .op(n6313) );
  nor2_1 U6914 ( .ip1(n6254), .ip2(n6253), .op(n6255) );
  nor2_1 U6915 ( .ip1(n6256), .ip2(n6255), .op(n6312) );
  nand2_1 U6916 ( .ip1(\STAGE_1/weightReg [5]), .ip2(m1Inputs[37]), .op(n6258)
         );
  nor3_1 U6917 ( .ip1(n11283), .ip2(n13835), .ip3(n6257), .op(n6279) );
  or2_1 U6918 ( .ip1(n6258), .ip2(n6279), .op(n6260) );
  nand2_1 U6919 ( .ip1(m1Inputs[38]), .ip2(n11974), .op(n6291) );
  or2_1 U6920 ( .ip1(n6291), .ip2(n6279), .op(n6259) );
  nand2_1 U6921 ( .ip1(n6260), .ip2(n6259), .op(n6278) );
  nor2_1 U6922 ( .ip1(n11549), .ip2(n13766), .op(n6280) );
  xnor2_1 U6923 ( .ip1(n6278), .ip2(n6280), .op(n6311) );
  or2_1 U6924 ( .ip1(n6261), .ip2(n6262), .op(n6265) );
  or2_1 U6925 ( .ip1(n6263), .ip2(n6262), .op(n6264) );
  nand2_1 U6926 ( .ip1(n6265), .ip2(n6264), .op(n6310) );
  or2_1 U6927 ( .ip1(n6266), .ip2(n6268), .op(n6271) );
  inv_1 U6928 ( .ip(n6267), .op(n6269) );
  or2_1 U6929 ( .ip1(n6269), .ip2(n6268), .op(n6270) );
  nand2_1 U6930 ( .ip1(n6271), .ip2(n6270), .op(n6309) );
  xor2_1 U6931 ( .ip1(n6273), .ip2(n6272), .op(n6308) );
  nor2_1 U6932 ( .ip1(n6275), .ip2(n6274), .op(n6276) );
  nor2_1 U6933 ( .ip1(n6277), .ip2(n6276), .op(n11107) );
  or2_1 U6934 ( .ip1(n6278), .ip2(n6279), .op(n6282) );
  or2_1 U6935 ( .ip1(n6280), .ip2(n6279), .op(n6281) );
  nand2_1 U6936 ( .ip1(n6282), .ip2(n6281), .op(n11106) );
  nand2_1 U6937 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[41]), .op(n6284)
         );
  nor3_1 U6938 ( .ip1(n13709), .ip2(n11511), .ip3(n6283), .op(n11126) );
  or2_1 U6939 ( .ip1(n6284), .ip2(n11126), .op(n6286) );
  nand2_1 U6940 ( .ip1(n12809), .ip2(m1Inputs[42]), .op(n11097) );
  or2_1 U6941 ( .ip1(n11097), .ip2(n11126), .op(n6285) );
  nand2_1 U6942 ( .ip1(n6286), .ip2(n6285), .op(n11124) );
  nand2_1 U6943 ( .ip1(column[35]), .ip2(n13039), .op(n11125) );
  xor2_1 U6944 ( .ip1(n11124), .ip2(n11125), .op(n11105) );
  nand2_1 U6945 ( .ip1(m1Inputs[36]), .ip2(n4627), .op(n6288) );
  and3_1 U6946 ( .ip1(n14835), .ip2(m1Inputs[37]), .ip3(n6287), .op(n11093) );
  or2_1 U6947 ( .ip1(n6288), .ip2(n11093), .op(n6290) );
  nand2_1 U6948 ( .ip1(n13749), .ip2(m1Inputs[37]), .op(n11117) );
  or2_1 U6949 ( .ip1(n11117), .ip2(n11093), .op(n6289) );
  nand2_1 U6950 ( .ip1(n6290), .ip2(n6289), .op(n11092) );
  nor2_1 U6951 ( .ip1(n11539), .ip2(n13766), .op(n11094) );
  xor2_1 U6952 ( .ip1(n11092), .ip2(n11094), .op(n11103) );
  nand2_1 U6953 ( .ip1(m1Inputs[38]), .ip2(n12699), .op(n6292) );
  inv_1 U6954 ( .ip(m1Inputs[39]), .op(n11534) );
  nor3_1 U6955 ( .ip1(n11534), .ip2(n13835), .ip3(n6291), .op(n11109) );
  or2_1 U6956 ( .ip1(n6292), .ip2(n11109), .op(n6294) );
  nand2_1 U6957 ( .ip1(m1Inputs[39]), .ip2(n11974), .op(n11113) );
  or2_1 U6958 ( .ip1(n11113), .ip2(n11109), .op(n6293) );
  nand2_1 U6959 ( .ip1(n6294), .ip2(n6293), .op(n11108) );
  nor2_1 U6960 ( .ip1(n11549), .ip2(n13594), .op(n11110) );
  xor2_1 U6961 ( .ip1(n11108), .ip2(n11110), .op(n11102) );
  nand2_1 U6962 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[40]), .op(n6296)
         );
  inv_1 U6963 ( .ip(m1Inputs[43]), .op(n11472) );
  nor3_1 U6964 ( .ip1(n13082), .ip2(n11472), .ip3(n6295), .op(n11088) );
  or2_1 U6965 ( .ip1(n6296), .ip2(n11088), .op(n6298) );
  nand2_1 U6966 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[43]), .op(n11471) );
  or2_1 U6967 ( .ip1(n11471), .ip2(n11088), .op(n6297) );
  nand2_1 U6968 ( .ip1(n6298), .ip2(n6297), .op(n11087) );
  nor2_1 U6969 ( .ip1(n11516), .ip2(n13579), .op(n11089) );
  xor2_1 U6970 ( .ip1(n11087), .ip2(n11089), .op(n11101) );
  inv_1 U6971 ( .ip(n6299), .op(n11138) );
  xnor2_1 U6972 ( .ip1(n6301), .ip2(n6300), .op(n6320) );
  fulladder U6973 ( .a(n6304), .b(n6303), .ci(n6302), .co(n6319), .s(n6222) );
  fulladder U6974 ( .a(n6307), .b(n6306), .ci(n6305), .co(n6318), .s(n6207) );
  fulladder U6975 ( .a(n6310), .b(n6309), .ci(n6308), .co(n11134), .s(n6324)
         );
  fulladder U6976 ( .a(n6313), .b(n6312), .ci(n6311), .co(n11135), .s(n6323)
         );
  fulladder U6977 ( .a(n6316), .b(n6315), .ci(n6314), .co(n6322), .s(n6201) );
  inv_1 U6978 ( .ip(n6317), .op(n11147) );
  fulladder U6979 ( .a(n6320), .b(n6319), .ci(n6318), .co(n11137), .s(n6321)
         );
  inv_1 U6980 ( .ip(n6321), .op(n6331) );
  fulladder U6981 ( .a(n6324), .b(n6323), .ci(n6322), .co(n11141), .s(n6325)
         );
  inv_1 U6982 ( .ip(n6325), .op(n6330) );
  fulladder U6983 ( .a(n6328), .b(n6327), .ci(n6326), .co(n6329), .s(n6336) );
  fulladder U6984 ( .a(n6331), .b(n6330), .ci(n6329), .co(n11146), .s(n6340)
         );
  fulladder U6985 ( .a(n6334), .b(n6333), .ci(n6332), .co(n6339), .s(
        \STAGE_1/M3/sum [1]) );
  fulladder U6986 ( .a(n6337), .b(n6336), .ci(n6335), .co(n6338), .s(n6334) );
  fulladder U6987 ( .a(n6340), .b(n6339), .ci(n6338), .co(n11145), .s(
        \STAGE_1/M3/sum [2]) );
  nand2_1 U6988 ( .ip1(m1Inputs[84]), .ip2(\STAGE_1/weightReg [5]), .op(n6342)
         );
  nor3_1 U6989 ( .ip1(n8942), .ip2(n13847), .ip3(n6341), .op(n6414) );
  or2_1 U6990 ( .ip1(n6342), .ip2(n6414), .op(n6344) );
  nand2_1 U6991 ( .ip1(n13637), .ip2(m1Inputs[85]), .op(n6409) );
  or2_1 U6992 ( .ip1(n6409), .ip2(n6414), .op(n6343) );
  nand2_1 U6993 ( .ip1(n6344), .ip2(n6343), .op(n6413) );
  nor2_1 U6994 ( .ip1(n13841), .ip2(n6504), .op(n6415) );
  xnor2_1 U6995 ( .ip1(n6413), .ip2(n6415), .op(n6468) );
  and3_1 U6996 ( .ip1(n12578), .ip2(m1Inputs[89]), .ip3(n6345), .op(n6408) );
  inv_1 U6997 ( .ip(m1Inputs[89]), .op(n13836) );
  nor2_1 U6998 ( .ip1(n10476), .ip2(n13836), .op(n6346) );
  or2_1 U6999 ( .ip1(m1Inputs[86]), .ip2(n6346), .op(n6348) );
  or2_1 U7000 ( .ip1(n9733), .ip2(n6346), .op(n6347) );
  nand2_1 U7001 ( .ip1(n6348), .ip2(n6347), .op(n6406) );
  nor2_1 U7002 ( .ip1(n6408), .ip2(n6406), .op(n6349) );
  nand2_1 U7003 ( .ip1(m1Inputs[80]), .ip2(n14994), .op(n6405) );
  xor2_1 U7004 ( .ip1(n6349), .ip2(n6405), .op(n6467) );
  fulladder U7005 ( .a(n6352), .b(n6351), .ci(n6350), .co(n6466), .s(n5416) );
  inv_1 U7006 ( .ip(n6353), .op(n6489) );
  inv_1 U7007 ( .ip(n6354), .op(n6358) );
  nor2_1 U7008 ( .ip1(n6356), .ip2(n6355), .op(n6357) );
  nor2_1 U7009 ( .ip1(n6358), .ip2(n6357), .op(n6459) );
  nand2_1 U7010 ( .ip1(m1Inputs[83]), .ip2(n12981), .op(n6458) );
  nand2_1 U7011 ( .ip1(m1Inputs[82]), .ip2(\STAGE_1/weightReg [7]), .op(n6457)
         );
  inv_1 U7012 ( .ip(n6359), .op(n6480) );
  or2_1 U7013 ( .ip1(n6360), .ip2(n6361), .op(n6364) );
  or2_1 U7014 ( .ip1(n6362), .ip2(n6361), .op(n6363) );
  nand2_1 U7015 ( .ip1(n6364), .ip2(n6363), .op(n6456) );
  or2_1 U7016 ( .ip1(n6365), .ip2(n6366), .op(n6369) );
  or2_1 U7017 ( .ip1(n6367), .ip2(n6366), .op(n6368) );
  nand2_1 U7018 ( .ip1(n6369), .ip2(n6368), .op(n6455) );
  nand2_1 U7019 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[87]), .op(n6371)
         );
  nor3_1 U7020 ( .ip1(n13709), .ip2(n13748), .ip3(n6370), .op(n6420) );
  or2_1 U7021 ( .ip1(n6371), .ip2(n6420), .op(n6373) );
  nand2_1 U7022 ( .ip1(n13707), .ip2(m1Inputs[88]), .op(n6387) );
  or2_1 U7023 ( .ip1(n6387), .ip2(n6420), .op(n6372) );
  nand2_1 U7024 ( .ip1(n6373), .ip2(n6372), .op(n6418) );
  nand2_1 U7025 ( .ip1(column[81]), .ip2(n13859), .op(n6419) );
  xor2_1 U7026 ( .ip1(n6418), .ip2(n6419), .op(n6454) );
  inv_1 U7027 ( .ip(n6374), .op(n6479) );
  fulladder U7028 ( .a(n6377), .b(n6376), .ci(n6375), .co(n6478), .s(n6381) );
  fulladder U7029 ( .a(n6380), .b(n6379), .ci(n6378), .co(n6487), .s(n6382) );
  fulladder U7030 ( .a(n6383), .b(n6382), .ci(n6381), .co(n6485), .s(n6386) );
  fulladder U7031 ( .a(n6386), .b(n6385), .ci(n6384), .co(n6484), .s(
        \STAGE_1/M6/sum [0]) );
  nand2_1 U7032 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[88]), .op(n6388)
         );
  nor3_1 U7033 ( .ip1(n13709), .ip2(n13836), .ip3(n6387), .op(n6391) );
  or2_1 U7034 ( .ip1(n6388), .ip2(n6391), .op(n6390) );
  nand2_1 U7035 ( .ip1(n13707), .ip2(m1Inputs[89]), .op(n6435) );
  or2_1 U7036 ( .ip1(n6435), .ip2(n6391), .op(n6389) );
  nand2_1 U7037 ( .ip1(n6390), .ip2(n6389), .op(n6425) );
  or2_1 U7038 ( .ip1(n6425), .ip2(n6391), .op(n6394) );
  nand2_1 U7039 ( .ip1(column[82]), .ip2(n13859), .op(n6424) );
  inv_1 U7040 ( .ip(n6424), .op(n6392) );
  or2_1 U7041 ( .ip1(n6392), .ip2(n6391), .op(n6393) );
  nand2_1 U7042 ( .ip1(n6394), .ip2(n6393), .op(n13393) );
  nand2_1 U7043 ( .ip1(n13614), .ip2(m1Inputs[87]), .op(n6396) );
  inv_1 U7044 ( .ip(m1Inputs[90]), .op(n13800) );
  nor3_1 U7045 ( .ip1(n13082), .ip2(n13800), .ip3(n6395), .op(n6399) );
  or2_1 U7046 ( .ip1(n6396), .ip2(n6399), .op(n6398) );
  nand2_1 U7047 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[90]), .op(n13799) );
  or2_1 U7048 ( .ip1(n13799), .ip2(n6399), .op(n6397) );
  nand2_1 U7049 ( .ip1(n6398), .ip2(n6397), .op(n6453) );
  or2_1 U7050 ( .ip1(n6453), .ip2(n6399), .op(n6401) );
  nor2_1 U7051 ( .ip1(n13807), .ip2(n13594), .op(n6452) );
  or2_1 U7052 ( .ip1(n6452), .ip2(n6399), .op(n6400) );
  nand2_1 U7053 ( .ip1(n6401), .ip2(n6400), .op(n13392) );
  nand2_1 U7054 ( .ip1(m1Inputs[83]), .ip2(n14975), .op(n13391) );
  nor3_1 U7055 ( .ip1(n13765), .ip2(n14384), .ip3(n6458), .op(n6429) );
  nor2_1 U7056 ( .ip1(n13765), .ip2(n14836), .op(n6439) );
  or2_1 U7057 ( .ip1(n14835), .ip2(n6439), .op(n6403) );
  or2_1 U7058 ( .ip1(m1Inputs[83]), .ip2(n6439), .op(n6402) );
  nand2_1 U7059 ( .ip1(n6403), .ip2(n6402), .op(n6427) );
  nor2_1 U7060 ( .ip1(n6429), .ip2(n6427), .op(n6404) );
  nand2_1 U7061 ( .ip1(m1Inputs[82]), .ip2(n14975), .op(n6426) );
  xor2_1 U7062 ( .ip1(n6404), .ip2(n6426), .op(n6465) );
  nor2_1 U7063 ( .ip1(n6406), .ip2(n6405), .op(n6407) );
  nor2_1 U7064 ( .ip1(n6408), .ip2(n6407), .op(n6464) );
  nand2_1 U7065 ( .ip1(n14369), .ip2(m1Inputs[85]), .op(n6410) );
  nor3_1 U7066 ( .ip1(n13578), .ip2(n13835), .ip3(n6409), .op(n6431) );
  or2_1 U7067 ( .ip1(n6410), .ip2(n6431), .op(n6412) );
  nand2_1 U7068 ( .ip1(m1Inputs[86]), .ip2(n13637), .op(n6443) );
  or2_1 U7069 ( .ip1(n6443), .ip2(n6431), .op(n6411) );
  nand2_1 U7070 ( .ip1(n6412), .ip2(n6411), .op(n6430) );
  nor2_1 U7071 ( .ip1(n13841), .ip2(n13766), .op(n6432) );
  xnor2_1 U7072 ( .ip1(n6430), .ip2(n6432), .op(n6463) );
  or2_1 U7073 ( .ip1(n6413), .ip2(n6414), .op(n6417) );
  or2_1 U7074 ( .ip1(n6415), .ip2(n6414), .op(n6416) );
  nand2_1 U7075 ( .ip1(n6417), .ip2(n6416), .op(n6462) );
  or2_1 U7076 ( .ip1(n6418), .ip2(n6420), .op(n6423) );
  inv_1 U7077 ( .ip(n6419), .op(n6421) );
  or2_1 U7078 ( .ip1(n6421), .ip2(n6420), .op(n6422) );
  nand2_1 U7079 ( .ip1(n6423), .ip2(n6422), .op(n6461) );
  xor2_1 U7080 ( .ip1(n6425), .ip2(n6424), .op(n6460) );
  nor2_1 U7081 ( .ip1(n6427), .ip2(n6426), .op(n6428) );
  nor2_1 U7082 ( .ip1(n6429), .ip2(n6428), .op(n13376) );
  or2_1 U7083 ( .ip1(n6430), .ip2(n6431), .op(n6434) );
  or2_1 U7084 ( .ip1(n6432), .ip2(n6431), .op(n6433) );
  nand2_1 U7085 ( .ip1(n6434), .ip2(n6433), .op(n13375) );
  nand2_1 U7086 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[89]), .op(n6436)
         );
  nor3_1 U7087 ( .ip1(n13709), .ip2(n13800), .ip3(n6435), .op(n13396) );
  or2_1 U7088 ( .ip1(n6436), .ip2(n13396), .op(n6438) );
  nand2_1 U7089 ( .ip1(n13707), .ip2(m1Inputs[90]), .op(n13366) );
  or2_1 U7090 ( .ip1(n13366), .ip2(n13396), .op(n6437) );
  nand2_1 U7091 ( .ip1(n6438), .ip2(n6437), .op(n13394) );
  nand2_1 U7092 ( .ip1(column[83]), .ip2(n13859), .op(n13395) );
  xor2_1 U7093 ( .ip1(n13394), .ip2(n13395), .op(n13374) );
  nand2_1 U7094 ( .ip1(m1Inputs[84]), .ip2(\STAGE_1/weightReg [7]), .op(n6440)
         );
  and3_1 U7095 ( .ip1(n4627), .ip2(m1Inputs[85]), .ip3(n6439), .op(n13362) );
  or2_1 U7096 ( .ip1(n6440), .ip2(n13362), .op(n6442) );
  nand2_1 U7097 ( .ip1(n13749), .ip2(m1Inputs[85]), .op(n13386) );
  or2_1 U7098 ( .ip1(n13386), .ip2(n13362), .op(n6441) );
  nand2_1 U7099 ( .ip1(n6442), .ip2(n6441), .op(n13361) );
  nor2_1 U7100 ( .ip1(n13830), .ip2(n12083), .op(n13363) );
  xor2_1 U7101 ( .ip1(n13361), .ip2(n13363), .op(n13372) );
  nand2_1 U7102 ( .ip1(m1Inputs[86]), .ip2(\STAGE_1/weightReg [5]), .op(n6444)
         );
  inv_1 U7103 ( .ip(m1Inputs[87]), .op(n13825) );
  nor3_1 U7104 ( .ip1(n13825), .ip2(n13835), .ip3(n6443), .op(n13378) );
  or2_1 U7105 ( .ip1(n6444), .ip2(n13378), .op(n6446) );
  nand2_1 U7106 ( .ip1(m1Inputs[87]), .ip2(n13637), .op(n13382) );
  or2_1 U7107 ( .ip1(n13382), .ip2(n13378), .op(n6445) );
  nand2_1 U7108 ( .ip1(n6446), .ip2(n6445), .op(n13377) );
  nor2_1 U7109 ( .ip1(n13841), .ip2(n13594), .op(n13379) );
  xor2_1 U7110 ( .ip1(n13377), .ip2(n13379), .op(n13371) );
  nand2_1 U7111 ( .ip1(n13614), .ip2(m1Inputs[88]), .op(n6448) );
  and3_1 U7112 ( .ip1(n12578), .ip2(m1Inputs[91]), .ip3(n6447), .op(n13357) );
  or2_1 U7113 ( .ip1(n6448), .ip2(n13357), .op(n6450) );
  nand2_1 U7114 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[91]), .op(n13759) );
  or2_1 U7115 ( .ip1(n13759), .ip2(n13357), .op(n6449) );
  nand2_1 U7116 ( .ip1(n6450), .ip2(n6449), .op(n13356) );
  buf_1 U7117 ( .ip(n13579), .op(n14824) );
  nor2_1 U7118 ( .ip1(n13807), .ip2(n14824), .op(n13358) );
  xor2_1 U7119 ( .ip1(n13356), .ip2(n13358), .op(n13370) );
  inv_1 U7120 ( .ip(n6451), .op(n13408) );
  xnor2_1 U7121 ( .ip1(n6453), .ip2(n6452), .op(n6472) );
  fulladder U7122 ( .a(n6456), .b(n6455), .ci(n6454), .co(n6471), .s(n6374) );
  fulladder U7123 ( .a(n6459), .b(n6458), .ci(n6457), .co(n6470), .s(n6359) );
  fulladder U7124 ( .a(n6462), .b(n6461), .ci(n6460), .co(n13404), .s(n6476)
         );
  fulladder U7125 ( .a(n6465), .b(n6464), .ci(n6463), .co(n13405), .s(n6475)
         );
  fulladder U7126 ( .a(n6468), .b(n6467), .ci(n6466), .co(n6474), .s(n6353) );
  inv_1 U7127 ( .ip(n6469), .op(n13417) );
  fulladder U7128 ( .a(n6472), .b(n6471), .ci(n6470), .co(n13407), .s(n6473)
         );
  inv_1 U7129 ( .ip(n6473), .op(n6483) );
  fulladder U7130 ( .a(n6476), .b(n6475), .ci(n6474), .co(n13411), .s(n6477)
         );
  inv_1 U7131 ( .ip(n6477), .op(n6482) );
  fulladder U7132 ( .a(n6480), .b(n6479), .ci(n6478), .co(n6481), .s(n6488) );
  fulladder U7133 ( .a(n6483), .b(n6482), .ci(n6481), .co(n13416), .s(n6492)
         );
  fulladder U7134 ( .a(n6486), .b(n6485), .ci(n6484), .co(n6491), .s(
        \STAGE_1/M6/sum [1]) );
  fulladder U7135 ( .a(n6489), .b(n6488), .ci(n6487), .co(n6490), .s(n6486) );
  fulladder U7136 ( .a(n6492), .b(n6491), .ci(n6490), .co(n13415), .s(
        \STAGE_1/M6/sum [2]) );
  nand2_1 U7137 ( .ip1(m1Inputs[23]), .ip2(n12699), .op(n6493) );
  nand2_1 U7138 ( .ip1(m1Inputs[23]), .ip2(n11974), .op(n6563) );
  nor3_1 U7139 ( .ip1(n10812), .ip2(n12746), .ip3(n6563), .op(n6496) );
  or2_1 U7140 ( .ip1(n6493), .ip2(n6496), .op(n6495) );
  nand2_1 U7141 ( .ip1(m1Inputs[24]), .ip2(n11974), .op(n6512) );
  or2_1 U7142 ( .ip1(n6512), .ip2(n6496), .op(n6494) );
  nand2_1 U7143 ( .ip1(n6495), .ip2(n6494), .op(n6570) );
  or2_1 U7144 ( .ip1(n6570), .ip2(n6496), .op(n6498) );
  nor2_1 U7145 ( .ip1(n10472), .ip2(n13579), .op(n6569) );
  or2_1 U7146 ( .ip1(n6569), .ip2(n6496), .op(n6497) );
  nand2_1 U7147 ( .ip1(n6498), .ip2(n6497), .op(n10652) );
  nand2_1 U7148 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[28]), .op(n10600) );
  nor3_1 U7149 ( .ip1(n10476), .ip2(n10753), .ip3(n10600), .op(n6593) );
  nor2_1 U7150 ( .ip1(n13801), .ip2(n10753), .op(n6499) );
  or2_1 U7151 ( .ip1(m1Inputs[28]), .ip2(n6499), .op(n6501) );
  or2_1 U7152 ( .ip1(n13803), .ip2(n6499), .op(n6500) );
  nand2_1 U7153 ( .ip1(n6501), .ip2(n6500), .op(n6592) );
  inv_1 U7154 ( .ip(\STAGE_1/weightReg [12]), .op(n14902) );
  inv_1 U7155 ( .ip(n14902), .op(n15025) );
  nand2_1 U7156 ( .ip1(m1Inputs[16]), .ip2(n15025), .op(n6594) );
  nor2_1 U7157 ( .ip1(n6592), .ip2(n6594), .op(n6502) );
  nor2_1 U7158 ( .ip1(n6593), .ip2(n6502), .op(n10651) );
  nand2_1 U7159 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[20]), .op(n6591)
         );
  nor3_1 U7160 ( .ip1(n13766), .ip2(n10866), .ip3(n6591), .op(n10578) );
  nor2_1 U7161 ( .ip1(n12083), .ip2(n10493), .op(n10525) );
  or2_1 U7162 ( .ip1(m1Inputs[21]), .ip2(n10525), .op(n6506) );
  buf_1 U7163 ( .ip(n6503), .op(n6504) );
  inv_1 U7164 ( .ip(n6504), .op(n14838) );
  or2_1 U7165 ( .ip1(n14838), .ip2(n10525), .op(n6505) );
  nand2_1 U7166 ( .ip1(n6506), .ip2(n6505), .op(n10576) );
  nor2_1 U7167 ( .ip1(n10578), .ip2(n10576), .op(n6507) );
  inv_1 U7168 ( .ip(n13594), .op(n14629) );
  buf_1 U7169 ( .ip(n14629), .op(n14876) );
  nand2_1 U7170 ( .ip1(m1Inputs[19]), .ip2(\STAGE_1/weightReg [10]), .op(
        n10575) );
  xor2_1 U7171 ( .ip1(n6507), .ip2(n10575), .op(n10650) );
  nand2_1 U7172 ( .ip1(n13803), .ip2(m1Inputs[26]), .op(n6582) );
  nand2_1 U7173 ( .ip1(n9733), .ip2(m1Inputs[29]), .op(n10501) );
  nor2_1 U7174 ( .ip1(n6582), .ip2(n10501), .op(n10521) );
  inv_1 U7175 ( .ip(m1Inputs[26]), .op(n10827) );
  nor2_1 U7176 ( .ip1(n13082), .ip2(n10827), .op(n6508) );
  or2_1 U7177 ( .ip1(m1Inputs[29]), .ip2(n6508), .op(n6510) );
  or2_1 U7178 ( .ip1(n13803), .ip2(n6508), .op(n6509) );
  nand2_1 U7179 ( .ip1(n6510), .ip2(n6509), .op(n6511) );
  nor2_1 U7180 ( .ip1(n10521), .ip2(n6511), .op(n10520) );
  inv_1 U7181 ( .ip(\STAGE_1/weightReg [13]), .op(n14340) );
  nor2_1 U7182 ( .ip1(n9995), .ip2(n14340), .op(n10522) );
  xor2_1 U7183 ( .ip1(n10520), .ip2(n10522), .op(n10680) );
  nand2_1 U7184 ( .ip1(m1Inputs[24]), .ip2(n12699), .op(n6513) );
  nor3_1 U7185 ( .ip1(n10753), .ip2(n4624), .ip3(n6512), .op(n10569) );
  or2_1 U7186 ( .ip1(n6513), .ip2(n10569), .op(n6515) );
  nand2_1 U7187 ( .ip1(m1Inputs[25]), .ip2(n11974), .op(n10530) );
  or2_1 U7188 ( .ip1(n10530), .ip2(n10569), .op(n6514) );
  nand2_1 U7189 ( .ip1(n6515), .ip2(n6514), .op(n10568) );
  buf_1 U7190 ( .ip(n14902), .op(n14188) );
  nor2_1 U7191 ( .ip1(n10472), .ip2(n14188), .op(n10570) );
  xor2_1 U7192 ( .ip1(n10568), .ip2(n10570), .op(n10679) );
  nand2_1 U7193 ( .ip1(m1Inputs[22]), .ip2(n14835), .op(n6516) );
  nand2_1 U7194 ( .ip1(m1Inputs[22]), .ip2(n13749), .op(n6528) );
  nor3_1 U7195 ( .ip1(n10734), .ip2(n14368), .ip3(n6528), .op(n10564) );
  or2_1 U7196 ( .ip1(n6516), .ip2(n10564), .op(n6518) );
  nand2_1 U7197 ( .ip1(m1Inputs[23]), .ip2(n12981), .op(n10777) );
  or2_1 U7198 ( .ip1(n10777), .ip2(n10564), .op(n6517) );
  nand2_1 U7199 ( .ip1(n6518), .ip2(n6517), .op(n10563) );
  nor2_1 U7200 ( .ip1(n10585), .ip2(n13579), .op(n10565) );
  xor2_1 U7201 ( .ip1(n10563), .ip2(n10565), .op(n10678) );
  inv_1 U7202 ( .ip(n6519), .op(n10693) );
  nand2_1 U7203 ( .ip1(n4672), .ip2(m1Inputs[26]), .op(n6520) );
  inv_1 U7204 ( .ip(m1Inputs[27]), .op(n10751) );
  nand2_1 U7205 ( .ip1(n10507), .ip2(m1Inputs[26]), .op(n6539) );
  nor3_1 U7206 ( .ip1(n10555), .ip2(n10751), .ip3(n6539), .op(n6523) );
  or2_1 U7207 ( .ip1(n6520), .ip2(n6523), .op(n6522) );
  nand2_1 U7208 ( .ip1(n13707), .ip2(m1Inputs[27]), .op(n6534) );
  or2_1 U7209 ( .ip1(n6534), .ip2(n6523), .op(n6521) );
  nand2_1 U7210 ( .ip1(n6522), .ip2(n6521), .op(n6561) );
  or2_1 U7211 ( .ip1(n6561), .ip2(n6523), .op(n6526) );
  nand2_1 U7212 ( .ip1(column[20]), .ip2(n13859), .op(n6560) );
  inv_1 U7213 ( .ip(n6560), .op(n6524) );
  or2_1 U7214 ( .ip1(n6524), .ip2(n6523), .op(n6525) );
  nand2_1 U7215 ( .ip1(n6526), .ip2(n6525), .op(n10635) );
  nand2_1 U7216 ( .ip1(\STAGE_1/weightReg [7]), .ip2(m1Inputs[21]), .op(n6527)
         );
  nand2_1 U7217 ( .ip1(n13749), .ip2(m1Inputs[21]), .op(n6554) );
  nor3_1 U7218 ( .ip1(n10867), .ip2(n14384), .ip3(n6554), .op(n6531) );
  or2_1 U7219 ( .ip1(n6527), .ip2(n6531), .op(n6530) );
  or2_1 U7220 ( .ip1(n6528), .ip2(n6531), .op(n6529) );
  nand2_1 U7221 ( .ip1(n6530), .ip2(n6529), .op(n6572) );
  or2_1 U7222 ( .ip1(n6572), .ip2(n6531), .op(n6533) );
  nor2_1 U7223 ( .ip1(n10585), .ip2(n13594), .op(n6571) );
  or2_1 U7224 ( .ip1(n6571), .ip2(n6531), .op(n6532) );
  nand2_1 U7225 ( .ip1(n6533), .ip2(n6532), .op(n10634) );
  nand2_1 U7226 ( .ip1(n4619), .ip2(m1Inputs[27]), .op(n6535) );
  inv_1 U7227 ( .ip(m1Inputs[28]), .op(n11033) );
  nor3_1 U7228 ( .ip1(n10555), .ip2(n11033), .ip3(n6534), .op(n10581) );
  or2_1 U7229 ( .ip1(n6535), .ip2(n10581), .op(n6537) );
  nand2_1 U7230 ( .ip1(n12809), .ip2(m1Inputs[28]), .op(n10505) );
  or2_1 U7231 ( .ip1(n10505), .ip2(n10581), .op(n6536) );
  nand2_1 U7232 ( .ip1(n6537), .ip2(n6536), .op(n10579) );
  nand2_1 U7233 ( .ip1(column[21]), .ip2(n13859), .op(n10580) );
  xor2_1 U7234 ( .ip1(n10579), .ip2(n10580), .op(n10633) );
  nand2_1 U7235 ( .ip1(n5056), .ip2(m1Inputs[25]), .op(n6538) );
  nand2_1 U7236 ( .ip1(n12809), .ip2(m1Inputs[25]), .op(n6575) );
  nor3_1 U7237 ( .ip1(n10555), .ip2(n10827), .ip3(n6575), .op(n6542) );
  or2_1 U7238 ( .ip1(n6538), .ip2(n6542), .op(n6541) );
  or2_1 U7239 ( .ip1(n6539), .ip2(n6542), .op(n6540) );
  nand2_1 U7240 ( .ip1(n6541), .ip2(n6540), .op(n6619) );
  or2_1 U7241 ( .ip1(n6619), .ip2(n6542), .op(n6545) );
  nand2_1 U7242 ( .ip1(column[19]), .ip2(n13859), .op(n6618) );
  inv_1 U7243 ( .ip(n6618), .op(n6543) );
  or2_1 U7244 ( .ip1(n6543), .ip2(n6542), .op(n6544) );
  nand2_1 U7245 ( .ip1(n6545), .ip2(n6544), .op(n6590) );
  nand2_1 U7246 ( .ip1(m1Inputs[19]), .ip2(n14994), .op(n6589) );
  nand2_1 U7247 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[24]), .op(n6547)
         );
  nor3_1 U7248 ( .ip1(n13082), .ip2(n10751), .ip3(n6546), .op(n6550) );
  or2_1 U7249 ( .ip1(n6547), .ip2(n6550), .op(n6549) );
  nand2_1 U7250 ( .ip1(n13803), .ip2(m1Inputs[27]), .op(n10545) );
  or2_1 U7251 ( .ip1(n10545), .ip2(n6550), .op(n6548) );
  nand2_1 U7252 ( .ip1(n6549), .ip2(n6548), .op(n6604) );
  or2_1 U7253 ( .ip1(n6604), .ip2(n6550), .op(n6552) );
  nor2_1 U7254 ( .ip1(n9995), .ip2(n13579), .op(n6603) );
  or2_1 U7255 ( .ip1(n6603), .ip2(n6550), .op(n6551) );
  nand2_1 U7256 ( .ip1(n6552), .ip2(n6551), .op(n6598) );
  nand2_1 U7257 ( .ip1(m1Inputs[20]), .ip2(n14835), .op(n6553) );
  nor2_1 U7258 ( .ip1(n10493), .ip2(n14289), .op(n6606) );
  and3_1 U7259 ( .ip1(n4627), .ip2(m1Inputs[21]), .ip3(n6606), .op(n6557) );
  or2_1 U7260 ( .ip1(n6553), .ip2(n6557), .op(n6556) );
  or2_1 U7261 ( .ip1(n6554), .ip2(n6557), .op(n6555) );
  nand2_1 U7262 ( .ip1(n6556), .ip2(n6555), .op(n6600) );
  or2_1 U7263 ( .ip1(n6600), .ip2(n6557), .op(n6559) );
  nor2_1 U7264 ( .ip1(n10585), .ip2(n13766), .op(n6599) );
  or2_1 U7265 ( .ip1(n6599), .ip2(n6557), .op(n6558) );
  nand2_1 U7266 ( .ip1(n6559), .ip2(n6558), .op(n6597) );
  xor2_1 U7267 ( .ip1(n6561), .ip2(n6560), .op(n6596) );
  nand2_1 U7268 ( .ip1(m1Inputs[22]), .ip2(n12699), .op(n6562) );
  nand2_1 U7269 ( .ip1(m1Inputs[22]), .ip2(n11974), .op(n6612) );
  nor3_1 U7270 ( .ip1(n10734), .ip2(n13835), .ip3(n6612), .op(n6566) );
  or2_1 U7271 ( .ip1(n6562), .ip2(n6566), .op(n6565) );
  or2_1 U7272 ( .ip1(n6563), .ip2(n6566), .op(n6564) );
  nand2_1 U7273 ( .ip1(n6565), .ip2(n6564), .op(n6602) );
  or2_1 U7274 ( .ip1(n6602), .ip2(n6566), .op(n6568) );
  nor2_1 U7275 ( .ip1(n10472), .ip2(n13594), .op(n6601) );
  or2_1 U7276 ( .ip1(n6601), .ip2(n6566), .op(n6567) );
  nand2_1 U7277 ( .ip1(n6568), .ip2(n6567), .op(n6622) );
  xnor2_1 U7278 ( .ip1(n6570), .ip2(n6569), .op(n6621) );
  xnor2_1 U7279 ( .ip1(n6572), .ip2(n6571), .op(n6620) );
  nand2_1 U7280 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[24]), .op(n6574)
         );
  nor3_1 U7281 ( .ip1(n10555), .ip2(n10753), .ip3(n6573), .op(n6578) );
  or2_1 U7282 ( .ip1(n6574), .ip2(n6578), .op(n6577) );
  or2_1 U7283 ( .ip1(n6575), .ip2(n6578), .op(n6576) );
  nand2_1 U7284 ( .ip1(n6577), .ip2(n6576), .op(n6651) );
  or2_1 U7285 ( .ip1(n6651), .ip2(n6578), .op(n6581) );
  nand2_1 U7286 ( .ip1(column[18]), .ip2(n13859), .op(n6650) );
  inv_1 U7287 ( .ip(n6650), .op(n6579) );
  or2_1 U7288 ( .ip1(n6579), .ip2(n6578), .op(n6580) );
  nand2_1 U7289 ( .ip1(n6581), .ip2(n6580), .op(n6628) );
  nor4_1 U7290 ( .ip1(n13646), .ip2(n13487), .ip3(n10827), .ip4(n10734), .op(
        n6586) );
  or2_1 U7291 ( .ip1(n6582), .ip2(n6586), .op(n6585) );
  or2_1 U7292 ( .ip1(n6583), .ip2(n6586), .op(n6584) );
  nand2_1 U7293 ( .ip1(n6585), .ip2(n6584), .op(n6669) );
  or2_1 U7294 ( .ip1(n6669), .ip2(n6586), .op(n6588) );
  nor2_1 U7295 ( .ip1(n9995), .ip2(n13594), .op(n6668) );
  or2_1 U7296 ( .ip1(n6668), .ip2(n6586), .op(n6587) );
  nand2_1 U7297 ( .ip1(n6588), .ip2(n6587), .op(n6627) );
  nand2_1 U7298 ( .ip1(m1Inputs[19]), .ip2(\STAGE_1/weightReg [8]), .op(n6626)
         );
  fulladder U7299 ( .a(n6591), .b(n6590), .ci(n6589), .co(n10697), .s(n6624)
         );
  nor2_1 U7300 ( .ip1(n6593), .ip2(n6592), .op(n6595) );
  xor2_1 U7301 ( .ip1(n6595), .ip2(n6594), .op(n6623) );
  fulladder U7302 ( .a(n6598), .b(n6597), .ci(n6596), .co(n10696), .s(n6659)
         );
  xor2_1 U7303 ( .ip1(n6600), .ip2(n6599), .op(n6667) );
  xor2_1 U7304 ( .ip1(n6602), .ip2(n6601), .op(n6666) );
  xor2_1 U7305 ( .ip1(n6604), .ip2(n6603), .op(n6665) );
  inv_1 U7306 ( .ip(n6605), .op(n6658) );
  and3_1 U7307 ( .ip1(m1Inputs[20]), .ip2(n14835), .ip3(n6675), .op(n6630) );
  or2_1 U7308 ( .ip1(n14835), .ip2(n6606), .op(n6608) );
  or2_1 U7309 ( .ip1(m1Inputs[19]), .ip2(n6606), .op(n6607) );
  nand2_1 U7310 ( .ip1(n6608), .ip2(n6607), .op(n6629) );
  nand2_1 U7311 ( .ip1(m1Inputs[18]), .ip2(n14975), .op(n6631) );
  nor2_1 U7312 ( .ip1(n6629), .ip2(n6631), .op(n6609) );
  nor2_1 U7313 ( .ip1(n6630), .ip2(n6609), .op(n6663) );
  nand2_1 U7314 ( .ip1(n14369), .ip2(m1Inputs[21]), .op(n6611) );
  nor3_1 U7315 ( .ip1(n10867), .ip2(n4624), .ip3(n6610), .op(n6615) );
  or2_1 U7316 ( .ip1(n6611), .ip2(n6615), .op(n6614) );
  or2_1 U7317 ( .ip1(n6612), .ip2(n6615), .op(n6613) );
  nand2_1 U7318 ( .ip1(n6614), .ip2(n6613), .op(n6638) );
  or2_1 U7319 ( .ip1(n6638), .ip2(n6615), .op(n6617) );
  nor2_1 U7320 ( .ip1(n10472), .ip2(n13766), .op(n6637) );
  or2_1 U7321 ( .ip1(n6637), .ip2(n6615), .op(n6616) );
  nand2_1 U7322 ( .ip1(n6617), .ip2(n6616), .op(n6662) );
  xor2_1 U7323 ( .ip1(n6619), .ip2(n6618), .op(n6661) );
  fulladder U7324 ( .a(n6622), .b(n6621), .ci(n6620), .co(n10695), .s(n6655)
         );
  fulladder U7325 ( .a(n6625), .b(n6624), .ci(n6623), .co(n10709), .s(n6654)
         );
  fulladder U7326 ( .a(n6628), .b(n6627), .ci(n6626), .co(n6625), .s(n6682) );
  nor2_1 U7327 ( .ip1(n6630), .ip2(n6629), .op(n6632) );
  xor2_1 U7328 ( .ip1(n6632), .ip2(n6631), .op(n6692) );
  nor2_1 U7329 ( .ip1(n6634), .ip2(n6633), .op(n6635) );
  nor2_1 U7330 ( .ip1(n6636), .ip2(n6635), .op(n6691) );
  xnor2_1 U7331 ( .ip1(n6638), .ip2(n6637), .op(n6690) );
  or2_1 U7332 ( .ip1(n6639), .ip2(n6640), .op(n6643) );
  or2_1 U7333 ( .ip1(n6641), .ip2(n6640), .op(n6642) );
  nand2_1 U7334 ( .ip1(n6643), .ip2(n6642), .op(n6689) );
  or2_1 U7335 ( .ip1(n6644), .ip2(n6646), .op(n6649) );
  inv_1 U7336 ( .ip(n6645), .op(n6647) );
  or2_1 U7337 ( .ip1(n6647), .ip2(n6646), .op(n6648) );
  nand2_1 U7338 ( .ip1(n6649), .ip2(n6648), .op(n6688) );
  xor2_1 U7339 ( .ip1(n6651), .ip2(n6650), .op(n6687) );
  inv_1 U7340 ( .ip(n6652), .op(n10716) );
  fulladder U7341 ( .a(n6655), .b(n6654), .ci(n6653), .co(n10718), .s(n6656)
         );
  inv_1 U7342 ( .ip(n6656), .op(n6679) );
  fulladder U7343 ( .a(n6659), .b(n6658), .ci(n6657), .co(n10708), .s(n6660)
         );
  inv_1 U7344 ( .ip(n6660), .op(n6678) );
  fulladder U7345 ( .a(n6663), .b(n6662), .ci(n6661), .co(n6657), .s(n6664) );
  inv_1 U7346 ( .ip(n6664), .op(n6685) );
  fulladder U7347 ( .a(n6667), .b(n6666), .ci(n6665), .co(n6605), .s(n6684) );
  xor2_1 U7348 ( .ip1(n6669), .ip2(n6668), .op(n6703) );
  fulladder U7349 ( .a(n6672), .b(n6671), .ci(n6670), .co(n6673), .s(n5927) );
  inv_1 U7350 ( .ip(n6673), .op(n6702) );
  fulladder U7351 ( .a(n6676), .b(n6675), .ci(n6674), .co(n6701), .s(n6710) );
  fulladder U7352 ( .a(n6679), .b(n6678), .ci(n6677), .co(n10715), .s(n6722)
         );
  fulladder U7353 ( .a(n6682), .b(n6681), .ci(n6680), .co(n6653), .s(n6699) );
  fulladder U7354 ( .a(n6685), .b(n6684), .ci(n6683), .co(n6677), .s(n6686) );
  inv_1 U7355 ( .ip(n6686), .op(n6698) );
  fulladder U7356 ( .a(n6689), .b(n6688), .ci(n6687), .co(n6680), .s(n6706) );
  fulladder U7357 ( .a(n6692), .b(n6691), .ci(n6690), .co(n6681), .s(n6705) );
  fulladder U7358 ( .a(n6695), .b(n6694), .ci(n6693), .co(n6704), .s(n5915) );
  inv_1 U7359 ( .ip(n6696), .op(n6721) );
  fulladder U7360 ( .a(n6699), .b(n6698), .ci(n6697), .co(n6696), .s(n6700) );
  inv_1 U7361 ( .ip(n6700), .op(n6725) );
  fulladder U7362 ( .a(n6703), .b(n6702), .ci(n6701), .co(n6683), .s(n6713) );
  fulladder U7363 ( .a(n6706), .b(n6705), .ci(n6704), .co(n6697), .s(n6707) );
  inv_1 U7364 ( .ip(n6707), .op(n6712) );
  fulladder U7365 ( .a(n6710), .b(n6709), .ci(n6708), .co(n6711), .s(n6718) );
  fulladder U7366 ( .a(n6713), .b(n6712), .ci(n6711), .co(n6724), .s(n6728) );
  fulladder U7367 ( .a(n6716), .b(n6715), .ci(n6714), .co(n6727), .s(
        \STAGE_1/M2/sum [1]) );
  fulladder U7368 ( .a(n6719), .b(n6718), .ci(n6717), .co(n6726), .s(n6716) );
  fulladder U7369 ( .a(n6722), .b(n6721), .ci(n6720), .co(n10714), .s(
        \STAGE_1/M2/sum [4]) );
  fulladder U7370 ( .a(n6725), .b(n6724), .ci(n6723), .co(n6720), .s(
        \STAGE_1/M2/sum [3]) );
  fulladder U7371 ( .a(n6728), .b(n6727), .ci(n6726), .co(n6723), .s(
        \STAGE_1/M2/sum [2]) );
  nand2_1 U7372 ( .ip1(m1Inputs[52]), .ip2(n12699), .op(n6730) );
  nor3_1 U7373 ( .ip1(n8942), .ip2(n12255), .ip3(n6729), .op(n6822) );
  or2_1 U7374 ( .ip1(n6730), .ip2(n6822), .op(n6732) );
  nand2_1 U7375 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[53]), .op(n6816)
         );
  or2_1 U7376 ( .ip1(n6816), .ip2(n6822), .op(n6731) );
  nand2_1 U7377 ( .ip1(n6732), .ip2(n6731), .op(n6821) );
  nor2_1 U7378 ( .ip1(n12126), .ip2(n6503), .op(n6823) );
  xnor2_1 U7379 ( .ip1(n6821), .ip2(n6823), .op(n6904) );
  and3_1 U7380 ( .ip1(n12578), .ip2(m1Inputs[57]), .ip3(n6733), .op(n6815) );
  inv_1 U7381 ( .ip(m1Inputs[57]), .op(n12231) );
  nor2_1 U7382 ( .ip1(n13646), .ip2(n12231), .op(n6734) );
  or2_1 U7383 ( .ip1(m1Inputs[54]), .ip2(n6734), .op(n6736) );
  or2_1 U7384 ( .ip1(n9733), .ip2(n6734), .op(n6735) );
  nand2_1 U7385 ( .ip1(n6736), .ip2(n6735), .op(n6813) );
  nor2_1 U7386 ( .ip1(n6815), .ip2(n6813), .op(n6737) );
  nand2_1 U7387 ( .ip1(m1Inputs[48]), .ip2(n14994), .op(n6812) );
  xor2_1 U7388 ( .ip1(n6737), .ip2(n6812), .op(n6903) );
  fulladder U7389 ( .a(n6740), .b(n6739), .ci(n6738), .co(n6902), .s(n5157) );
  inv_1 U7390 ( .ip(n6741), .op(n6928) );
  nor2_1 U7391 ( .ip1(n12032), .ip2(n14368), .op(n6888) );
  nor2_1 U7392 ( .ip1(n12138), .ip2(n14289), .op(n6887) );
  nand3_1 U7393 ( .ip1(column[48]), .ip2(n15042), .ip3(n6742), .op(n6743) );
  nand2_1 U7394 ( .ip1(n6744), .ip2(n6743), .op(n6886) );
  nand2_1 U7395 ( .ip1(n12809), .ip2(m1Inputs[56]), .op(n6780) );
  inv_1 U7396 ( .ip(m1Inputs[56]), .op(n12237) );
  nor4_1 U7397 ( .ip1(n6745), .ip2(n9047), .ip3(n12237), .ip4(n12155), .op(
        n6828) );
  or2_1 U7398 ( .ip1(n6780), .ip2(n6828), .op(n6748) );
  nand2_1 U7399 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[55]), .op(n6746)
         );
  or2_1 U7400 ( .ip1(n6746), .ip2(n6828), .op(n6747) );
  nand2_1 U7401 ( .ip1(n6748), .ip2(n6747), .op(n6826) );
  nand2_1 U7402 ( .ip1(column[49]), .ip2(n14768), .op(n6827) );
  xor2_1 U7403 ( .ip1(n6826), .ip2(n6827), .op(n6884) );
  inv_1 U7404 ( .ip(n6749), .op(n6751) );
  nor2_1 U7405 ( .ip1(n6751), .ip2(n6750), .op(n6883) );
  nor2_1 U7406 ( .ip1(n6753), .ip2(n6752), .op(n6882) );
  inv_1 U7407 ( .ip(n6754), .op(n6918) );
  fulladder U7408 ( .a(n6757), .b(n6756), .ci(n6755), .co(n6917), .s(n6761) );
  fulladder U7409 ( .a(n6760), .b(n6759), .ci(n6758), .co(n6926), .s(n6762) );
  fulladder U7410 ( .a(n6763), .b(n6762), .ci(n6761), .co(n6924), .s(n6766) );
  fulladder U7411 ( .a(n6766), .b(n6765), .ci(n6764), .co(n6923), .s(
        \STAGE_1/M4/sum [0]) );
  nand2_1 U7412 ( .ip1(m1Inputs[54]), .ip2(n12699), .op(n6767) );
  nand2_1 U7413 ( .ip1(m1Inputs[54]), .ip2(\STAGE_1/weightReg [4]), .op(n6818)
         );
  nor3_1 U7414 ( .ip1(n12155), .ip2(n13835), .ip3(n6818), .op(n6770) );
  or2_1 U7415 ( .ip1(n6767), .ip2(n6770), .op(n6769) );
  nand2_1 U7416 ( .ip1(m1Inputs[55]), .ip2(\STAGE_1/weightReg [4]), .op(n6773)
         );
  or2_1 U7417 ( .ip1(n6773), .ip2(n6770), .op(n6768) );
  nand2_1 U7418 ( .ip1(n6769), .ip2(n6768), .op(n6857) );
  or2_1 U7419 ( .ip1(n6857), .ip2(n6770), .op(n6772) );
  nor2_1 U7420 ( .ip1(n12126), .ip2(n13390), .op(n6856) );
  or2_1 U7421 ( .ip1(n6856), .ip2(n6770), .op(n6771) );
  nand2_1 U7422 ( .ip1(n6772), .ip2(n6771), .op(n11891) );
  nand2_1 U7423 ( .ip1(m1Inputs[55]), .ip2(n12699), .op(n6774) );
  nor3_1 U7424 ( .ip1(n12237), .ip2(n13835), .ip3(n6773), .op(n11842) );
  or2_1 U7425 ( .ip1(n6774), .ip2(n11842), .op(n6776) );
  nand2_1 U7426 ( .ip1(m1Inputs[56]), .ip2(n11974), .op(n11859) );
  or2_1 U7427 ( .ip1(n11859), .ip2(n11842), .op(n6775) );
  nand2_1 U7428 ( .ip1(n6776), .ip2(n6775), .op(n11841) );
  nor2_1 U7429 ( .ip1(n12126), .ip2(n13579), .op(n11843) );
  xnor2_1 U7430 ( .ip1(n11841), .ip2(n11843), .op(n11890) );
  nand2_1 U7431 ( .ip1(n14835), .ip2(m1Inputs[53]), .op(n6777) );
  nand2_1 U7432 ( .ip1(n13749), .ip2(m1Inputs[53]), .op(n6844) );
  nor3_1 U7433 ( .ip1(n12063), .ip2(n14384), .ip3(n6844), .op(n11875) );
  or2_1 U7434 ( .ip1(n6777), .ip2(n11875), .op(n6779) );
  nand2_1 U7435 ( .ip1(m1Inputs[54]), .ip2(n12981), .op(n11863) );
  or2_1 U7436 ( .ip1(n11863), .ip2(n11875), .op(n6778) );
  nand2_1 U7437 ( .ip1(n6779), .ip2(n6778), .op(n11874) );
  nor2_1 U7438 ( .ip1(n12032), .ip2(n13390), .op(n11876) );
  xnor2_1 U7439 ( .ip1(n11874), .ip2(n11876), .op(n11889) );
  nand2_1 U7440 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[56]), .op(n6781)
         );
  nor3_1 U7441 ( .ip1(n13854), .ip2(n12231), .ip3(n6780), .op(n6784) );
  or2_1 U7442 ( .ip1(n6781), .ip2(n6784), .op(n6783) );
  nand2_1 U7443 ( .ip1(n12809), .ip2(m1Inputs[57]), .op(n6794) );
  or2_1 U7444 ( .ip1(n6794), .ip2(n6784), .op(n6782) );
  nand2_1 U7445 ( .ip1(n6783), .ip2(n6782), .op(n6833) );
  or2_1 U7446 ( .ip1(n6833), .ip2(n6784), .op(n6787) );
  nand2_1 U7447 ( .ip1(column[50]), .ip2(n13039), .op(n6832) );
  inv_1 U7448 ( .ip(n6832), .op(n6785) );
  or2_1 U7449 ( .ip1(n6785), .ip2(n6784), .op(n6786) );
  nand2_1 U7450 ( .ip1(n6787), .ip2(n6786), .op(n6808) );
  nand2_1 U7451 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[58]), .op(n11853) );
  inv_1 U7452 ( .ip(m1Inputs[58]), .op(n12230) );
  nor4_1 U7453 ( .ip1(n10476), .ip2(n13801), .ip3(n12230), .ip4(n12155), .op(
        n6791) );
  or2_1 U7454 ( .ip1(n11853), .ip2(n6791), .op(n6790) );
  or2_1 U7455 ( .ip1(n6788), .ip2(n6791), .op(n6789) );
  nand2_1 U7456 ( .ip1(n6790), .ip2(n6789), .op(n6881) );
  or2_1 U7457 ( .ip1(n6881), .ip2(n6791), .op(n6793) );
  nor2_1 U7458 ( .ip1(n11858), .ip2(n13594), .op(n6880) );
  or2_1 U7459 ( .ip1(n6880), .ip2(n6791), .op(n6792) );
  nand2_1 U7460 ( .ip1(n6793), .ip2(n6792), .op(n6807) );
  nand2_1 U7461 ( .ip1(m1Inputs[51]), .ip2(n14975), .op(n6806) );
  nand2_1 U7462 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[52]), .op(n11885) );
  nand2_1 U7463 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[57]), .op(n6795)
         );
  nor3_1 U7464 ( .ip1(n13709), .ip2(n12230), .ip3(n6794), .op(n6798) );
  or2_1 U7465 ( .ip1(n6795), .ip2(n6798), .op(n6797) );
  nand2_1 U7466 ( .ip1(n13707), .ip2(m1Inputs[58]), .op(n6850) );
  or2_1 U7467 ( .ip1(n6850), .ip2(n6798), .op(n6796) );
  nand2_1 U7468 ( .ip1(n6797), .ip2(n6796), .op(n6871) );
  or2_1 U7469 ( .ip1(n6871), .ip2(n6798), .op(n6801) );
  nand2_1 U7470 ( .ip1(column[51]), .ip2(n13039), .op(n6870) );
  inv_1 U7471 ( .ip(n6870), .op(n6799) );
  or2_1 U7472 ( .ip1(n6799), .ip2(n6798), .op(n6800) );
  nand2_1 U7473 ( .ip1(n6801), .ip2(n6800), .op(n11884) );
  nand2_1 U7474 ( .ip1(m1Inputs[51]), .ip2(n14994), .op(n11883) );
  nand2_1 U7475 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[60]), .op(n12212) );
  nor3_1 U7476 ( .ip1(n13646), .ip2(n12231), .ip3(n12212), .op(n11849) );
  nor2_1 U7477 ( .ip1(n13082), .ip2(n12231), .op(n6802) );
  or2_1 U7478 ( .ip1(m1Inputs[60]), .ip2(n6802), .op(n6804) );
  or2_1 U7479 ( .ip1(n13803), .ip2(n6802), .op(n6803) );
  nand2_1 U7480 ( .ip1(n6804), .ip2(n6803), .op(n11847) );
  nor2_1 U7481 ( .ip1(n11849), .ip2(n11847), .op(n6805) );
  nand2_1 U7482 ( .ip1(m1Inputs[48]), .ip2(n15025), .op(n11846) );
  xor2_1 U7483 ( .ip1(n6805), .ip2(n11846), .op(n11892) );
  fulladder U7484 ( .a(n6808), .b(n6807), .ci(n6806), .co(n11894), .s(n6891)
         );
  and3_1 U7485 ( .ip1(m1Inputs[52]), .ip2(n14835), .ip3(n6887), .op(n6864) );
  nor2_1 U7486 ( .ip1(n12066), .ip2(n14289), .op(n6842) );
  or2_1 U7487 ( .ip1(n14835), .ip2(n6842), .op(n6810) );
  or2_1 U7488 ( .ip1(m1Inputs[51]), .ip2(n6842), .op(n6809) );
  nand2_1 U7489 ( .ip1(n6810), .ip2(n6809), .op(n6862) );
  nor2_1 U7490 ( .ip1(n6864), .ip2(n6862), .op(n6811) );
  nand2_1 U7491 ( .ip1(m1Inputs[50]), .ip2(n14975), .op(n6861) );
  xor2_1 U7492 ( .ip1(n6811), .ip2(n6861), .op(n6901) );
  nor2_1 U7493 ( .ip1(n6813), .ip2(n6812), .op(n6814) );
  nor2_1 U7494 ( .ip1(n6815), .ip2(n6814), .op(n6900) );
  nand2_1 U7495 ( .ip1(n14369), .ip2(m1Inputs[53]), .op(n6817) );
  nor3_1 U7496 ( .ip1(n12063), .ip2(n13835), .ip3(n6816), .op(n6866) );
  or2_1 U7497 ( .ip1(n6817), .ip2(n6866), .op(n6820) );
  or2_1 U7498 ( .ip1(n6818), .ip2(n6866), .op(n6819) );
  nand2_1 U7499 ( .ip1(n6820), .ip2(n6819), .op(n6865) );
  nor2_1 U7500 ( .ip1(n12126), .ip2(n12083), .op(n6867) );
  xnor2_1 U7501 ( .ip1(n6865), .ip2(n6867), .op(n6899) );
  or2_1 U7502 ( .ip1(n6821), .ip2(n6822), .op(n6825) );
  or2_1 U7503 ( .ip1(n6823), .ip2(n6822), .op(n6824) );
  nand2_1 U7504 ( .ip1(n6825), .ip2(n6824), .op(n6898) );
  or2_1 U7505 ( .ip1(n6826), .ip2(n6828), .op(n6831) );
  inv_1 U7506 ( .ip(n6827), .op(n6829) );
  or2_1 U7507 ( .ip1(n6829), .ip2(n6828), .op(n6830) );
  nand2_1 U7508 ( .ip1(n6831), .ip2(n6830), .op(n6897) );
  xor2_1 U7509 ( .ip1(n6833), .ip2(n6832), .op(n6896) );
  inv_1 U7510 ( .ip(n6834), .op(n11904) );
  nand2_1 U7511 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[56]), .op(n6836)
         );
  inv_1 U7512 ( .ip(m1Inputs[59]), .op(n12248) );
  nor3_1 U7513 ( .ip1(n13082), .ip2(n12248), .ip3(n6835), .op(n6839) );
  or2_1 U7514 ( .ip1(n6836), .ip2(n6839), .op(n6838) );
  nand2_1 U7515 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[59]), .op(n12247) );
  or2_1 U7516 ( .ip1(n12247), .ip2(n6839), .op(n6837) );
  nand2_1 U7517 ( .ip1(n6838), .ip2(n6837), .op(n6859) );
  or2_1 U7518 ( .ip1(n6859), .ip2(n6839), .op(n6841) );
  nor2_1 U7519 ( .ip1(n11858), .ip2(n13579), .op(n6858) );
  or2_1 U7520 ( .ip1(n6858), .ip2(n6839), .op(n6840) );
  nand2_1 U7521 ( .ip1(n6841), .ip2(n6840), .op(n11888) );
  nand2_1 U7522 ( .ip1(m1Inputs[52]), .ip2(n4627), .op(n6843) );
  and3_1 U7523 ( .ip1(n4627), .ip2(m1Inputs[53]), .ip3(n6842), .op(n6847) );
  or2_1 U7524 ( .ip1(n6843), .ip2(n6847), .op(n6846) );
  or2_1 U7525 ( .ip1(n6844), .ip2(n6847), .op(n6845) );
  nand2_1 U7526 ( .ip1(n6846), .ip2(n6845), .op(n6855) );
  or2_1 U7527 ( .ip1(n6855), .ip2(n6847), .op(n6849) );
  nor2_1 U7528 ( .ip1(n12032), .ip2(n13766), .op(n6854) );
  or2_1 U7529 ( .ip1(n6854), .ip2(n6847), .op(n6848) );
  nand2_1 U7530 ( .ip1(n6849), .ip2(n6848), .op(n11887) );
  nand2_1 U7531 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[58]), .op(n6851)
         );
  nor3_1 U7532 ( .ip1(n13709), .ip2(n12248), .ip3(n6850), .op(n11870) );
  or2_1 U7533 ( .ip1(n6851), .ip2(n11870), .op(n6853) );
  nand2_1 U7534 ( .ip1(n12809), .ip2(m1Inputs[59]), .op(n11879) );
  or2_1 U7535 ( .ip1(n11879), .ip2(n11870), .op(n6852) );
  nand2_1 U7536 ( .ip1(n6853), .ip2(n6852), .op(n11868) );
  nand2_1 U7537 ( .ip1(column[52]), .ip2(n13039), .op(n11869) );
  xor2_1 U7538 ( .ip1(n11868), .ip2(n11869), .op(n11886) );
  xor2_1 U7539 ( .ip1(n6855), .ip2(n6854), .op(n6879) );
  xor2_1 U7540 ( .ip1(n6857), .ip2(n6856), .op(n6878) );
  xor2_1 U7541 ( .ip1(n6859), .ip2(n6858), .op(n6877) );
  inv_1 U7542 ( .ip(n6860), .op(n11896) );
  nor2_1 U7543 ( .ip1(n6862), .ip2(n6861), .op(n6863) );
  nor2_1 U7544 ( .ip1(n6864), .ip2(n6863), .op(n6875) );
  or2_1 U7545 ( .ip1(n6865), .ip2(n6866), .op(n6869) );
  or2_1 U7546 ( .ip1(n6867), .ip2(n6866), .op(n6868) );
  nand2_1 U7547 ( .ip1(n6869), .ip2(n6868), .op(n6874) );
  xor2_1 U7548 ( .ip1(n6871), .ip2(n6870), .op(n6873) );
  inv_1 U7549 ( .ip(n6872), .op(n11903) );
  fulladder U7550 ( .a(n6875), .b(n6874), .ci(n6873), .co(n11895), .s(n6876)
         );
  inv_1 U7551 ( .ip(n6876), .op(n6894) );
  fulladder U7552 ( .a(n6879), .b(n6878), .ci(n6877), .co(n6860), .s(n6893) );
  xor2_1 U7553 ( .ip1(n6881), .ip2(n6880), .op(n6912) );
  fulladder U7554 ( .a(n6884), .b(n6883), .ci(n6882), .co(n6885), .s(n6754) );
  inv_1 U7555 ( .ip(n6885), .op(n6911) );
  fulladder U7556 ( .a(n6888), .b(n6887), .ci(n6886), .co(n6910), .s(n6919) );
  fulladder U7557 ( .a(n6891), .b(n6890), .ci(n6889), .co(n11898), .s(n6908)
         );
  fulladder U7558 ( .a(n6894), .b(n6893), .ci(n6892), .co(n11902), .s(n6895)
         );
  inv_1 U7559 ( .ip(n6895), .op(n6907) );
  fulladder U7560 ( .a(n6898), .b(n6897), .ci(n6896), .co(n6889), .s(n6915) );
  fulladder U7561 ( .a(n6901), .b(n6900), .ci(n6899), .co(n6890), .s(n6914) );
  fulladder U7562 ( .a(n6904), .b(n6903), .ci(n6902), .co(n6913), .s(n6741) );
  inv_1 U7563 ( .ip(n6905), .op(n11906) );
  fulladder U7564 ( .a(n6908), .b(n6907), .ci(n6906), .co(n6905), .s(n6909) );
  inv_1 U7565 ( .ip(n6909), .op(n6931) );
  fulladder U7566 ( .a(n6912), .b(n6911), .ci(n6910), .co(n6892), .s(n6922) );
  fulladder U7567 ( .a(n6915), .b(n6914), .ci(n6913), .co(n6906), .s(n6916) );
  inv_1 U7568 ( .ip(n6916), .op(n6921) );
  fulladder U7569 ( .a(n6919), .b(n6918), .ci(n6917), .co(n6920), .s(n6927) );
  fulladder U7570 ( .a(n6922), .b(n6921), .ci(n6920), .co(n6930), .s(n6934) );
  fulladder U7571 ( .a(n6925), .b(n6924), .ci(n6923), .co(n6933), .s(
        \STAGE_1/M4/sum [1]) );
  fulladder U7572 ( .a(n6928), .b(n6927), .ci(n6926), .co(n6932), .s(n6925) );
  fulladder U7573 ( .a(n6931), .b(n6930), .ci(n6929), .co(n11905), .s(
        \STAGE_1/M4/sum [3]) );
  fulladder U7574 ( .a(n6934), .b(n6933), .ci(n6932), .co(n6929), .s(
        \STAGE_1/M4/sum [2]) );
  nand2_1 U7575 ( .ip1(n11974), .ip2(m1Inputs[101]), .op(n7558) );
  nor4_1 U7576 ( .ip1(n14783), .ip2(n7553), .ip3(n13835), .ip4(n7326), .op(
        n7597) );
  or2_1 U7577 ( .ip1(n7558), .ip2(n7597), .op(n6937) );
  or2_1 U7578 ( .ip1(n6935), .ip2(n7597), .op(n6936) );
  nand2_1 U7579 ( .ip1(n6937), .ip2(n6936), .op(n7596) );
  nor2_1 U7580 ( .ip1(n7564), .ip2(n6503), .op(n7598) );
  xnor2_1 U7581 ( .ip1(n7596), .ip2(n7598), .op(n7654) );
  and3_1 U7582 ( .ip1(n12578), .ip2(m1Inputs[105]), .ip3(n6938), .op(n7593) );
  inv_1 U7583 ( .ip(m1Inputs[105]), .op(n7518) );
  nor2_1 U7584 ( .ip1(n10476), .ip2(n7518), .op(n6939) );
  or2_1 U7585 ( .ip1(m1Inputs[102]), .ip2(n6939), .op(n6941) );
  or2_1 U7586 ( .ip1(n9733), .ip2(n6939), .op(n6940) );
  nand2_1 U7587 ( .ip1(n6941), .ip2(n6940), .op(n7591) );
  nor2_1 U7588 ( .ip1(n7593), .ip2(n7591), .op(n6942) );
  nand2_1 U7589 ( .ip1(m1Inputs[96]), .ip2(\STAGE_1/weightReg [9]), .op(n7590)
         );
  xor2_1 U7590 ( .ip1(n6942), .ip2(n7590), .op(n7653) );
  fulladder U7591 ( .a(n6945), .b(n6944), .ci(n6943), .co(n7652), .s(n5034) );
  inv_1 U7592 ( .ip(n6946), .op(n7679) );
  inv_1 U7593 ( .ip(n6947), .op(n6951) );
  nor2_1 U7594 ( .ip1(n6949), .ip2(n6948), .op(n6950) );
  nor2_1 U7595 ( .ip1(n6951), .ip2(n6950), .op(n7634) );
  nand2_1 U7596 ( .ip1(m1Inputs[99]), .ip2(n12981), .op(n7633) );
  nand2_1 U7597 ( .ip1(m1Inputs[98]), .ip2(\STAGE_1/weightReg [7]), .op(n7632)
         );
  inv_1 U7598 ( .ip(n6952), .op(n7670) );
  or2_1 U7599 ( .ip1(n6953), .ip2(n6954), .op(n6957) );
  or2_1 U7600 ( .ip1(n6955), .ip2(n6954), .op(n6956) );
  nand2_1 U7601 ( .ip1(n6957), .ip2(n6956), .op(n7631) );
  or2_1 U7602 ( .ip1(n6958), .ip2(n6959), .op(n6962) );
  or2_1 U7603 ( .ip1(n6960), .ip2(n6959), .op(n6961) );
  nand2_1 U7604 ( .ip1(n6962), .ip2(n6961), .op(n7630) );
  nand2_1 U7605 ( .ip1(n4619), .ip2(m1Inputs[103]), .op(n6964) );
  nor3_1 U7606 ( .ip1(n13709), .ip2(n14169), .ip3(n6963), .op(n7603) );
  or2_1 U7607 ( .ip1(n6964), .ip2(n7603), .op(n6966) );
  nand2_1 U7608 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[104]), .op(n7517) );
  or2_1 U7609 ( .ip1(n7517), .ip2(n7603), .op(n6965) );
  nand2_1 U7610 ( .ip1(n6966), .ip2(n6965), .op(n7601) );
  nand2_1 U7611 ( .ip1(column[97]), .ip2(n13498), .op(n7602) );
  xor2_1 U7612 ( .ip1(n7601), .ip2(n7602), .op(n7629) );
  inv_1 U7613 ( .ip(n6967), .op(n7669) );
  fulladder U7614 ( .a(n6970), .b(n6969), .ci(n6968), .co(n7668), .s(n6974) );
  fulladder U7615 ( .a(n6973), .b(n6972), .ci(n6971), .co(n7677), .s(n6975) );
  fulladder U7616 ( .a(n6976), .b(n6975), .ci(n6974), .co(n7675), .s(n6979) );
  fulladder U7617 ( .a(n6979), .b(n6978), .ci(n6977), .co(n7674), .s(
        \STAGE_1/M7/sum [0]) );
  buf_1 U7618 ( .ip(n14340), .op(n14373) );
  nand2_1 U7619 ( .ip1(m1Inputs[103]), .ip2(\STAGE_1/weightReg [13]), .op(
        n6981) );
  inv_1 U7620 ( .ip(n14824), .op(n14847) );
  buf_1 U7621 ( .ip(n14847), .op(n13718) );
  nand2_1 U7622 ( .ip1(m1Inputs[105]), .ip2(\STAGE_1/weightReg [11]), .op(
        n6980) );
  xor2_1 U7623 ( .ip1(n6981), .ip2(n6980), .op(n7036) );
  inv_1 U7624 ( .ip(\STAGE_1/weightReg [14]), .op(n14842) );
  nor2_1 U7625 ( .ip1(n14842), .ip2(n7559), .op(n6982) );
  xor2_1 U7626 ( .ip1(n7036), .ip2(n6982), .op(n7030) );
  nor2_1 U7627 ( .ip1(n14188), .ip2(n14169), .op(n7047) );
  nand3_1 U7628 ( .ip1(n14847), .ip2(m1Inputs[103]), .ip3(n7047), .op(n6986)
         );
  buf_1 U7629 ( .ip(n14842), .op(n14883) );
  inv_1 U7630 ( .ip(n14883), .op(n14816) );
  nand2_1 U7631 ( .ip1(m1Inputs[103]), .ip2(\STAGE_1/weightReg [12]), .op(
        n6984) );
  nand2_1 U7632 ( .ip1(m1Inputs[104]), .ip2(\STAGE_1/weightReg [11]), .op(
        n6983) );
  xor2_1 U7633 ( .ip1(n6984), .ip2(n6983), .op(n7058) );
  nand3_1 U7634 ( .ip1(n14816), .ip2(n7058), .ip3(m1Inputs[101]), .op(n6985)
         );
  nand2_1 U7635 ( .ip1(n6986), .ip2(n6985), .op(n7029) );
  inv_1 U7636 ( .ip(m1Inputs[108]), .op(n7331) );
  nor2_1 U7637 ( .ip1(n7331), .ip2(n14384), .op(n7061) );
  inv_1 U7638 ( .ip(m1Inputs[110]), .op(n14189) );
  nor2_1 U7639 ( .ip1(n14189), .ip2(n12746), .op(n7060) );
  nand2_1 U7640 ( .ip1(m1Inputs[111]), .ip2(n13637), .op(n7059) );
  inv_1 U7641 ( .ip(m1Inputs[109]), .op(n14170) );
  nor2_1 U7642 ( .ip1(n14170), .ip2(n14368), .op(n7048) );
  inv_1 U7643 ( .ip(\STAGE_1/weightReg [15]), .op(n14853) );
  inv_1 U7644 ( .ip(n14853), .op(n14976) );
  nand2_1 U7645 ( .ip1(n14976), .ip2(m1Inputs[101]), .op(n7046) );
  inv_1 U7646 ( .ip(n6987), .op(n7052) );
  nor2_1 U7647 ( .ip1(n14189), .ip2(n14289), .op(n7034) );
  nor2_1 U7648 ( .ip1(n6504), .ip2(n7331), .op(n7033) );
  nand2_1 U7649 ( .ip1(m1Inputs[111]), .ip2(n14369), .op(n7032) );
  inv_1 U7650 ( .ip(n6988), .op(n7051) );
  nand2_1 U7651 ( .ip1(n14629), .ip2(m1Inputs[106]), .op(n7039) );
  nand2_1 U7652 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[104]), .op(n7209) );
  nor2_1 U7653 ( .ip1(n7039), .ip2(n7209), .op(n6992) );
  nand2_1 U7654 ( .ip1(m1Inputs[106]), .ip2(n14975), .op(n6990) );
  nand2_1 U7655 ( .ip1(m1Inputs[104]), .ip2(\STAGE_1/weightReg [10]), .op(
        n6989) );
  xor2_1 U7656 ( .ip1(n6990), .ip2(n6989), .op(n7006) );
  and3_1 U7657 ( .ip1(column[106]), .ip2(n13498), .ip3(n7006), .op(n6991) );
  nor2_1 U7658 ( .ip1(n6992), .ip2(n6991), .op(n7010) );
  nand2_1 U7659 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[102]), .op(
        n7009) );
  nand2_1 U7660 ( .ip1(n13718), .ip2(m1Inputs[108]), .op(n14259) );
  nand2_1 U7661 ( .ip1(m1Inputs[103]), .ip2(n12981), .op(n7311) );
  nor2_1 U7662 ( .ip1(n14259), .ip2(n7311), .op(n6997) );
  inv_1 U7663 ( .ip(m1Inputs[103]), .op(n7492) );
  nor2_1 U7664 ( .ip1(n13579), .ip2(n7492), .op(n7078) );
  or2_1 U7665 ( .ip1(n13749), .ip2(n7078), .op(n6994) );
  or2_1 U7666 ( .ip1(m1Inputs[108]), .ip2(n7078), .op(n6993) );
  nand2_1 U7667 ( .ip1(n6994), .ip2(n6993), .op(n6995) );
  or2_1 U7668 ( .ip1(n6997), .ip2(n6995), .op(n7076) );
  nor3_1 U7669 ( .ip1(n14842), .ip2(n7553), .ip3(n7076), .op(n6996) );
  nor2_1 U7670 ( .ip1(n6997), .ip2(n6996), .op(n7008) );
  inv_1 U7671 ( .ip(n6998), .op(n7126) );
  inv_1 U7672 ( .ip(m1Inputs[106]), .op(n14187) );
  nand2_1 U7673 ( .ip1(m1Inputs[107]), .ip2(n4627), .op(n7113) );
  nor3_1 U7674 ( .ip1(n14187), .ip2(n14289), .ip3(n7113), .op(n7004) );
  inv_1 U7675 ( .ip(n7004), .op(n7002) );
  nand2_1 U7676 ( .ip1(m1Inputs[107]), .ip2(n12981), .op(n7000) );
  nand2_1 U7677 ( .ip1(m1Inputs[106]), .ip2(\STAGE_1/weightReg [7]), .op(n6999) );
  nand2_1 U7678 ( .ip1(n7000), .ip2(n6999), .op(n7001) );
  nand2_1 U7679 ( .ip1(n7002), .ip2(n7001), .op(n7099) );
  nor3_1 U7680 ( .ip1(n7331), .ip2(n4624), .ip3(n7099), .op(n7003) );
  nor2_1 U7681 ( .ip1(n7004), .ip2(n7003), .op(n7137) );
  nand2_1 U7682 ( .ip1(m1Inputs[109]), .ip2(n13637), .op(n7143) );
  nor2_1 U7683 ( .ip1(n7486), .ip2(n14853), .op(n7142) );
  nand2_1 U7684 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[105]), .op(n7141) );
  nand2_1 U7685 ( .ip1(column[106]), .ip2(n14768), .op(n7005) );
  xor2_1 U7686 ( .ip1(n7006), .ip2(n7005), .op(n7135) );
  inv_1 U7687 ( .ip(n7007), .op(n7090) );
  fulladder U7688 ( .a(n7010), .b(n7009), .ci(n7008), .co(n7050), .s(n7011) );
  inv_1 U7689 ( .ip(n7011), .op(n7089) );
  nor2_1 U7690 ( .ip1(n14902), .ip2(n7559), .op(n7093) );
  nor2_1 U7691 ( .ip1(n14340), .ip2(n7326), .op(n7092) );
  and2_1 U7692 ( .ip1(column[105]), .ip2(n13498), .op(n7103) );
  nand2_1 U7693 ( .ip1(column[104]), .ip2(n13498), .op(n7177) );
  inv_1 U7694 ( .ip(n7177), .op(n7102) );
  nor2_1 U7695 ( .ip1(n12083), .ip2(n14169), .op(n7101) );
  nor2_1 U7696 ( .ip1(n14842), .ip2(n7492), .op(n14186) );
  nor2_1 U7697 ( .ip1(n14373), .ip2(n14169), .op(n14185) );
  nand4_1 U7698 ( .ip1(\STAGE_1/weightReg [10]), .ip2(n14994), .ip3(
        m1Inputs[107]), .ip4(m1Inputs[106]), .op(n7017) );
  inv_1 U7699 ( .ip(n7017), .op(n7012) );
  or2_1 U7700 ( .ip1(n7039), .ip2(n7012), .op(n7015) );
  nand2_1 U7701 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[107]), .op(n7013) );
  or2_1 U7702 ( .ip1(n7013), .ip2(n7012), .op(n7014) );
  nand2_1 U7703 ( .ip1(n7015), .ip2(n7014), .op(n7026) );
  nand3_1 U7704 ( .ip1(column[108]), .ip2(n15042), .ip3(n7026), .op(n7016) );
  nand2_1 U7705 ( .ip1(n7017), .ip2(n7016), .op(n14184) );
  nand2_1 U7706 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[105]), .op(n7117) );
  nor2_1 U7707 ( .ip1(n7039), .ip2(n7117), .op(n7019) );
  inv_1 U7708 ( .ip(n7019), .op(n7024) );
  nand2_1 U7709 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[106]), .op(n7018) );
  or2_1 U7710 ( .ip1(n7018), .ip2(n7019), .op(n7022) );
  nand2_1 U7711 ( .ip1(n14629), .ip2(m1Inputs[105]), .op(n7020) );
  or2_1 U7712 ( .ip1(n7020), .ip2(n7019), .op(n7021) );
  nand2_1 U7713 ( .ip1(n7022), .ip2(n7021), .op(n7067) );
  nand3_1 U7714 ( .ip1(column[107]), .ip2(n15042), .ip3(n7067), .op(n7023) );
  nand2_1 U7715 ( .ip1(n7024), .ip2(n7023), .op(n7055) );
  inv_1 U7716 ( .ip(m1Inputs[107]), .op(n7474) );
  nor2_1 U7717 ( .ip1(n6503), .ip2(n7474), .op(n7064) );
  nor2_1 U7718 ( .ip1(n14170), .ip2(n14289), .op(n7063) );
  nand2_1 U7719 ( .ip1(n14976), .ip2(m1Inputs[100]), .op(n7062) );
  inv_1 U7720 ( .ip(n7026), .op(n7027) );
  nand2_1 U7721 ( .ip1(column[108]), .ip2(n13859), .op(n7025) );
  mux2_1 U7722 ( .ip1(n7027), .ip2(n7026), .s(n7025), .op(n7053) );
  fulladder U7723 ( .a(n7030), .b(n7029), .ci(n7028), .co(n14193), .s(n7127)
         );
  inv_1 U7724 ( .ip(n7031), .op(n14199) );
  nor2_1 U7725 ( .ip1(n12083), .ip2(n7331), .op(n14180) );
  nor2_1 U7726 ( .ip1(n14189), .ip2(n14368), .op(n14179) );
  nand2_1 U7727 ( .ip1(n14976), .ip2(m1Inputs[102]), .op(n14178) );
  nor2_1 U7728 ( .ip1(n14188), .ip2(n7518), .op(n14173) );
  nor2_1 U7729 ( .ip1(n6503), .ip2(n14170), .op(n14172) );
  nand2_1 U7730 ( .ip1(m1Inputs[111]), .ip2(n12981), .op(n14171) );
  fulladder U7731 ( .a(n7034), .b(n7033), .ci(n7032), .co(n14181), .s(n6988)
         );
  inv_1 U7732 ( .ip(n7035), .op(n14161) );
  nor2_1 U7733 ( .ip1(n14340), .ip2(n7518), .op(n14236) );
  nand3_1 U7734 ( .ip1(n14847), .ip2(m1Inputs[103]), .ip3(n14236), .op(n7038)
         );
  nand3_1 U7735 ( .ip1(n14816), .ip2(m1Inputs[102]), .ip3(n7036), .op(n7037)
         );
  nand2_1 U7736 ( .ip1(n7038), .ip2(n7037), .op(n14192) );
  nand2_1 U7737 ( .ip1(n14629), .ip2(m1Inputs[107]), .op(n7040) );
  nand2_1 U7738 ( .ip1(n13718), .ip2(m1Inputs[107]), .op(n14162) );
  nor2_1 U7739 ( .ip1(n14162), .ip2(n7039), .op(n14174) );
  or2_1 U7740 ( .ip1(n7040), .ip2(n14174), .op(n7043) );
  nand2_1 U7741 ( .ip1(n13718), .ip2(m1Inputs[106]), .op(n7041) );
  or2_1 U7742 ( .ip1(n7041), .ip2(n14174), .op(n7042) );
  nand2_1 U7743 ( .ip1(n7043), .ip2(n7042), .op(n14175) );
  inv_1 U7744 ( .ip(n14175), .op(n7045) );
  nand2_1 U7745 ( .ip1(column[109]), .ip2(n14768), .op(n7044) );
  mux2_1 U7746 ( .ip1(n7045), .ip2(n14175), .s(n7044), .op(n14191) );
  fulladder U7747 ( .a(n7048), .b(n7047), .ci(n7046), .co(n14190), .s(n6987)
         );
  inv_1 U7748 ( .ip(n7049), .op(n14160) );
  fulladder U7749 ( .a(n7052), .b(n7051), .ci(n7050), .co(n14159), .s(n6998)
         );
  fulladder U7750 ( .a(n7055), .b(n7054), .ci(n7053), .co(n14194), .s(n7056)
         );
  inv_1 U7751 ( .ip(n7056), .op(n7086) );
  nor2_1 U7752 ( .ip1(n14842), .ip2(n7326), .op(n7057) );
  xor2_1 U7753 ( .ip1(n7058), .ip2(n7057), .op(n7074) );
  fulladder U7754 ( .a(n7061), .b(n7060), .ci(n7059), .co(n7028), .s(n7073) );
  fulladder U7755 ( .a(n7064), .b(n7063), .ci(n7062), .co(n7054), .s(n7072) );
  inv_1 U7756 ( .ip(n7065), .op(n7085) );
  nand2_1 U7757 ( .ip1(column[107]), .ip2(n13498), .op(n7066) );
  xor2_1 U7758 ( .ip1(n7067), .ip2(n7066), .op(n7071) );
  nand2_1 U7759 ( .ip1(m1Inputs[109]), .ip2(\STAGE_1/weightReg [5]), .op(n7119) );
  nor2_1 U7760 ( .ip1(n7184), .ip2(n14853), .op(n7118) );
  inv_1 U7761 ( .ip(m1Inputs[111]), .op(n7176) );
  nor2_1 U7762 ( .ip1(n13801), .ip2(n7176), .op(n7115) );
  nand2_1 U7763 ( .ip1(m1Inputs[110]), .ip2(n13637), .op(n7114) );
  inv_1 U7764 ( .ip(n7068), .op(n14202) );
  fulladder U7765 ( .a(n7071), .b(n7070), .ci(n7069), .co(n7084), .s(n7133) );
  fulladder U7766 ( .a(n7074), .b(n7073), .ci(n7072), .co(n7065), .s(n7075) );
  inv_1 U7767 ( .ip(n7075), .op(n7132) );
  nor2_1 U7768 ( .ip1(n14842), .ip2(n7553), .op(n7077) );
  xor2_1 U7769 ( .ip1(n7077), .ip2(n7076), .op(n7140) );
  nor2_1 U7770 ( .ip1(n13594), .ip2(n7559), .op(n7121) );
  and2_1 U7771 ( .ip1(n7078), .ip2(n7121), .op(n7096) );
  nor2_1 U7772 ( .ip1(n14824), .ip2(n7559), .op(n7079) );
  or2_1 U7773 ( .ip1(m1Inputs[103]), .ip2(n7079), .op(n7081) );
  or2_1 U7774 ( .ip1(n14876), .ip2(n7079), .op(n7080) );
  nand2_1 U7775 ( .ip1(n7081), .ip2(n7080), .op(n7095) );
  nand2_1 U7776 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[100]), .op(
        n7097) );
  nor2_1 U7777 ( .ip1(n7095), .ip2(n7097), .op(n7082) );
  nor2_1 U7778 ( .ip1(n7096), .ip2(n7082), .op(n7139) );
  nor2_1 U7779 ( .ip1(n13854), .ip2(n7176), .op(n7145) );
  nand2_1 U7780 ( .ip1(n13614), .ip2(m1Inputs[110]), .op(n7253) );
  nand2_1 U7781 ( .ip1(m1Inputs[99]), .ip2(\STAGE_1/weightReg [14]), .op(n7144) );
  inv_1 U7782 ( .ip(n7083), .op(n7130) );
  fulladder U7783 ( .a(n7086), .b(n7085), .ci(n7084), .co(n14197), .s(n7087)
         );
  inv_1 U7784 ( .ip(n7087), .op(n7129) );
  fulladder U7785 ( .a(n7090), .b(n7089), .ci(n7088), .co(n7125), .s(n7192) );
  fulladder U7786 ( .a(n7093), .b(n7092), .ci(n7091), .co(n7088), .s(n7094) );
  inv_1 U7787 ( .ip(n7094), .op(n7164) );
  nor2_1 U7788 ( .ip1(n7096), .ip2(n7095), .op(n7098) );
  xor2_1 U7789 ( .ip1(n7098), .ip2(n7097), .op(n7206) );
  nand2_1 U7790 ( .ip1(m1Inputs[108]), .ip2(n13637), .op(n7211) );
  nor2_1 U7791 ( .ip1(n7564), .ip2(n14853), .op(n7210) );
  nor2_1 U7792 ( .ip1(n7331), .ip2(n12746), .op(n7100) );
  xor2_1 U7793 ( .ip1(n7100), .ip2(n7099), .op(n7204) );
  fulladder U7794 ( .a(n7103), .b(n7102), .ci(n7101), .co(n7091), .s(n7104) );
  inv_1 U7795 ( .ip(n7104), .op(n7203) );
  nor2_1 U7796 ( .ip1(n7518), .ip2(n14289), .op(n7169) );
  and3_1 U7797 ( .ip1(m1Inputs[106]), .ip2(n14835), .ip3(n7169), .op(n7109) );
  nor2_1 U7798 ( .ip1(n14187), .ip2(n14289), .op(n7105) );
  or2_1 U7799 ( .ip1(\STAGE_1/weightReg [7]), .ip2(n7105), .op(n7107) );
  or2_1 U7800 ( .ip1(m1Inputs[105]), .ip2(n7105), .op(n7106) );
  nand2_1 U7801 ( .ip1(n7107), .ip2(n7106), .op(n7108) );
  nor2_1 U7802 ( .ip1(n7109), .ip2(n7108), .op(n7188) );
  or2_1 U7803 ( .ip1(n7188), .ip2(n7109), .op(n7111) );
  nor2_1 U7804 ( .ip1(n7474), .ip2(n12746), .op(n7187) );
  or2_1 U7805 ( .ip1(n7187), .ip2(n7109), .op(n7110) );
  nand2_1 U7806 ( .ip1(n7111), .ip2(n7110), .op(n7202) );
  nor2_1 U7807 ( .ip1(n13570), .ip2(n7176), .op(n7208) );
  nand2_1 U7808 ( .ip1(n13614), .ip2(m1Inputs[109]), .op(n7289) );
  nand2_1 U7809 ( .ip1(m1Inputs[98]), .ip2(\STAGE_1/weightReg [14]), .op(n7207) );
  inv_1 U7810 ( .ip(n7112), .op(n7191) );
  fulladder U7811 ( .a(n7115), .b(n7114), .ci(n7113), .co(n7069), .s(n7116) );
  inv_1 U7812 ( .ip(n7116), .op(n7161) );
  fulladder U7813 ( .a(n7119), .b(n7118), .ci(n7117), .co(n7070), .s(n7120) );
  inv_1 U7814 ( .ip(n7120), .op(n7160) );
  nor2_1 U7815 ( .ip1(n14902), .ip2(n7326), .op(n7168) );
  or2_1 U7816 ( .ip1(m1Inputs[101]), .ip2(n7121), .op(n7123) );
  or2_1 U7817 ( .ip1(\STAGE_1/weightReg [11]), .ip2(n7121), .op(n7122) );
  nand2_1 U7818 ( .ip1(n7123), .ip2(n7122), .op(n7182) );
  nor3_1 U7819 ( .ip1(n7182), .ip2(n7184), .ip3(n14340), .op(n7124) );
  nor2_1 U7820 ( .ip1(n13594), .ip2(n7326), .op(n7258) );
  and3_1 U7821 ( .ip1(\STAGE_1/weightReg [11]), .ip2(m1Inputs[102]), .ip3(
        n7258), .op(n7183) );
  or2_1 U7822 ( .ip1(n7124), .ip2(n7183), .op(n7167) );
  nor2_1 U7823 ( .ip1(n12083), .ip2(n7492), .op(n7179) );
  nor2_1 U7824 ( .ip1(n13854), .ip2(n14189), .op(n7178) );
  fulladder U7825 ( .a(n7127), .b(n7126), .ci(n7125), .co(n14203), .s(n7687)
         );
  fulladder U7826 ( .a(n7130), .b(n7129), .ci(n7128), .co(n14201), .s(n7686)
         );
  fulladder U7827 ( .a(n7133), .b(n7132), .ci(n7131), .co(n7083), .s(n7134) );
  inv_1 U7828 ( .ip(n7134), .op(n7196) );
  fulladder U7829 ( .a(n7137), .b(n7136), .ci(n7135), .co(n7007), .s(n7200) );
  fulladder U7830 ( .a(n7140), .b(n7139), .ci(n7138), .co(n7131), .s(n7199) );
  fulladder U7831 ( .a(n7143), .b(n7142), .ci(n7141), .co(n7136), .s(n7222) );
  fulladder U7832 ( .a(n7145), .b(n7253), .ci(n7144), .co(n7138), .s(n7221) );
  nor3_1 U7833 ( .ip1(n7492), .ip2(n7209), .ip3(n14384), .op(n7250) );
  nor2_1 U7834 ( .ip1(n14169), .ip2(n14368), .op(n7146) );
  or2_1 U7835 ( .ip1(m1Inputs[103]), .ip2(n7146), .op(n7148) );
  or2_1 U7836 ( .ip1(n14838), .ip2(n7146), .op(n7147) );
  nand2_1 U7837 ( .ip1(n7148), .ip2(n7147), .op(n7249) );
  nand2_1 U7838 ( .ip1(m1Inputs[98]), .ip2(\STAGE_1/weightReg [13]), .op(n7251) );
  nor2_1 U7839 ( .ip1(n7249), .ip2(n7251), .op(n7149) );
  nor2_1 U7840 ( .ip1(n7250), .ip2(n7149), .op(n7240) );
  nand2_1 U7841 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[109]), .op(n7150) );
  nand2_1 U7842 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[109]), .op(n7213) );
  nor3_1 U7843 ( .ip1(n13709), .ip2(n14189), .ip3(n7213), .op(n7154) );
  or2_1 U7844 ( .ip1(n7150), .ip2(n7154), .op(n7153) );
  nand2_1 U7845 ( .ip1(n13707), .ip2(m1Inputs[110]), .op(n7151) );
  or2_1 U7846 ( .ip1(n7151), .ip2(n7154), .op(n7152) );
  nand2_1 U7847 ( .ip1(n7153), .ip2(n7152), .op(n7264) );
  or2_1 U7848 ( .ip1(n7264), .ip2(n7154), .op(n7157) );
  nand2_1 U7849 ( .ip1(column[103]), .ip2(n13498), .op(n7263) );
  inv_1 U7850 ( .ip(n7263), .op(n7155) );
  or2_1 U7851 ( .ip1(n7155), .ip2(n7154), .op(n7156) );
  nand2_1 U7852 ( .ip1(n7157), .ip2(n7156), .op(n7239) );
  nand2_1 U7853 ( .ip1(n15025), .ip2(m1Inputs[100]), .op(n7238) );
  inv_1 U7854 ( .ip(n7158), .op(n7195) );
  fulladder U7855 ( .a(n7161), .b(n7160), .ci(n7159), .co(n7190), .s(n7273) );
  fulladder U7856 ( .a(n7164), .b(n7163), .ci(n7162), .co(n7112), .s(n7165) );
  inv_1 U7857 ( .ip(n7165), .op(n7272) );
  fulladder U7858 ( .a(n7168), .b(n7167), .ci(n7166), .co(n7159), .s(n7277) );
  nand2_1 U7859 ( .ip1(m1Inputs[105]), .ip2(\STAGE_1/weightReg [4]), .op(n7318) );
  nor3_1 U7860 ( .ip1(n7474), .ip2(n14836), .ip3(n7318), .op(n7173) );
  or2_1 U7861 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n7169), .op(n7171) );
  or2_1 U7862 ( .ip1(m1Inputs[107]), .ip2(n7169), .op(n7170) );
  nand2_1 U7863 ( .ip1(n7171), .ip2(n7170), .op(n7172) );
  nor2_1 U7864 ( .ip1(n7173), .ip2(n7172), .op(n7229) );
  or2_1 U7865 ( .ip1(n7229), .ip2(n7173), .op(n7175) );
  nor2_1 U7866 ( .ip1(n7564), .ip2(n14842), .op(n7228) );
  or2_1 U7867 ( .ip1(n7228), .ip2(n7173), .op(n7174) );
  nand2_1 U7868 ( .ip1(n7175), .ip2(n7174), .op(n7235) );
  nand2_1 U7869 ( .ip1(n13614), .ip2(m1Inputs[108]), .op(n7398) );
  nor2_1 U7870 ( .ip1(n10476), .ip2(n7176), .op(n7224) );
  nand2_1 U7871 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[102]), .op(n7223) );
  fulladder U7872 ( .a(n7179), .b(n7178), .ci(n7177), .co(n7166), .s(n7180) );
  inv_1 U7873 ( .ip(n7180), .op(n7233) );
  inv_1 U7874 ( .ip(n7181), .op(n7276) );
  nor2_1 U7875 ( .ip1(n7183), .ip2(n7182), .op(n7186) );
  nor2_1 U7876 ( .ip1(n7184), .ip2(n14340), .op(n7185) );
  xor2_1 U7877 ( .ip1(n7186), .ip2(n7185), .op(n7232) );
  xor2_1 U7878 ( .ip1(n7188), .ip2(n7187), .op(n7231) );
  nor2_1 U7879 ( .ip1(n14187), .ip2(n4624), .op(n7227) );
  nand2_1 U7880 ( .ip1(m1Inputs[96]), .ip2(\STAGE_1/weightReg [15]), .op(n7226) );
  inv_1 U7881 ( .ip(n7189), .op(n14137) );
  fulladder U7882 ( .a(n7192), .b(n7191), .ci(n7190), .co(n7128), .s(n7193) );
  inv_1 U7883 ( .ip(n7193), .op(n7267) );
  fulladder U7884 ( .a(n7196), .b(n7195), .ci(n7194), .co(n7685), .s(n7197) );
  inv_1 U7885 ( .ip(n7197), .op(n7266) );
  fulladder U7886 ( .a(n7200), .b(n7199), .ci(n7198), .co(n7158), .s(n7270) );
  fulladder U7887 ( .a(n7203), .b(n7202), .ci(n7201), .co(n7162), .s(n7281) );
  fulladder U7888 ( .a(n7206), .b(n7205), .ci(n7204), .co(n7163), .s(n7280) );
  fulladder U7889 ( .a(n7208), .b(n7289), .ci(n7207), .co(n7201), .s(n7284) );
  fulladder U7890 ( .a(n7211), .b(n7210), .ci(n7209), .co(n7205), .s(n7283) );
  nand2_1 U7891 ( .ip1(n4672), .ip2(m1Inputs[108]), .op(n7212) );
  nand2_1 U7892 ( .ip1(n13707), .ip2(m1Inputs[108]), .op(n7333) );
  nor3_1 U7893 ( .ip1(n13709), .ip2(n14170), .ip3(n7333), .op(n7216) );
  or2_1 U7894 ( .ip1(n7212), .ip2(n7216), .op(n7215) );
  or2_1 U7895 ( .ip1(n7213), .ip2(n7216), .op(n7214) );
  nand2_1 U7896 ( .ip1(n7215), .ip2(n7214), .op(n7325) );
  or2_1 U7897 ( .ip1(n7325), .ip2(n7216), .op(n7219) );
  nand2_1 U7898 ( .ip1(column[102]), .ip2(n13498), .op(n7324) );
  inv_1 U7899 ( .ip(n7324), .op(n7217) );
  or2_1 U7900 ( .ip1(n7217), .ip2(n7216), .op(n7218) );
  nand2_1 U7901 ( .ip1(n7219), .ip2(n7218), .op(n7309) );
  nand2_1 U7902 ( .ip1(m1Inputs[99]), .ip2(\STAGE_1/weightReg [12]), .op(n7308) );
  nand2_1 U7903 ( .ip1(n13718), .ip2(m1Inputs[100]), .op(n7307) );
  fulladder U7904 ( .a(n7222), .b(n7221), .ci(n7220), .co(n7198), .s(n7345) );
  fulladder U7905 ( .a(n7398), .b(n7224), .ci(n7223), .co(n7234), .s(n7225) );
  inv_1 U7906 ( .ip(n7225), .op(n7358) );
  fulladder U7907 ( .a(n7227), .b(n7258), .ci(n7226), .co(n7230), .s(n7357) );
  xor2_1 U7908 ( .ip1(n7229), .ip2(n7228), .op(n7356) );
  fulladder U7909 ( .a(n7232), .b(n7231), .ci(n7230), .co(n7275), .s(n7353) );
  fulladder U7910 ( .a(n7235), .b(n7234), .ci(n7233), .co(n7181), .s(n7236) );
  inv_1 U7911 ( .ip(n7236), .op(n7352) );
  inv_1 U7912 ( .ip(n7237), .op(n7344) );
  fulladder U7913 ( .a(n7240), .b(n7239), .ci(n7238), .co(n7220), .s(n7351) );
  nor3_1 U7914 ( .ip1(n14187), .ip2(n4624), .ip3(n7318), .op(n7378) );
  nor2_1 U7915 ( .ip1(n7518), .ip2(n12746), .op(n7241) );
  or2_1 U7916 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n7241), .op(n7243) );
  or2_1 U7917 ( .ip1(m1Inputs[106]), .ip2(n7241), .op(n7242) );
  nand2_1 U7918 ( .ip1(n7243), .ip2(n7242), .op(n7377) );
  nand2_1 U7919 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[102]), .op(n7379) );
  nor2_1 U7920 ( .ip1(n7377), .ip2(n7379), .op(n7244) );
  nor2_1 U7921 ( .ip1(n7378), .ip2(n7244), .op(n7303) );
  nor3_1 U7922 ( .ip1(n14169), .ip2(n14368), .ip3(n7311), .op(n7286) );
  nor2_1 U7923 ( .ip1(n7492), .ip2(n14384), .op(n7245) );
  or2_1 U7924 ( .ip1(n13749), .ip2(n7245), .op(n7247) );
  or2_1 U7925 ( .ip1(m1Inputs[104]), .ip2(n7245), .op(n7246) );
  nand2_1 U7926 ( .ip1(n7247), .ip2(n7246), .op(n7285) );
  nand2_1 U7927 ( .ip1(m1Inputs[97]), .ip2(\STAGE_1/weightReg [13]), .op(n7287) );
  nor2_1 U7928 ( .ip1(n7285), .ip2(n7287), .op(n7248) );
  nor2_1 U7929 ( .ip1(n7286), .ip2(n7248), .op(n7302) );
  nor2_1 U7930 ( .ip1(n7250), .ip2(n7249), .op(n7252) );
  xor2_1 U7931 ( .ip1(n7252), .ip2(n7251), .op(n7301) );
  nand2_1 U7932 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[107]), .op(n7476) );
  nor2_1 U7933 ( .ip1(n7476), .ip2(n7253), .op(n7382) );
  nor2_1 U7934 ( .ip1(n13801), .ip2(n7474), .op(n7254) );
  or2_1 U7935 ( .ip1(m1Inputs[110]), .ip2(n7254), .op(n7256) );
  or2_1 U7936 ( .ip1(n13803), .ip2(n7254), .op(n7255) );
  nand2_1 U7937 ( .ip1(n7256), .ip2(n7255), .op(n7381) );
  nand2_1 U7938 ( .ip1(m1Inputs[96]), .ip2(n14816), .op(n7383) );
  nor2_1 U7939 ( .ip1(n7381), .ip2(n7383), .op(n7257) );
  nor2_1 U7940 ( .ip1(n7382), .ip2(n7257), .op(n7306) );
  nor2_1 U7941 ( .ip1(n13766), .ip2(n7553), .op(n7327) );
  and2_1 U7942 ( .ip1(n7327), .ip2(n7258), .op(n7298) );
  nor2_1 U7943 ( .ip1(n13766), .ip2(n7326), .op(n7259) );
  or2_1 U7944 ( .ip1(m1Inputs[100]), .ip2(n7259), .op(n7261) );
  or2_1 U7945 ( .ip1(n14876), .ip2(n7259), .op(n7260) );
  nand2_1 U7946 ( .ip1(n7261), .ip2(n7260), .op(n7297) );
  nand2_1 U7947 ( .ip1(m1Inputs[98]), .ip2(\STAGE_1/weightReg [12]), .op(n7299) );
  nor2_1 U7948 ( .ip1(n7297), .ip2(n7299), .op(n7262) );
  nor2_1 U7949 ( .ip1(n7298), .ip2(n7262), .op(n7305) );
  xor2_1 U7950 ( .ip1(n7264), .ip2(n7263), .op(n7304) );
  fulladder U7951 ( .a(n7267), .b(n7266), .ci(n7265), .co(n14136), .s(n14141)
         );
  fulladder U7952 ( .a(n7270), .b(n7269), .ci(n7268), .co(n7265), .s(n7342) );
  fulladder U7953 ( .a(n7273), .b(n7272), .ci(n7271), .co(n7194), .s(n7274) );
  inv_1 U7954 ( .ip(n7274), .op(n7341) );
  fulladder U7955 ( .a(n7277), .b(n7276), .ci(n7275), .co(n7271), .s(n7278) );
  inv_1 U7956 ( .ip(n7278), .op(n7348) );
  fulladder U7957 ( .a(n7281), .b(n7280), .ci(n7279), .co(n7269), .s(n7347) );
  fulladder U7958 ( .a(n7284), .b(n7283), .ci(n7282), .co(n7279), .s(n7416) );
  nor2_1 U7959 ( .ip1(n7286), .ip2(n7285), .op(n7288) );
  xor2_1 U7960 ( .ip1(n7288), .ip2(n7287), .op(n7428) );
  nand2_1 U7961 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[106]), .op(n7529) );
  nor2_1 U7962 ( .ip1(n7529), .ip2(n7289), .op(n7294) );
  nor2_1 U7963 ( .ip1(n13487), .ip2(n14187), .op(n7290) );
  or2_1 U7964 ( .ip1(m1Inputs[109]), .ip2(n7290), .op(n7292) );
  or2_1 U7965 ( .ip1(n13803), .ip2(n7290), .op(n7291) );
  nand2_1 U7966 ( .ip1(n7292), .ip2(n7291), .op(n7293) );
  nor2_1 U7967 ( .ip1(n7294), .ip2(n7293), .op(n7435) );
  or2_1 U7968 ( .ip1(n7435), .ip2(n7294), .op(n7296) );
  nor2_1 U7969 ( .ip1(n7532), .ip2(n14340), .op(n7434) );
  or2_1 U7970 ( .ip1(n7434), .ip2(n7294), .op(n7295) );
  nand2_1 U7971 ( .ip1(n7296), .ip2(n7295), .op(n7427) );
  nor2_1 U7972 ( .ip1(n7298), .ip2(n7297), .op(n7300) );
  xor2_1 U7973 ( .ip1(n7300), .ip2(n7299), .op(n7426) );
  fulladder U7974 ( .a(n7303), .b(n7302), .ci(n7301), .co(n7350), .s(n7423) );
  fulladder U7975 ( .a(n7306), .b(n7305), .ci(n7304), .co(n7349), .s(n7422) );
  fulladder U7976 ( .a(n7309), .b(n7308), .ci(n7307), .co(n7282), .s(n7420) );
  nand2_1 U7977 ( .ip1(m1Inputs[102]), .ip2(\STAGE_1/weightReg [7]), .op(n7310) );
  nand2_1 U7978 ( .ip1(m1Inputs[102]), .ip2(n12981), .op(n7369) );
  nor3_1 U7979 ( .ip1(n7492), .ip2(n14368), .ip3(n7369), .op(n7314) );
  or2_1 U7980 ( .ip1(n7310), .ip2(n7314), .op(n7313) );
  or2_1 U7981 ( .ip1(n7311), .ip2(n7314), .op(n7312) );
  nand2_1 U7982 ( .ip1(n7313), .ip2(n7312), .op(n7439) );
  or2_1 U7983 ( .ip1(n7439), .ip2(n7314), .op(n7316) );
  nor2_1 U7984 ( .ip1(n7486), .ip2(n14824), .op(n7438) );
  or2_1 U7985 ( .ip1(n7438), .ip2(n7314), .op(n7315) );
  nand2_1 U7986 ( .ip1(n7316), .ip2(n7315), .op(n7390) );
  nand2_1 U7987 ( .ip1(m1Inputs[104]), .ip2(n14369), .op(n7317) );
  nand2_1 U7988 ( .ip1(m1Inputs[104]), .ip2(n11974), .op(n7392) );
  nor3_1 U7989 ( .ip1(n7518), .ip2(n4624), .ip3(n7392), .op(n7321) );
  or2_1 U7990 ( .ip1(n7317), .ip2(n7321), .op(n7320) );
  or2_1 U7991 ( .ip1(n7318), .ip2(n7321), .op(n7319) );
  nand2_1 U7992 ( .ip1(n7320), .ip2(n7319), .op(n7437) );
  or2_1 U7993 ( .ip1(n7437), .ip2(n7321), .op(n7323) );
  nor2_1 U7994 ( .ip1(n7564), .ip2(n14902), .op(n7436) );
  or2_1 U7995 ( .ip1(n7436), .ip2(n7321), .op(n7322) );
  nand2_1 U7996 ( .ip1(n7323), .ip2(n7322), .op(n7389) );
  xor2_1 U7997 ( .ip1(n7325), .ip2(n7324), .op(n7388) );
  nand2_1 U7998 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[100]), .op(n7538) );
  nor3_1 U7999 ( .ip1(n12083), .ip2(n7326), .ip3(n7538), .op(n7404) );
  or2_1 U8000 ( .ip1(m1Inputs[101]), .ip2(n7327), .op(n7329) );
  or2_1 U8001 ( .ip1(n14838), .ip2(n7327), .op(n7328) );
  nand2_1 U8002 ( .ip1(n7329), .ip2(n7328), .op(n7403) );
  nand2_1 U8003 ( .ip1(m1Inputs[99]), .ip2(\STAGE_1/weightReg [10]), .op(n7405) );
  nor2_1 U8004 ( .ip1(n7403), .ip2(n7405), .op(n7330) );
  nor2_1 U8005 ( .ip1(n7404), .ip2(n7330), .op(n7387) );
  nand2_1 U8006 ( .ip1(n4619), .ip2(m1Inputs[107]), .op(n7332) );
  nand2_1 U8007 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[107]), .op(n7361) );
  nor3_1 U8008 ( .ip1(n13709), .ip2(n7331), .ip3(n7361), .op(n7336) );
  or2_1 U8009 ( .ip1(n7332), .ip2(n7336), .op(n7335) );
  or2_1 U8010 ( .ip1(n7333), .ip2(n7336), .op(n7334) );
  nand2_1 U8011 ( .ip1(n7335), .ip2(n7334), .op(n7376) );
  or2_1 U8012 ( .ip1(n7376), .ip2(n7336), .op(n7339) );
  nand2_1 U8013 ( .ip1(column[101]), .ip2(n13859), .op(n7375) );
  inv_1 U8014 ( .ip(n7375), .op(n7337) );
  or2_1 U8015 ( .ip1(n7337), .ip2(n7336), .op(n7338) );
  nand2_1 U8016 ( .ip1(n7339), .ip2(n7338), .op(n7386) );
  nand2_1 U8017 ( .ip1(m1Inputs[99]), .ip2(\STAGE_1/weightReg [11]), .op(n7385) );
  fulladder U8018 ( .a(n7342), .b(n7341), .ci(n7340), .co(n14140), .s(n14145)
         );
  fulladder U8019 ( .a(n7345), .b(n7344), .ci(n7343), .co(n7268), .s(n7409) );
  fulladder U8020 ( .a(n7348), .b(n7347), .ci(n7346), .co(n7340), .s(n7408) );
  fulladder U8021 ( .a(n7351), .b(n7350), .ci(n7349), .co(n7343), .s(n7412) );
  fulladder U8022 ( .a(n7354), .b(n7353), .ci(n7352), .co(n7237), .s(n7355) );
  inv_1 U8023 ( .ip(n7355), .op(n7411) );
  fulladder U8024 ( .a(n7358), .b(n7357), .ci(n7356), .co(n7354), .s(n7359) );
  inv_1 U8025 ( .ip(n7359), .op(n7447) );
  nand2_1 U8026 ( .ip1(n4619), .ip2(m1Inputs[106]), .op(n7360) );
  nand2_1 U8027 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[106]), .op(n7466) );
  nor3_1 U8028 ( .ip1(n13709), .ip2(n7474), .ip3(n7466), .op(n7364) );
  or2_1 U8029 ( .ip1(n7360), .ip2(n7364), .op(n7363) );
  or2_1 U8030 ( .ip1(n7361), .ip2(n7364), .op(n7362) );
  nand2_1 U8031 ( .ip1(n7363), .ip2(n7362), .op(n7491) );
  or2_1 U8032 ( .ip1(n7491), .ip2(n7364), .op(n7367) );
  nand2_1 U8033 ( .ip1(column[100]), .ip2(n13498), .op(n7490) );
  inv_1 U8034 ( .ip(n7490), .op(n7365) );
  or2_1 U8035 ( .ip1(n7365), .ip2(n7364), .op(n7366) );
  nand2_1 U8036 ( .ip1(n7367), .ip2(n7366), .op(n7464) );
  nand2_1 U8037 ( .ip1(n4627), .ip2(m1Inputs[101]), .op(n7368) );
  nand2_1 U8038 ( .ip1(n13749), .ip2(m1Inputs[101]), .op(n7483) );
  nor3_1 U8039 ( .ip1(n7559), .ip2(n14384), .ip3(n7483), .op(n7372) );
  or2_1 U8040 ( .ip1(n7368), .ip2(n7372), .op(n7371) );
  or2_1 U8041 ( .ip1(n7369), .ip2(n7372), .op(n7370) );
  nand2_1 U8042 ( .ip1(n7371), .ip2(n7370), .op(n7503) );
  or2_1 U8043 ( .ip1(n7503), .ip2(n7372), .op(n7374) );
  nor2_1 U8044 ( .ip1(n7486), .ip2(n13390), .op(n7502) );
  or2_1 U8045 ( .ip1(n7502), .ip2(n7372), .op(n7373) );
  nand2_1 U8046 ( .ip1(n7374), .ip2(n7373), .op(n7463) );
  xor2_1 U8047 ( .ip1(n7376), .ip2(n7375), .op(n7462) );
  nor2_1 U8048 ( .ip1(n7378), .ip2(n7377), .op(n7380) );
  xor2_1 U8049 ( .ip1(n7380), .ip2(n7379), .op(n7431) );
  nor2_1 U8050 ( .ip1(n7382), .ip2(n7381), .op(n7384) );
  xor2_1 U8051 ( .ip1(n7384), .ip2(n7383), .op(n7430) );
  fulladder U8052 ( .a(n7387), .b(n7386), .ci(n7385), .co(n7418), .s(n7454) );
  fulladder U8053 ( .a(n7390), .b(n7389), .ci(n7388), .co(n7419), .s(n7453) );
  nand2_1 U8054 ( .ip1(m1Inputs[103]), .ip2(n14369), .op(n7391) );
  nand2_1 U8055 ( .ip1(m1Inputs[103]), .ip2(n13637), .op(n7494) );
  nor3_1 U8056 ( .ip1(n14169), .ip2(n12746), .ip3(n7494), .op(n7395) );
  or2_1 U8057 ( .ip1(n7391), .ip2(n7395), .op(n7394) );
  or2_1 U8058 ( .ip1(n7392), .ip2(n7395), .op(n7393) );
  nand2_1 U8059 ( .ip1(n7394), .ip2(n7393), .op(n7501) );
  or2_1 U8060 ( .ip1(n7501), .ip2(n7395), .op(n7397) );
  nor2_1 U8061 ( .ip1(n7564), .ip2(n13579), .op(n7500) );
  or2_1 U8062 ( .ip1(n7500), .ip2(n7395), .op(n7396) );
  nand2_1 U8063 ( .ip1(n7397), .ip2(n7396), .op(n7457) );
  nor3_1 U8064 ( .ip1(n10476), .ip2(n7518), .ip3(n7398), .op(n7540) );
  nor2_1 U8065 ( .ip1(n13801), .ip2(n7518), .op(n7399) );
  or2_1 U8066 ( .ip1(m1Inputs[108]), .ip2(n7399), .op(n7401) );
  or2_1 U8067 ( .ip1(n13803), .ip2(n7399), .op(n7400) );
  nand2_1 U8068 ( .ip1(n7401), .ip2(n7400), .op(n7539) );
  nand2_1 U8069 ( .ip1(m1Inputs[96]), .ip2(\STAGE_1/weightReg [12]), .op(n7541) );
  nor2_1 U8070 ( .ip1(n7539), .ip2(n7541), .op(n7402) );
  nor2_1 U8071 ( .ip1(n7540), .ip2(n7402), .op(n7456) );
  nor2_1 U8072 ( .ip1(n7404), .ip2(n7403), .op(n7406) );
  xor2_1 U8073 ( .ip1(n7406), .ip2(n7405), .op(n7455) );
  fulladder U8074 ( .a(n7409), .b(n7408), .ci(n7407), .co(n14144), .s(n14149)
         );
  fulladder U8075 ( .a(n7412), .b(n7411), .ci(n7410), .co(n7407), .s(n7413) );
  inv_1 U8076 ( .ip(n7413), .op(n7443) );
  fulladder U8077 ( .a(n7416), .b(n7415), .ci(n7414), .co(n7346), .s(n7417) );
  inv_1 U8078 ( .ip(n7417), .op(n7442) );
  fulladder U8079 ( .a(n7420), .b(n7419), .ci(n7418), .co(n7414), .s(n7421) );
  inv_1 U8080 ( .ip(n7421), .op(n7450) );
  fulladder U8081 ( .a(n7424), .b(n7423), .ci(n7422), .co(n7415), .s(n7425) );
  inv_1 U8082 ( .ip(n7425), .op(n7449) );
  fulladder U8083 ( .a(n7428), .b(n7427), .ci(n7426), .co(n7424), .s(n7429) );
  inv_1 U8084 ( .ip(n7429), .op(n7512) );
  fulladder U8085 ( .a(n7432), .b(n7431), .ci(n7430), .co(n7446), .s(n7433) );
  inv_1 U8086 ( .ip(n7433), .op(n7511) );
  xor2_1 U8087 ( .ip1(n7435), .ip2(n7434), .op(n7460) );
  xor2_1 U8088 ( .ip1(n7437), .ip2(n7436), .op(n7459) );
  xor2_1 U8089 ( .ip1(n7439), .ip2(n7438), .op(n7458) );
  inv_1 U8090 ( .ip(n7440), .op(n14148) );
  fulladder U8091 ( .a(n7443), .b(n7442), .ci(n7441), .co(n7440), .s(n7444) );
  inv_1 U8092 ( .ip(n7444), .op(n14153) );
  fulladder U8093 ( .a(n7447), .b(n7446), .ci(n7445), .co(n7410), .s(n7506) );
  fulladder U8094 ( .a(n7450), .b(n7449), .ci(n7448), .co(n7441), .s(n7451) );
  inv_1 U8095 ( .ip(n7451), .op(n7505) );
  fulladder U8096 ( .a(n7454), .b(n7453), .ci(n7452), .co(n7445), .s(n7509) );
  fulladder U8097 ( .a(n7457), .b(n7456), .ci(n7455), .co(n7452), .s(n7573) );
  fulladder U8098 ( .a(n7460), .b(n7459), .ci(n7458), .co(n7510), .s(n7461) );
  inv_1 U8099 ( .ip(n7461), .op(n7572) );
  fulladder U8100 ( .a(n7464), .b(n7463), .ci(n7462), .co(n7432), .s(n7571) );
  nand2_1 U8101 ( .ip1(n4619), .ip2(m1Inputs[105]), .op(n7465) );
  nand2_1 U8102 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[105]), .op(n7520) );
  nor3_1 U8103 ( .ip1(n13709), .ip2(n14187), .ip3(n7520), .op(n7469) );
  or2_1 U8104 ( .ip1(n7465), .ip2(n7469), .op(n7468) );
  or2_1 U8105 ( .ip1(n7466), .ip2(n7469), .op(n7467) );
  nand2_1 U8106 ( .ip1(n7468), .ip2(n7467), .op(n7569) );
  or2_1 U8107 ( .ip1(n7569), .ip2(n7469), .op(n7472) );
  nand2_1 U8108 ( .ip1(column[99]), .ip2(n13498), .op(n7568) );
  inv_1 U8109 ( .ip(n7568), .op(n7470) );
  or2_1 U8110 ( .ip1(n7470), .ip2(n7469), .op(n7471) );
  nand2_1 U8111 ( .ip1(n7472), .ip2(n7471), .op(n7537) );
  nand2_1 U8112 ( .ip1(m1Inputs[99]), .ip2(n14994), .op(n7536) );
  nand2_1 U8113 ( .ip1(n13614), .ip2(m1Inputs[104]), .op(n7475) );
  nor3_1 U8114 ( .ip1(n13801), .ip2(n7474), .ip3(n7473), .op(n7479) );
  or2_1 U8115 ( .ip1(n7475), .ip2(n7479), .op(n7478) );
  or2_1 U8116 ( .ip1(n7476), .ip2(n7479), .op(n7477) );
  nand2_1 U8117 ( .ip1(n7478), .ip2(n7477), .op(n7551) );
  or2_1 U8118 ( .ip1(n7551), .ip2(n7479), .op(n7481) );
  nor2_1 U8119 ( .ip1(n7532), .ip2(n14824), .op(n7550) );
  or2_1 U8120 ( .ip1(n7550), .ip2(n7479), .op(n7480) );
  nand2_1 U8121 ( .ip1(n7481), .ip2(n7480), .op(n7545) );
  nand2_1 U8122 ( .ip1(m1Inputs[100]), .ip2(\STAGE_1/weightReg [7]), .op(n7482) );
  nor2_1 U8123 ( .ip1(n7553), .ip2(n14289), .op(n7554) );
  and3_1 U8124 ( .ip1(n4627), .ip2(m1Inputs[101]), .ip3(n7554), .op(n7487) );
  or2_1 U8125 ( .ip1(n7482), .ip2(n7487), .op(n7485) );
  or2_1 U8126 ( .ip1(n7483), .ip2(n7487), .op(n7484) );
  nand2_1 U8127 ( .ip1(n7485), .ip2(n7484), .op(n7547) );
  or2_1 U8128 ( .ip1(n7547), .ip2(n7487), .op(n7489) );
  nor2_1 U8129 ( .ip1(n7486), .ip2(n12083), .op(n7546) );
  or2_1 U8130 ( .ip1(n7546), .ip2(n7487), .op(n7488) );
  nand2_1 U8131 ( .ip1(n7489), .ip2(n7488), .op(n7544) );
  xor2_1 U8132 ( .ip1(n7491), .ip2(n7490), .op(n7543) );
  nand2_1 U8133 ( .ip1(m1Inputs[102]), .ip2(n14369), .op(n7493) );
  nand2_1 U8134 ( .ip1(m1Inputs[102]), .ip2(n11974), .op(n7561) );
  nor3_1 U8135 ( .ip1(n7492), .ip2(n4624), .ip3(n7561), .op(n7497) );
  or2_1 U8136 ( .ip1(n7493), .ip2(n7497), .op(n7496) );
  or2_1 U8137 ( .ip1(n7494), .ip2(n7497), .op(n7495) );
  nand2_1 U8138 ( .ip1(n7496), .ip2(n7495), .op(n7549) );
  or2_1 U8139 ( .ip1(n7549), .ip2(n7497), .op(n7499) );
  nor2_1 U8140 ( .ip1(n7564), .ip2(n13390), .op(n7548) );
  or2_1 U8141 ( .ip1(n7548), .ip2(n7497), .op(n7498) );
  nand2_1 U8142 ( .ip1(n7499), .ip2(n7498), .op(n7579) );
  xnor2_1 U8143 ( .ip1(n7501), .ip2(n7500), .op(n7578) );
  xnor2_1 U8144 ( .ip1(n7503), .ip2(n7502), .op(n7577) );
  fulladder U8145 ( .a(n7506), .b(n7505), .ci(n7504), .co(n14152), .s(n14157)
         );
  fulladder U8146 ( .a(n7509), .b(n7508), .ci(n7507), .co(n7504), .s(n7683) );
  fulladder U8147 ( .a(n7512), .b(n7511), .ci(n7510), .co(n7448), .s(n7513) );
  inv_1 U8148 ( .ip(n7513), .op(n7682) );
  fulladder U8149 ( .a(n7516), .b(n7515), .ci(n7514), .co(n7507), .s(n7576) );
  nand2_1 U8150 ( .ip1(n4619), .ip2(m1Inputs[104]), .op(n7519) );
  nor3_1 U8151 ( .ip1(n13709), .ip2(n7518), .ip3(n7517), .op(n7523) );
  or2_1 U8152 ( .ip1(n7519), .ip2(n7523), .op(n7522) );
  or2_1 U8153 ( .ip1(n7520), .ip2(n7523), .op(n7521) );
  nand2_1 U8154 ( .ip1(n7522), .ip2(n7521), .op(n7608) );
  or2_1 U8155 ( .ip1(n7608), .ip2(n7523), .op(n7526) );
  nand2_1 U8156 ( .ip1(column[98]), .ip2(n13498), .op(n7607) );
  inv_1 U8157 ( .ip(n7607), .op(n7524) );
  or2_1 U8158 ( .ip1(n7524), .ip2(n7523), .op(n7525) );
  nand2_1 U8159 ( .ip1(n7526), .ip2(n7525), .op(n7585) );
  nand2_1 U8160 ( .ip1(n13614), .ip2(m1Inputs[103]), .op(n7528) );
  nor3_1 U8161 ( .ip1(n13082), .ip2(n14187), .ip3(n7527), .op(n7533) );
  or2_1 U8162 ( .ip1(n7528), .ip2(n7533), .op(n7531) );
  or2_1 U8163 ( .ip1(n7529), .ip2(n7533), .op(n7530) );
  nand2_1 U8164 ( .ip1(n7531), .ip2(n7530), .op(n7628) );
  or2_1 U8165 ( .ip1(n7628), .ip2(n7533), .op(n7535) );
  nor2_1 U8166 ( .ip1(n7532), .ip2(n13594), .op(n7627) );
  or2_1 U8167 ( .ip1(n7627), .ip2(n7533), .op(n7534) );
  nand2_1 U8168 ( .ip1(n7535), .ip2(n7534), .op(n7584) );
  nand2_1 U8169 ( .ip1(m1Inputs[99]), .ip2(n14975), .op(n7583) );
  fulladder U8170 ( .a(n7538), .b(n7537), .ci(n7536), .co(n7516), .s(n7581) );
  nor2_1 U8171 ( .ip1(n7540), .ip2(n7539), .op(n7542) );
  xor2_1 U8172 ( .ip1(n7542), .ip2(n7541), .op(n7580) );
  fulladder U8173 ( .a(n7545), .b(n7544), .ci(n7543), .co(n7515), .s(n7616) );
  xor2_1 U8174 ( .ip1(n7547), .ip2(n7546), .op(n7625) );
  xor2_1 U8175 ( .ip1(n7549), .ip2(n7548), .op(n7624) );
  xor2_1 U8176 ( .ip1(n7551), .ip2(n7550), .op(n7623) );
  inv_1 U8177 ( .ip(n7552), .op(n7615) );
  nor3_1 U8178 ( .ip1(n7553), .ip2(n14368), .ip3(n7633), .op(n7587) );
  or2_1 U8179 ( .ip1(n14835), .ip2(n7554), .op(n7556) );
  or2_1 U8180 ( .ip1(m1Inputs[99]), .ip2(n7554), .op(n7555) );
  nand2_1 U8181 ( .ip1(n7556), .ip2(n7555), .op(n7586) );
  nand2_1 U8182 ( .ip1(m1Inputs[98]), .ip2(n14975), .op(n7588) );
  nor2_1 U8183 ( .ip1(n7586), .ip2(n7588), .op(n7557) );
  nor2_1 U8184 ( .ip1(n7587), .ip2(n7557), .op(n7622) );
  nand2_1 U8185 ( .ip1(n14369), .ip2(m1Inputs[101]), .op(n7560) );
  nor3_1 U8186 ( .ip1(n7559), .ip2(n4624), .ip3(n7558), .op(n7565) );
  or2_1 U8187 ( .ip1(n7560), .ip2(n7565), .op(n7563) );
  or2_1 U8188 ( .ip1(n7561), .ip2(n7565), .op(n7562) );
  nand2_1 U8189 ( .ip1(n7563), .ip2(n7562), .op(n7595) );
  or2_1 U8190 ( .ip1(n7595), .ip2(n7565), .op(n7567) );
  nor2_1 U8191 ( .ip1(n7564), .ip2(n13766), .op(n7594) );
  or2_1 U8192 ( .ip1(n7594), .ip2(n7565), .op(n7566) );
  nand2_1 U8193 ( .ip1(n7567), .ip2(n7566), .op(n7621) );
  xor2_1 U8194 ( .ip1(n7569), .ip2(n7568), .op(n7620) );
  inv_1 U8195 ( .ip(n7570), .op(n7690) );
  fulladder U8196 ( .a(n7573), .b(n7572), .ci(n7571), .co(n7508), .s(n7612) );
  fulladder U8197 ( .a(n7576), .b(n7575), .ci(n7574), .co(n7681), .s(n7611) );
  fulladder U8198 ( .a(n7579), .b(n7578), .ci(n7577), .co(n7514), .s(n7619) );
  fulladder U8199 ( .a(n7582), .b(n7581), .ci(n7580), .co(n7575), .s(n7618) );
  fulladder U8200 ( .a(n7585), .b(n7584), .ci(n7583), .co(n7582), .s(n7642) );
  nor2_1 U8201 ( .ip1(n7587), .ip2(n7586), .op(n7589) );
  xor2_1 U8202 ( .ip1(n7589), .ip2(n7588), .op(n7651) );
  nor2_1 U8203 ( .ip1(n7591), .ip2(n7590), .op(n7592) );
  nor2_1 U8204 ( .ip1(n7593), .ip2(n7592), .op(n7650) );
  xnor2_1 U8205 ( .ip1(n7595), .ip2(n7594), .op(n7649) );
  or2_1 U8206 ( .ip1(n7596), .ip2(n7597), .op(n7600) );
  or2_1 U8207 ( .ip1(n7598), .ip2(n7597), .op(n7599) );
  nand2_1 U8208 ( .ip1(n7600), .ip2(n7599), .op(n7648) );
  or2_1 U8209 ( .ip1(n7601), .ip2(n7603), .op(n7606) );
  inv_1 U8210 ( .ip(n7602), .op(n7604) );
  or2_1 U8211 ( .ip1(n7604), .ip2(n7603), .op(n7605) );
  nand2_1 U8212 ( .ip1(n7606), .ip2(n7605), .op(n7647) );
  xor2_1 U8213 ( .ip1(n7608), .ip2(n7607), .op(n7646) );
  inv_1 U8214 ( .ip(n7609), .op(n7689) );
  fulladder U8215 ( .a(n7612), .b(n7611), .ci(n7610), .co(n7609), .s(n7613) );
  inv_1 U8216 ( .ip(n7613), .op(n7693) );
  fulladder U8217 ( .a(n7616), .b(n7615), .ci(n7614), .co(n7574), .s(n7638) );
  fulladder U8218 ( .a(n7619), .b(n7618), .ci(n7617), .co(n7610), .s(n7637) );
  fulladder U8219 ( .a(n7622), .b(n7621), .ci(n7620), .co(n7614), .s(n7645) );
  fulladder U8220 ( .a(n7625), .b(n7624), .ci(n7623), .co(n7552), .s(n7626) );
  inv_1 U8221 ( .ip(n7626), .op(n7644) );
  xnor2_1 U8222 ( .ip1(n7628), .ip2(n7627), .op(n7662) );
  fulladder U8223 ( .a(n7631), .b(n7630), .ci(n7629), .co(n7661), .s(n6967) );
  fulladder U8224 ( .a(n7634), .b(n7633), .ci(n7632), .co(n7660), .s(n6952) );
  inv_1 U8225 ( .ip(n7635), .op(n7692) );
  fulladder U8226 ( .a(n7638), .b(n7637), .ci(n7636), .co(n7635), .s(n7639) );
  inv_1 U8227 ( .ip(n7639), .op(n7696) );
  fulladder U8228 ( .a(n7642), .b(n7641), .ci(n7640), .co(n7617), .s(n7658) );
  fulladder U8229 ( .a(n7645), .b(n7644), .ci(n7643), .co(n7636), .s(n7657) );
  fulladder U8230 ( .a(n7648), .b(n7647), .ci(n7646), .co(n7640), .s(n7666) );
  fulladder U8231 ( .a(n7651), .b(n7650), .ci(n7649), .co(n7641), .s(n7665) );
  fulladder U8232 ( .a(n7654), .b(n7653), .ci(n7652), .co(n7664), .s(n6946) );
  inv_1 U8233 ( .ip(n7655), .op(n7695) );
  fulladder U8234 ( .a(n7658), .b(n7657), .ci(n7656), .co(n7655), .s(n7659) );
  inv_1 U8235 ( .ip(n7659), .op(n7699) );
  fulladder U8236 ( .a(n7662), .b(n7661), .ci(n7660), .co(n7643), .s(n7663) );
  inv_1 U8237 ( .ip(n7663), .op(n7673) );
  fulladder U8238 ( .a(n7666), .b(n7665), .ci(n7664), .co(n7656), .s(n7667) );
  inv_1 U8239 ( .ip(n7667), .op(n7672) );
  fulladder U8240 ( .a(n7670), .b(n7669), .ci(n7668), .co(n7671), .s(n7678) );
  fulladder U8241 ( .a(n7673), .b(n7672), .ci(n7671), .co(n7698), .s(n7702) );
  fulladder U8242 ( .a(n7676), .b(n7675), .ci(n7674), .co(n7701), .s(
        \STAGE_1/M7/sum [1]) );
  fulladder U8243 ( .a(n7679), .b(n7678), .ci(n7677), .co(n7700), .s(n7676) );
  inv_1 U8244 ( .ip(n7680), .op(n14156) );
  fulladder U8245 ( .a(n7683), .b(n7682), .ci(n7681), .co(n14155), .s(n7570)
         );
  inv_1 U8246 ( .ip(n7684), .op(n14205) );
  fulladder U8247 ( .a(n7687), .b(n7686), .ci(n7685), .co(n14204), .s(n7189)
         );
  fulladder U8248 ( .a(n7690), .b(n7689), .ci(n7688), .co(n7680), .s(
        \STAGE_1/M7/sum [6]) );
  fulladder U8249 ( .a(n7693), .b(n7692), .ci(n7691), .co(n7688), .s(
        \STAGE_1/M7/sum [5]) );
  fulladder U8250 ( .a(n7696), .b(n7695), .ci(n7694), .co(n7691), .s(
        \STAGE_1/M7/sum [4]) );
  fulladder U8251 ( .a(n7699), .b(n7698), .ci(n7697), .co(n7694), .s(
        \STAGE_1/M7/sum [3]) );
  fulladder U8252 ( .a(n7702), .b(n7701), .ci(n7700), .co(n7697), .s(
        \STAGE_1/M7/sum [2]) );
  nand2_1 U8253 ( .ip1(\STAGE_1/weightReg [4]), .ip2(m1Inputs[117]), .op(n8171) );
  nor4_1 U8254 ( .ip1(n14783), .ip2(n8166), .ip3(n4624), .ip4(n14286), .op(
        n8214) );
  or2_1 U8255 ( .ip1(n8171), .ip2(n8214), .op(n7705) );
  or2_1 U8256 ( .ip1(n7703), .ip2(n8214), .op(n7704) );
  nand2_1 U8257 ( .ip1(n7705), .ip2(n7704), .op(n8213) );
  nor2_1 U8258 ( .ip1(n8177), .ip2(n6503), .op(n8215) );
  xnor2_1 U8259 ( .ip1(n8213), .ip2(n8215), .op(n8271) );
  and3_1 U8260 ( .ip1(n12578), .ip2(m1Inputs[121]), .ip3(n7706), .op(n8210) );
  inv_1 U8261 ( .ip(m1Inputs[121]), .op(n14372) );
  nor2_1 U8262 ( .ip1(n13646), .ip2(n14372), .op(n7707) );
  or2_1 U8263 ( .ip1(m1Inputs[118]), .ip2(n7707), .op(n7709) );
  or2_1 U8264 ( .ip1(n9733), .ip2(n7707), .op(n7708) );
  nand2_1 U8265 ( .ip1(n7709), .ip2(n7708), .op(n8208) );
  nor2_1 U8266 ( .ip1(n8210), .ip2(n8208), .op(n7710) );
  nand2_1 U8267 ( .ip1(m1Inputs[112]), .ip2(n14994), .op(n8207) );
  xor2_1 U8268 ( .ip1(n7710), .ip2(n8207), .op(n8270) );
  fulladder U8269 ( .a(n7713), .b(n7712), .ci(n7711), .co(n8269), .s(n4899) );
  inv_1 U8270 ( .ip(n7714), .op(n8296) );
  inv_1 U8271 ( .ip(n7715), .op(n7719) );
  nor2_1 U8272 ( .ip1(n7717), .ip2(n7716), .op(n7718) );
  nor2_1 U8273 ( .ip1(n7719), .ip2(n7718), .op(n8251) );
  nand2_1 U8274 ( .ip1(m1Inputs[115]), .ip2(n12981), .op(n8250) );
  nand2_1 U8275 ( .ip1(m1Inputs[114]), .ip2(\STAGE_1/weightReg [7]), .op(n8249) );
  inv_1 U8276 ( .ip(n7720), .op(n8287) );
  or2_1 U8277 ( .ip1(n7721), .ip2(n7722), .op(n7725) );
  or2_1 U8278 ( .ip1(n7723), .ip2(n7722), .op(n7724) );
  nand2_1 U8279 ( .ip1(n7725), .ip2(n7724), .op(n8248) );
  or2_1 U8280 ( .ip1(n7726), .ip2(n7727), .op(n7730) );
  or2_1 U8281 ( .ip1(n7728), .ip2(n7727), .op(n7729) );
  nand2_1 U8282 ( .ip1(n7730), .ip2(n7729), .op(n8247) );
  nand2_1 U8283 ( .ip1(n4619), .ip2(m1Inputs[119]), .op(n7732) );
  nor3_1 U8284 ( .ip1(n13709), .ip2(n14418), .ip3(n7731), .op(n8220) );
  or2_1 U8285 ( .ip1(n7732), .ip2(n8220), .op(n7734) );
  nand2_1 U8286 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[120]), .op(n8131) );
  or2_1 U8287 ( .ip1(n8131), .ip2(n8220), .op(n7733) );
  nand2_1 U8288 ( .ip1(n7734), .ip2(n7733), .op(n8218) );
  nand2_1 U8289 ( .ip1(column[113]), .ip2(n14768), .op(n8219) );
  xor2_1 U8290 ( .ip1(n8218), .ip2(n8219), .op(n8246) );
  inv_1 U8291 ( .ip(n7735), .op(n8286) );
  fulladder U8292 ( .a(n7738), .b(n7737), .ci(n7736), .co(n8285), .s(n7742) );
  fulladder U8293 ( .a(n7741), .b(n7740), .ci(n7739), .co(n8294), .s(n7743) );
  fulladder U8294 ( .a(n7744), .b(n7743), .ci(n7742), .co(n8292), .s(n7747) );
  fulladder U8295 ( .a(n7747), .b(n7746), .ci(n7745), .co(n8291), .s(
        \STAGE_1/M8/sum [0]) );
  inv_1 U8296 ( .ip(m1Inputs[126]), .op(n14434) );
  nor2_1 U8297 ( .ip1(n14434), .ip2(n14783), .op(n14282) );
  inv_1 U8298 ( .ip(m1Inputs[123]), .op(n14290) );
  nor2_1 U8299 ( .ip1(n14290), .ip2(n14384), .op(n14281) );
  nand2_1 U8300 ( .ip1(n12578), .ip2(m1Inputs[127]), .op(n14280) );
  nand2_1 U8301 ( .ip1(m1Inputs[125]), .ip2(n14369), .op(n14278) );
  nor2_1 U8302 ( .ip1(n7790), .ip2(n14853), .op(n14277) );
  nand2_1 U8303 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[121]), .op(
        n14276) );
  inv_1 U8304 ( .ip(n7748), .op(n14325) );
  nor2_1 U8305 ( .ip1(n14902), .ip2(n14286), .op(n7775) );
  nor2_1 U8306 ( .ip1(n13594), .ip2(n8172), .op(n7768) );
  or2_1 U8307 ( .ip1(m1Inputs[117]), .ip2(n7768), .op(n7750) );
  or2_1 U8308 ( .ip1(n14847), .ip2(n7768), .op(n7749) );
  nand2_1 U8309 ( .ip1(n7750), .ip2(n7749), .op(n7788) );
  nor3_1 U8310 ( .ip1(n7788), .ip2(n7790), .ip3(n14340), .op(n7751) );
  nor2_1 U8311 ( .ip1(n13594), .ip2(n14286), .op(n7886) );
  and3_1 U8312 ( .ip1(\STAGE_1/weightReg [11]), .ip2(m1Inputs[118]), .ip3(
        n7886), .op(n7789) );
  or2_1 U8313 ( .ip1(n7751), .ip2(n7789), .op(n7774) );
  nor2_1 U8314 ( .ip1(n13854), .ip2(n14434), .op(n7785) );
  nand2_1 U8315 ( .ip1(column[120]), .ip2(n14768), .op(n7784) );
  inv_1 U8316 ( .ip(m1Inputs[119]), .op(n14339) );
  nor2_1 U8317 ( .ip1(n13766), .ip2(n14339), .op(n7783) );
  nor2_1 U8318 ( .ip1(n14373), .ip2(n14286), .op(n14320) );
  nor2_1 U8319 ( .ip1(n14902), .ip2(n8172), .op(n14319) );
  nor2_1 U8320 ( .ip1(n12083), .ip2(n14418), .op(n7760) );
  and2_1 U8321 ( .ip1(column[121]), .ip2(n13498), .op(n7759) );
  inv_1 U8322 ( .ip(n7784), .op(n7758) );
  nor2_1 U8323 ( .ip1(n14372), .ip2(n14289), .op(n7776) );
  and3_1 U8324 ( .ip1(m1Inputs[122]), .ip2(n14835), .ip3(n7776), .op(n7755) );
  inv_1 U8325 ( .ip(m1Inputs[122]), .op(n14433) );
  nor2_1 U8326 ( .ip1(n14433), .ip2(n14836), .op(n7763) );
  or2_1 U8327 ( .ip1(n4627), .ip2(n7763), .op(n7753) );
  or2_1 U8328 ( .ip1(m1Inputs[121]), .ip2(n7763), .op(n7752) );
  nand2_1 U8329 ( .ip1(n7753), .ip2(n7752), .op(n7754) );
  nor2_1 U8330 ( .ip1(n7755), .ip2(n7754), .op(n7794) );
  or2_1 U8331 ( .ip1(n7794), .ip2(n7755), .op(n7757) );
  nor2_1 U8332 ( .ip1(n14290), .ip2(n4624), .op(n7793) );
  or2_1 U8333 ( .ip1(n7793), .ip2(n7755), .op(n7756) );
  nand2_1 U8334 ( .ip1(n7757), .ip2(n7756), .op(n7798) );
  nand2_1 U8335 ( .ip1(n13614), .ip2(m1Inputs[125]), .op(n7907) );
  inv_1 U8336 ( .ip(m1Inputs[127]), .op(n14287) );
  nor2_1 U8337 ( .ip1(n13570), .ip2(n14287), .op(n7804) );
  nand2_1 U8338 ( .ip1(m1Inputs[114]), .ip2(\STAGE_1/weightReg [14]), .op(
        n7803) );
  fulladder U8339 ( .a(n7760), .b(n7759), .ci(n7758), .co(n14318), .s(n7761)
         );
  inv_1 U8340 ( .ip(n7761), .op(n7796) );
  inv_1 U8341 ( .ip(n7762), .op(n14322) );
  nand2_1 U8342 ( .ip1(m1Inputs[123]), .ip2(\STAGE_1/weightReg [6]), .op(n7764) );
  and2_1 U8343 ( .ip1(n7763), .ip2(n14281), .op(n7816) );
  or2_1 U8344 ( .ip1(n7764), .ip2(n7816), .op(n7767) );
  nand2_1 U8345 ( .ip1(m1Inputs[122]), .ip2(n14835), .op(n7765) );
  or2_1 U8346 ( .ip1(n7765), .ip2(n7816), .op(n7766) );
  nand2_1 U8347 ( .ip1(n7767), .ip2(n7766), .op(n7815) );
  inv_1 U8348 ( .ip(m1Inputs[124]), .op(n14517) );
  nor2_1 U8349 ( .ip1(n14517), .ip2(n12746), .op(n7817) );
  xor2_1 U8350 ( .ip1(n7815), .ip2(n7817), .op(n7801) );
  and3_1 U8351 ( .ip1(\STAGE_1/weightReg [11]), .ip2(m1Inputs[119]), .ip3(
        n7768), .op(n7826) );
  nor2_1 U8352 ( .ip1(n13579), .ip2(n8172), .op(n7769) );
  or2_1 U8353 ( .ip1(m1Inputs[119]), .ip2(n7769), .op(n7771) );
  or2_1 U8354 ( .ip1(n14876), .ip2(n7769), .op(n7770) );
  nand2_1 U8355 ( .ip1(n7771), .ip2(n7770), .op(n7772) );
  nor2_1 U8356 ( .ip1(n7826), .ip2(n7772), .op(n7825) );
  nor2_1 U8357 ( .ip1(n14340), .ip2(n8166), .op(n7827) );
  xor2_1 U8358 ( .ip1(n7825), .ip2(n7827), .op(n7800) );
  nor2_1 U8359 ( .ip1(n14517), .ip2(n14783), .op(n7806) );
  nor2_1 U8360 ( .ip1(n6503), .ip2(n14418), .op(n14302) );
  nand2_1 U8361 ( .ip1(m1Inputs[113]), .ip2(\STAGE_1/weightReg [15]), .op(
        n7805) );
  fulladder U8362 ( .a(n7775), .b(n7774), .ci(n7773), .co(n14324), .s(n7895)
         );
  nand2_1 U8363 ( .ip1(m1Inputs[121]), .ip2(\STAGE_1/weightReg [4]), .op(n7936) );
  nor3_1 U8364 ( .ip1(n14290), .ip2(n14289), .ip3(n7936), .op(n7780) );
  or2_1 U8365 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n7776), .op(n7778) );
  or2_1 U8366 ( .ip1(m1Inputs[123]), .ip2(n7776), .op(n7777) );
  nand2_1 U8367 ( .ip1(n7778), .ip2(n7777), .op(n7779) );
  nor2_1 U8368 ( .ip1(n7780), .ip2(n7779), .op(n7857) );
  or2_1 U8369 ( .ip1(n7857), .ip2(n7780), .op(n7782) );
  nor2_1 U8370 ( .ip1(n8177), .ip2(n14842), .op(n7856) );
  or2_1 U8371 ( .ip1(n7856), .ip2(n7780), .op(n7781) );
  nand2_1 U8372 ( .ip1(n7782), .ip2(n7781), .op(n7863) );
  nand2_1 U8373 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[124]), .op(n8012) );
  nor2_1 U8374 ( .ip1(n10476), .ip2(n14287), .op(n7852) );
  nand2_1 U8375 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[118]), .op(n7851) );
  fulladder U8376 ( .a(n7785), .b(n7784), .ci(n7783), .co(n7773), .s(n7786) );
  inv_1 U8377 ( .ip(n7786), .op(n7861) );
  inv_1 U8378 ( .ip(n7787), .op(n7894) );
  nor2_1 U8379 ( .ip1(n7789), .ip2(n7788), .op(n7792) );
  nor2_1 U8380 ( .ip1(n7790), .ip2(n14340), .op(n7791) );
  xor2_1 U8381 ( .ip1(n7792), .ip2(n7791), .op(n7860) );
  xor2_1 U8382 ( .ip1(n7794), .ip2(n7793), .op(n7859) );
  nor2_1 U8383 ( .ip1(n14433), .ip2(n12746), .op(n7855) );
  nand2_1 U8384 ( .ip1(m1Inputs[112]), .ip2(\STAGE_1/weightReg [15]), .op(
        n7854) );
  inv_1 U8385 ( .ip(n7795), .op(n14334) );
  fulladder U8386 ( .a(n7798), .b(n7797), .ci(n7796), .co(n7762), .s(n7899) );
  fulladder U8387 ( .a(n7801), .b(n7800), .ci(n7799), .co(n14321), .s(n7802)
         );
  inv_1 U8388 ( .ip(n7802), .op(n7898) );
  fulladder U8389 ( .a(n7907), .b(n7804), .ci(n7803), .co(n7797), .s(n7902) );
  fulladder U8390 ( .a(n7806), .b(n14302), .ci(n7805), .co(n7799), .s(n7807)
         );
  inv_1 U8391 ( .ip(n7807), .op(n7901) );
  nand2_1 U8392 ( .ip1(n4619), .ip2(m1Inputs[124]), .op(n7808) );
  inv_1 U8393 ( .ip(m1Inputs[125]), .op(n14419) );
  nand2_1 U8394 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[124]), .op(n7949) );
  nor3_1 U8395 ( .ip1(n13709), .ip2(n14419), .ip3(n7949), .op(n7811) );
  or2_1 U8396 ( .ip1(n7808), .ip2(n7811), .op(n7810) );
  nand2_1 U8397 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[125]), .op(n7839) );
  or2_1 U8398 ( .ip1(n7839), .ip2(n7811), .op(n7809) );
  nand2_1 U8399 ( .ip1(n7810), .ip2(n7809), .op(n7943) );
  or2_1 U8400 ( .ip1(n7943), .ip2(n7811), .op(n7814) );
  nand2_1 U8401 ( .ip1(column[118]), .ip2(n13498), .op(n7942) );
  inv_1 U8402 ( .ip(n7942), .op(n7812) );
  or2_1 U8403 ( .ip1(n7812), .ip2(n7811), .op(n7813) );
  nand2_1 U8404 ( .ip1(n7814), .ip2(n7813), .op(n7927) );
  nand2_1 U8405 ( .ip1(m1Inputs[115]), .ip2(\STAGE_1/weightReg [12]), .op(
        n7926) );
  nand2_1 U8406 ( .ip1(n14847), .ip2(m1Inputs[116]), .op(n7925) );
  or2_1 U8407 ( .ip1(n7815), .ip2(n7816), .op(n7819) );
  or2_1 U8408 ( .ip1(n7817), .ip2(n7816), .op(n7818) );
  nand2_1 U8409 ( .ip1(n7819), .ip2(n7818), .op(n14316) );
  nand2_1 U8410 ( .ip1(m1Inputs[125]), .ip2(n13637), .op(n7832) );
  nor2_1 U8411 ( .ip1(n8099), .ip2(n14853), .op(n7831) );
  nand2_1 U8412 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[121]), .op(n7830) );
  nand2_1 U8413 ( .ip1(m1Inputs[122]), .ip2(n14975), .op(n7821) );
  nand2_1 U8414 ( .ip1(m1Inputs[120]), .ip2(\STAGE_1/weightReg [10]), .op(
        n7820) );
  xor2_1 U8415 ( .ip1(n7821), .ip2(n7820), .op(n14303) );
  nand2_1 U8416 ( .ip1(column[122]), .ip2(n14768), .op(n14304) );
  xor2_1 U8417 ( .ip1(n14303), .ip2(n14304), .op(n14314) );
  nand2_1 U8418 ( .ip1(m1Inputs[119]), .ip2(n12981), .op(n7929) );
  nor3_1 U8419 ( .ip1(n14824), .ip2(n14517), .ip3(n7929), .op(n14312) );
  nor2_1 U8420 ( .ip1(n14824), .ip2(n14339), .op(n14374) );
  or2_1 U8421 ( .ip1(n13749), .ip2(n14374), .op(n7823) );
  or2_1 U8422 ( .ip1(m1Inputs[124]), .ip2(n14374), .op(n7822) );
  nand2_1 U8423 ( .ip1(n7823), .ip2(n7822), .op(n14310) );
  nor2_1 U8424 ( .ip1(n14312), .ip2(n14310), .op(n7824) );
  nand2_1 U8425 ( .ip1(n14816), .ip2(m1Inputs[116]), .op(n14309) );
  xor2_1 U8426 ( .ip1(n7824), .ip2(n14309), .op(n14294) );
  or2_1 U8427 ( .ip1(n7825), .ip2(n7826), .op(n7829) );
  or2_1 U8428 ( .ip1(n7827), .ip2(n7826), .op(n7828) );
  nand2_1 U8429 ( .ip1(n7829), .ip2(n7828), .op(n14293) );
  nor2_1 U8430 ( .ip1(n13854), .ip2(n14287), .op(n7834) );
  nand2_1 U8431 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[126]), .op(n7881) );
  nand2_1 U8432 ( .ip1(m1Inputs[115]), .ip2(\STAGE_1/weightReg [14]), .op(
        n7833) );
  fulladder U8433 ( .a(n7832), .b(n7831), .ci(n7830), .co(n14315), .s(n7850)
         );
  fulladder U8434 ( .a(n7834), .b(n7881), .ci(n7833), .co(n14292), .s(n7849)
         );
  nor2_1 U8435 ( .ip1(n14339), .ip2(n14368), .op(n7873) );
  and2_1 U8436 ( .ip1(n14302), .ip2(n7873), .op(n7878) );
  nor2_1 U8437 ( .ip1(n14418), .ip2(n14384), .op(n7835) );
  or2_1 U8438 ( .ip1(m1Inputs[119]), .ip2(n7835), .op(n7837) );
  or2_1 U8439 ( .ip1(n14838), .ip2(n7835), .op(n7836) );
  nand2_1 U8440 ( .ip1(n7837), .ip2(n7836), .op(n7877) );
  nand2_1 U8441 ( .ip1(m1Inputs[114]), .ip2(\STAGE_1/weightReg [13]), .op(
        n7879) );
  nor2_1 U8442 ( .ip1(n7877), .ip2(n7879), .op(n7838) );
  nor2_1 U8443 ( .ip1(n7878), .ip2(n7838), .op(n7868) );
  nand2_1 U8444 ( .ip1(n4672), .ip2(m1Inputs[125]), .op(n7840) );
  nor3_1 U8445 ( .ip1(n13709), .ip2(n14434), .ip3(n7839), .op(n7844) );
  or2_1 U8446 ( .ip1(n7840), .ip2(n7844), .op(n7843) );
  nand2_1 U8447 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[126]), .op(n7841) );
  or2_1 U8448 ( .ip1(n7841), .ip2(n7844), .op(n7842) );
  nand2_1 U8449 ( .ip1(n7843), .ip2(n7842), .op(n7892) );
  or2_1 U8450 ( .ip1(n7892), .ip2(n7844), .op(n7847) );
  nand2_1 U8451 ( .ip1(column[119]), .ip2(n13498), .op(n7891) );
  inv_1 U8452 ( .ip(n7891), .op(n7845) );
  or2_1 U8453 ( .ip1(n7845), .ip2(n7844), .op(n7846) );
  nand2_1 U8454 ( .ip1(n7847), .ip2(n7846), .op(n7867) );
  nand2_1 U8455 ( .ip1(n15025), .ip2(m1Inputs[116]), .op(n7866) );
  fulladder U8456 ( .a(n7850), .b(n7849), .ci(n7848), .co(n14299), .s(n7959)
         );
  fulladder U8457 ( .a(n8012), .b(n7852), .ci(n7851), .co(n7862), .s(n7853) );
  inv_1 U8458 ( .ip(n7853), .op(n7972) );
  fulladder U8459 ( .a(n7855), .b(n7886), .ci(n7854), .co(n7858), .s(n7971) );
  xor2_1 U8460 ( .ip1(n7857), .ip2(n7856), .op(n7970) );
  fulladder U8461 ( .a(n7860), .b(n7859), .ci(n7858), .co(n7893), .s(n7967) );
  fulladder U8462 ( .a(n7863), .b(n7862), .ci(n7861), .co(n7787), .s(n7864) );
  inv_1 U8463 ( .ip(n7864), .op(n7966) );
  inv_1 U8464 ( .ip(n7865), .op(n7958) );
  fulladder U8465 ( .a(n7868), .b(n7867), .ci(n7866), .co(n7848), .s(n7965) );
  nor3_1 U8466 ( .ip1(n14433), .ip2(n4624), .ip3(n7936), .op(n7992) );
  nor2_1 U8467 ( .ip1(n14372), .ip2(n12746), .op(n7869) );
  or2_1 U8468 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n7869), .op(n7871) );
  or2_1 U8469 ( .ip1(m1Inputs[122]), .ip2(n7869), .op(n7870) );
  nand2_1 U8470 ( .ip1(n7871), .ip2(n7870), .op(n7991) );
  nand2_1 U8471 ( .ip1(n14838), .ip2(m1Inputs[118]), .op(n7993) );
  nor2_1 U8472 ( .ip1(n7991), .ip2(n7993), .op(n7872) );
  nor2_1 U8473 ( .ip1(n7992), .ip2(n7872), .op(n7921) );
  nor3_1 U8474 ( .ip1(n14418), .ip2(n14384), .ip3(n7929), .op(n7904) );
  or2_1 U8475 ( .ip1(n13749), .ip2(n7873), .op(n7875) );
  or2_1 U8476 ( .ip1(m1Inputs[120]), .ip2(n7873), .op(n7874) );
  nand2_1 U8477 ( .ip1(n7875), .ip2(n7874), .op(n7903) );
  nand2_1 U8478 ( .ip1(m1Inputs[113]), .ip2(\STAGE_1/weightReg [13]), .op(
        n7905) );
  nor2_1 U8479 ( .ip1(n7903), .ip2(n7905), .op(n7876) );
  nor2_1 U8480 ( .ip1(n7904), .ip2(n7876), .op(n7920) );
  nor2_1 U8481 ( .ip1(n7878), .ip2(n7877), .op(n7880) );
  xor2_1 U8482 ( .ip1(n7880), .ip2(n7879), .op(n7919) );
  nand2_1 U8483 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[123]), .op(n8089) );
  nor2_1 U8484 ( .ip1(n8089), .ip2(n7881), .op(n7996) );
  nor2_1 U8485 ( .ip1(n13487), .ip2(n14290), .op(n7882) );
  or2_1 U8486 ( .ip1(m1Inputs[126]), .ip2(n7882), .op(n7884) );
  or2_1 U8487 ( .ip1(n13803), .ip2(n7882), .op(n7883) );
  nand2_1 U8488 ( .ip1(n7884), .ip2(n7883), .op(n7995) );
  nand2_1 U8489 ( .ip1(m1Inputs[112]), .ip2(\STAGE_1/weightReg [14]), .op(
        n7997) );
  nor2_1 U8490 ( .ip1(n7995), .ip2(n7997), .op(n7885) );
  nor2_1 U8491 ( .ip1(n7996), .ip2(n7885), .op(n7924) );
  nor2_1 U8492 ( .ip1(n13766), .ip2(n8166), .op(n7944) );
  and2_1 U8493 ( .ip1(n7944), .ip2(n7886), .op(n7916) );
  nor2_1 U8494 ( .ip1(n13766), .ip2(n14286), .op(n7887) );
  or2_1 U8495 ( .ip1(m1Inputs[116]), .ip2(n7887), .op(n7889) );
  or2_1 U8496 ( .ip1(n14876), .ip2(n7887), .op(n7888) );
  nand2_1 U8497 ( .ip1(n7889), .ip2(n7888), .op(n7915) );
  nand2_1 U8498 ( .ip1(m1Inputs[114]), .ip2(\STAGE_1/weightReg [12]), .op(
        n7917) );
  nor2_1 U8499 ( .ip1(n7915), .ip2(n7917), .op(n7890) );
  nor2_1 U8500 ( .ip1(n7916), .ip2(n7890), .op(n7923) );
  xor2_1 U8501 ( .ip1(n7892), .ip2(n7891), .op(n7922) );
  fulladder U8502 ( .a(n7895), .b(n7894), .ci(n7893), .co(n14295), .s(n7896)
         );
  inv_1 U8503 ( .ip(n7896), .op(n7962) );
  fulladder U8504 ( .a(n7899), .b(n7898), .ci(n7897), .co(n14330), .s(n7961)
         );
  fulladder U8505 ( .a(n7902), .b(n7901), .ci(n7900), .co(n7897), .s(n8028) );
  nor2_1 U8506 ( .ip1(n7904), .ip2(n7903), .op(n7906) );
  xor2_1 U8507 ( .ip1(n7906), .ip2(n7905), .op(n8044) );
  nand2_1 U8508 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[122]), .op(n8142) );
  nor2_1 U8509 ( .ip1(n8142), .ip2(n7907), .op(n7912) );
  nor2_1 U8510 ( .ip1(n13082), .ip2(n14433), .op(n7908) );
  or2_1 U8511 ( .ip1(m1Inputs[125]), .ip2(n7908), .op(n7910) );
  or2_1 U8512 ( .ip1(n13803), .ip2(n7908), .op(n7909) );
  nand2_1 U8513 ( .ip1(n7910), .ip2(n7909), .op(n7911) );
  nor2_1 U8514 ( .ip1(n7912), .ip2(n7911), .op(n8051) );
  or2_1 U8515 ( .ip1(n8051), .ip2(n7912), .op(n7914) );
  nor2_1 U8516 ( .ip1(n8145), .ip2(n14340), .op(n8050) );
  or2_1 U8517 ( .ip1(n8050), .ip2(n7912), .op(n7913) );
  nand2_1 U8518 ( .ip1(n7914), .ip2(n7913), .op(n8043) );
  nor2_1 U8519 ( .ip1(n7916), .ip2(n7915), .op(n7918) );
  xor2_1 U8520 ( .ip1(n7918), .ip2(n7917), .op(n8042) );
  fulladder U8521 ( .a(n7921), .b(n7920), .ci(n7919), .co(n7964), .s(n8039) );
  fulladder U8522 ( .a(n7924), .b(n7923), .ci(n7922), .co(n7963), .s(n8038) );
  fulladder U8523 ( .a(n7927), .b(n7926), .ci(n7925), .co(n7900), .s(n8036) );
  nand2_1 U8524 ( .ip1(m1Inputs[118]), .ip2(\STAGE_1/weightReg [7]), .op(n7928) );
  nand2_1 U8525 ( .ip1(m1Inputs[118]), .ip2(n12981), .op(n7983) );
  nor3_1 U8526 ( .ip1(n14339), .ip2(n14368), .ip3(n7983), .op(n7932) );
  or2_1 U8527 ( .ip1(n7928), .ip2(n7932), .op(n7931) );
  or2_1 U8528 ( .ip1(n7929), .ip2(n7932), .op(n7930) );
  nand2_1 U8529 ( .ip1(n7931), .ip2(n7930), .op(n8055) );
  or2_1 U8530 ( .ip1(n8055), .ip2(n7932), .op(n7934) );
  nor2_1 U8531 ( .ip1(n8099), .ip2(n14824), .op(n8054) );
  or2_1 U8532 ( .ip1(n8054), .ip2(n7932), .op(n7933) );
  nand2_1 U8533 ( .ip1(n7934), .ip2(n7933), .op(n8004) );
  nand2_1 U8534 ( .ip1(m1Inputs[120]), .ip2(n14369), .op(n7935) );
  nand2_1 U8535 ( .ip1(m1Inputs[120]), .ip2(n13637), .op(n8006) );
  nor3_1 U8536 ( .ip1(n14372), .ip2(n12746), .ip3(n8006), .op(n7939) );
  or2_1 U8537 ( .ip1(n7935), .ip2(n7939), .op(n7938) );
  or2_1 U8538 ( .ip1(n7936), .ip2(n7939), .op(n7937) );
  nand2_1 U8539 ( .ip1(n7938), .ip2(n7937), .op(n8053) );
  or2_1 U8540 ( .ip1(n8053), .ip2(n7939), .op(n7941) );
  nor2_1 U8541 ( .ip1(n8177), .ip2(n14188), .op(n8052) );
  or2_1 U8542 ( .ip1(n8052), .ip2(n7939), .op(n7940) );
  nand2_1 U8543 ( .ip1(n7941), .ip2(n7940), .op(n8003) );
  xor2_1 U8544 ( .ip1(n7943), .ip2(n7942), .op(n8002) );
  nand2_1 U8545 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[116]), .op(n8151) );
  nor3_1 U8546 ( .ip1(n12083), .ip2(n14286), .ip3(n8151), .op(n8018) );
  or2_1 U8547 ( .ip1(m1Inputs[117]), .ip2(n7944), .op(n7946) );
  or2_1 U8548 ( .ip1(n14838), .ip2(n7944), .op(n7945) );
  nand2_1 U8549 ( .ip1(n7946), .ip2(n7945), .op(n8017) );
  nand2_1 U8550 ( .ip1(m1Inputs[115]), .ip2(\STAGE_1/weightReg [10]), .op(
        n8019) );
  nor2_1 U8551 ( .ip1(n8017), .ip2(n8019), .op(n7947) );
  nor2_1 U8552 ( .ip1(n8018), .ip2(n7947), .op(n8001) );
  nand2_1 U8553 ( .ip1(n4619), .ip2(m1Inputs[123]), .op(n7948) );
  nand2_1 U8554 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[123]), .op(n7975) );
  nor3_1 U8555 ( .ip1(n13709), .ip2(n14517), .ip3(n7975), .op(n7952) );
  or2_1 U8556 ( .ip1(n7948), .ip2(n7952), .op(n7951) );
  or2_1 U8557 ( .ip1(n7949), .ip2(n7952), .op(n7950) );
  nand2_1 U8558 ( .ip1(n7951), .ip2(n7950), .op(n7990) );
  or2_1 U8559 ( .ip1(n7990), .ip2(n7952), .op(n7955) );
  nand2_1 U8560 ( .ip1(column[117]), .ip2(n14768), .op(n7989) );
  inv_1 U8561 ( .ip(n7989), .op(n7953) );
  or2_1 U8562 ( .ip1(n7953), .ip2(n7952), .op(n7954) );
  nand2_1 U8563 ( .ip1(n7955), .ip2(n7954), .op(n8000) );
  nand2_1 U8564 ( .ip1(m1Inputs[115]), .ip2(\STAGE_1/weightReg [11]), .op(
        n7999) );
  inv_1 U8565 ( .ip(n7956), .op(n14338) );
  fulladder U8566 ( .a(n7959), .b(n7958), .ci(n7957), .co(n14328), .s(n8024)
         );
  fulladder U8567 ( .a(n7962), .b(n7961), .ci(n7960), .co(n14332), .s(n8023)
         );
  fulladder U8568 ( .a(n7965), .b(n7964), .ci(n7963), .co(n7957), .s(n8032) );
  fulladder U8569 ( .a(n7968), .b(n7967), .ci(n7966), .co(n7865), .s(n7969) );
  inv_1 U8570 ( .ip(n7969), .op(n8031) );
  fulladder U8571 ( .a(n7972), .b(n7971), .ci(n7970), .co(n7968), .s(n7973) );
  inv_1 U8572 ( .ip(n7973), .op(n8061) );
  nand2_1 U8573 ( .ip1(n4619), .ip2(m1Inputs[122]), .op(n7974) );
  nand2_1 U8574 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[122]), .op(n8080) );
  nor3_1 U8575 ( .ip1(n13709), .ip2(n14290), .ip3(n8080), .op(n7978) );
  or2_1 U8576 ( .ip1(n7974), .ip2(n7978), .op(n7977) );
  or2_1 U8577 ( .ip1(n7975), .ip2(n7978), .op(n7976) );
  nand2_1 U8578 ( .ip1(n7977), .ip2(n7976), .op(n8104) );
  or2_1 U8579 ( .ip1(n8104), .ip2(n7978), .op(n7981) );
  nand2_1 U8580 ( .ip1(column[116]), .ip2(n13859), .op(n8103) );
  inv_1 U8581 ( .ip(n8103), .op(n7979) );
  or2_1 U8582 ( .ip1(n7979), .ip2(n7978), .op(n7980) );
  nand2_1 U8583 ( .ip1(n7981), .ip2(n7980), .op(n8078) );
  nand2_1 U8584 ( .ip1(n14835), .ip2(m1Inputs[117]), .op(n7982) );
  nand2_1 U8585 ( .ip1(n13749), .ip2(m1Inputs[117]), .op(n8096) );
  nor3_1 U8586 ( .ip1(n8172), .ip2(n14368), .ip3(n8096), .op(n7986) );
  or2_1 U8587 ( .ip1(n7982), .ip2(n7986), .op(n7985) );
  or2_1 U8588 ( .ip1(n7983), .ip2(n7986), .op(n7984) );
  nand2_1 U8589 ( .ip1(n7985), .ip2(n7984), .op(n8115) );
  or2_1 U8590 ( .ip1(n8115), .ip2(n7986), .op(n7988) );
  nor2_1 U8591 ( .ip1(n8099), .ip2(n13594), .op(n8114) );
  or2_1 U8592 ( .ip1(n8114), .ip2(n7986), .op(n7987) );
  nand2_1 U8593 ( .ip1(n7988), .ip2(n7987), .op(n8077) );
  xor2_1 U8594 ( .ip1(n7990), .ip2(n7989), .op(n8076) );
  nor2_1 U8595 ( .ip1(n7992), .ip2(n7991), .op(n7994) );
  xor2_1 U8596 ( .ip1(n7994), .ip2(n7993), .op(n8047) );
  nor2_1 U8597 ( .ip1(n7996), .ip2(n7995), .op(n7998) );
  xor2_1 U8598 ( .ip1(n7998), .ip2(n7997), .op(n8046) );
  fulladder U8599 ( .a(n8001), .b(n8000), .ci(n7999), .co(n8034), .s(n8068) );
  fulladder U8600 ( .a(n8004), .b(n8003), .ci(n8002), .co(n8035), .s(n8067) );
  nand2_1 U8601 ( .ip1(m1Inputs[119]), .ip2(n14369), .op(n8005) );
  nand2_1 U8602 ( .ip1(m1Inputs[119]), .ip2(n13637), .op(n8106) );
  nor3_1 U8603 ( .ip1(n14418), .ip2(n13835), .ip3(n8106), .op(n8009) );
  or2_1 U8604 ( .ip1(n8005), .ip2(n8009), .op(n8008) );
  or2_1 U8605 ( .ip1(n8006), .ip2(n8009), .op(n8007) );
  nand2_1 U8606 ( .ip1(n8008), .ip2(n8007), .op(n8113) );
  or2_1 U8607 ( .ip1(n8113), .ip2(n8009), .op(n8011) );
  nor2_1 U8608 ( .ip1(n8177), .ip2(n14824), .op(n8112) );
  or2_1 U8609 ( .ip1(n8112), .ip2(n8009), .op(n8010) );
  nand2_1 U8610 ( .ip1(n8011), .ip2(n8010), .op(n8071) );
  nor3_1 U8611 ( .ip1(n10476), .ip2(n14372), .ip3(n8012), .op(n8153) );
  nor2_1 U8612 ( .ip1(n13487), .ip2(n14372), .op(n8013) );
  or2_1 U8613 ( .ip1(m1Inputs[124]), .ip2(n8013), .op(n8015) );
  or2_1 U8614 ( .ip1(n13803), .ip2(n8013), .op(n8014) );
  nand2_1 U8615 ( .ip1(n8015), .ip2(n8014), .op(n8152) );
  nand2_1 U8616 ( .ip1(m1Inputs[112]), .ip2(\STAGE_1/weightReg [12]), .op(
        n8154) );
  nor2_1 U8617 ( .ip1(n8152), .ip2(n8154), .op(n8016) );
  nor2_1 U8618 ( .ip1(n8153), .ip2(n8016), .op(n8070) );
  nor2_1 U8619 ( .ip1(n8018), .ip2(n8017), .op(n8020) );
  xor2_1 U8620 ( .ip1(n8020), .ip2(n8019), .op(n8069) );
  inv_1 U8621 ( .ip(n8021), .op(n14337) );
  fulladder U8622 ( .a(n8024), .b(n8023), .ci(n8022), .co(n8021), .s(n8025) );
  inv_1 U8623 ( .ip(n8025), .op(n8299) );
  fulladder U8624 ( .a(n8028), .b(n8027), .ci(n8026), .co(n7960), .s(n8029) );
  inv_1 U8625 ( .ip(n8029), .op(n8058) );
  fulladder U8626 ( .a(n8032), .b(n8031), .ci(n8030), .co(n8022), .s(n8033) );
  inv_1 U8627 ( .ip(n8033), .op(n8057) );
  fulladder U8628 ( .a(n8036), .b(n8035), .ci(n8034), .co(n8026), .s(n8037) );
  inv_1 U8629 ( .ip(n8037), .op(n8064) );
  fulladder U8630 ( .a(n8040), .b(n8039), .ci(n8038), .co(n8027), .s(n8041) );
  inv_1 U8631 ( .ip(n8041), .op(n8063) );
  fulladder U8632 ( .a(n8044), .b(n8043), .ci(n8042), .co(n8040), .s(n8045) );
  inv_1 U8633 ( .ip(n8045), .op(n8123) );
  fulladder U8634 ( .a(n8048), .b(n8047), .ci(n8046), .co(n8060), .s(n8049) );
  inv_1 U8635 ( .ip(n8049), .op(n8122) );
  xor2_1 U8636 ( .ip1(n8051), .ip2(n8050), .op(n8074) );
  xor2_1 U8637 ( .ip1(n8053), .ip2(n8052), .op(n8073) );
  xor2_1 U8638 ( .ip1(n8055), .ip2(n8054), .op(n8072) );
  fulladder U8639 ( .a(n8058), .b(n8057), .ci(n8056), .co(n8298), .s(n8302) );
  fulladder U8640 ( .a(n8061), .b(n8060), .ci(n8059), .co(n8030), .s(n8119) );
  fulladder U8641 ( .a(n8064), .b(n8063), .ci(n8062), .co(n8056), .s(n8065) );
  inv_1 U8642 ( .ip(n8065), .op(n8118) );
  fulladder U8643 ( .a(n8068), .b(n8067), .ci(n8066), .co(n8059), .s(n8127) );
  fulladder U8644 ( .a(n8071), .b(n8070), .ci(n8069), .co(n8066), .s(n8190) );
  fulladder U8645 ( .a(n8074), .b(n8073), .ci(n8072), .co(n8121), .s(n8075) );
  inv_1 U8646 ( .ip(n8075), .op(n8189) );
  fulladder U8647 ( .a(n8078), .b(n8077), .ci(n8076), .co(n8048), .s(n8188) );
  nand2_1 U8648 ( .ip1(n4619), .ip2(m1Inputs[121]), .op(n8079) );
  nand2_1 U8649 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[121]), .op(n8133) );
  nor3_1 U8650 ( .ip1(n13709), .ip2(n14433), .ip3(n8133), .op(n8083) );
  or2_1 U8651 ( .ip1(n8079), .ip2(n8083), .op(n8082) );
  or2_1 U8652 ( .ip1(n8080), .ip2(n8083), .op(n8081) );
  nand2_1 U8653 ( .ip1(n8082), .ip2(n8081), .op(n8182) );
  or2_1 U8654 ( .ip1(n8182), .ip2(n8083), .op(n8086) );
  nand2_1 U8655 ( .ip1(column[115]), .ip2(n14768), .op(n8181) );
  inv_1 U8656 ( .ip(n8181), .op(n8084) );
  or2_1 U8657 ( .ip1(n8084), .ip2(n8083), .op(n8085) );
  nand2_1 U8658 ( .ip1(n8086), .ip2(n8085), .op(n8150) );
  nand2_1 U8659 ( .ip1(m1Inputs[115]), .ip2(n14994), .op(n8149) );
  nand2_1 U8660 ( .ip1(n13614), .ip2(m1Inputs[120]), .op(n8088) );
  nor3_1 U8661 ( .ip1(n13082), .ip2(n14290), .ip3(n8087), .op(n8092) );
  or2_1 U8662 ( .ip1(n8088), .ip2(n8092), .op(n8091) );
  or2_1 U8663 ( .ip1(n8089), .ip2(n8092), .op(n8090) );
  nand2_1 U8664 ( .ip1(n8091), .ip2(n8090), .op(n8164) );
  or2_1 U8665 ( .ip1(n8164), .ip2(n8092), .op(n8094) );
  nor2_1 U8666 ( .ip1(n8145), .ip2(n14824), .op(n8163) );
  or2_1 U8667 ( .ip1(n8163), .ip2(n8092), .op(n8093) );
  nand2_1 U8668 ( .ip1(n8094), .ip2(n8093), .op(n8158) );
  nand2_1 U8669 ( .ip1(m1Inputs[116]), .ip2(n14835), .op(n8095) );
  nor2_1 U8670 ( .ip1(n8166), .ip2(n14836), .op(n8167) );
  and3_1 U8671 ( .ip1(n4627), .ip2(m1Inputs[117]), .ip3(n8167), .op(n8100) );
  or2_1 U8672 ( .ip1(n8095), .ip2(n8100), .op(n8098) );
  or2_1 U8673 ( .ip1(n8096), .ip2(n8100), .op(n8097) );
  nand2_1 U8674 ( .ip1(n8098), .ip2(n8097), .op(n8160) );
  or2_1 U8675 ( .ip1(n8160), .ip2(n8100), .op(n8102) );
  nor2_1 U8676 ( .ip1(n8099), .ip2(n13766), .op(n8159) );
  or2_1 U8677 ( .ip1(n8159), .ip2(n8100), .op(n8101) );
  nand2_1 U8678 ( .ip1(n8102), .ip2(n8101), .op(n8157) );
  xor2_1 U8679 ( .ip1(n8104), .ip2(n8103), .op(n8156) );
  nand2_1 U8680 ( .ip1(m1Inputs[118]), .ip2(n12699), .op(n8105) );
  nand2_1 U8681 ( .ip1(m1Inputs[118]), .ip2(n11974), .op(n8174) );
  nor3_1 U8682 ( .ip1(n14339), .ip2(n13835), .ip3(n8174), .op(n8109) );
  or2_1 U8683 ( .ip1(n8105), .ip2(n8109), .op(n8108) );
  or2_1 U8684 ( .ip1(n8106), .ip2(n8109), .op(n8107) );
  nand2_1 U8685 ( .ip1(n8108), .ip2(n8107), .op(n8162) );
  or2_1 U8686 ( .ip1(n8162), .ip2(n8109), .op(n8111) );
  nor2_1 U8687 ( .ip1(n8177), .ip2(n13594), .op(n8161) );
  or2_1 U8688 ( .ip1(n8161), .ip2(n8109), .op(n8110) );
  nand2_1 U8689 ( .ip1(n8111), .ip2(n8110), .op(n8196) );
  xnor2_1 U8690 ( .ip1(n8113), .ip2(n8112), .op(n8195) );
  xnor2_1 U8691 ( .ip1(n8115), .ip2(n8114), .op(n8194) );
  inv_1 U8692 ( .ip(n8116), .op(n8301) );
  fulladder U8693 ( .a(n8119), .b(n8118), .ci(n8117), .co(n8116), .s(n8120) );
  inv_1 U8694 ( .ip(n8120), .op(n8305) );
  fulladder U8695 ( .a(n8123), .b(n8122), .ci(n8121), .co(n8062), .s(n8124) );
  inv_1 U8696 ( .ip(n8124), .op(n8186) );
  fulladder U8697 ( .a(n8127), .b(n8126), .ci(n8125), .co(n8117), .s(n8185) );
  fulladder U8698 ( .a(n8130), .b(n8129), .ci(n8128), .co(n8125), .s(n8193) );
  nand2_1 U8699 ( .ip1(n4619), .ip2(m1Inputs[120]), .op(n8132) );
  nor3_1 U8700 ( .ip1(n13709), .ip2(n14372), .ip3(n8131), .op(n8136) );
  or2_1 U8701 ( .ip1(n8132), .ip2(n8136), .op(n8135) );
  or2_1 U8702 ( .ip1(n8133), .ip2(n8136), .op(n8134) );
  nand2_1 U8703 ( .ip1(n8135), .ip2(n8134), .op(n8225) );
  or2_1 U8704 ( .ip1(n8225), .ip2(n8136), .op(n8139) );
  nand2_1 U8705 ( .ip1(column[114]), .ip2(n14768), .op(n8224) );
  inv_1 U8706 ( .ip(n8224), .op(n8137) );
  or2_1 U8707 ( .ip1(n8137), .ip2(n8136), .op(n8138) );
  nand2_1 U8708 ( .ip1(n8139), .ip2(n8138), .op(n8202) );
  nand2_1 U8709 ( .ip1(n13614), .ip2(m1Inputs[119]), .op(n8141) );
  nor3_1 U8710 ( .ip1(n13082), .ip2(n14433), .ip3(n8140), .op(n8146) );
  or2_1 U8711 ( .ip1(n8141), .ip2(n8146), .op(n8144) );
  or2_1 U8712 ( .ip1(n8142), .ip2(n8146), .op(n8143) );
  nand2_1 U8713 ( .ip1(n8144), .ip2(n8143), .op(n8245) );
  or2_1 U8714 ( .ip1(n8245), .ip2(n8146), .op(n8148) );
  nor2_1 U8715 ( .ip1(n8145), .ip2(n13594), .op(n8244) );
  or2_1 U8716 ( .ip1(n8244), .ip2(n8146), .op(n8147) );
  nand2_1 U8717 ( .ip1(n8148), .ip2(n8147), .op(n8201) );
  nand2_1 U8718 ( .ip1(m1Inputs[115]), .ip2(n14975), .op(n8200) );
  fulladder U8719 ( .a(n8151), .b(n8150), .ci(n8149), .co(n8130), .s(n8198) );
  nor2_1 U8720 ( .ip1(n8153), .ip2(n8152), .op(n8155) );
  xor2_1 U8721 ( .ip1(n8155), .ip2(n8154), .op(n8197) );
  fulladder U8722 ( .a(n8158), .b(n8157), .ci(n8156), .co(n8129), .s(n8233) );
  xor2_1 U8723 ( .ip1(n8160), .ip2(n8159), .op(n8242) );
  xor2_1 U8724 ( .ip1(n8162), .ip2(n8161), .op(n8241) );
  xor2_1 U8725 ( .ip1(n8164), .ip2(n8163), .op(n8240) );
  inv_1 U8726 ( .ip(n8165), .op(n8232) );
  nor3_1 U8727 ( .ip1(n8166), .ip2(n14384), .ip3(n8250), .op(n8204) );
  or2_1 U8728 ( .ip1(\STAGE_1/weightReg [7]), .ip2(n8167), .op(n8169) );
  or2_1 U8729 ( .ip1(m1Inputs[115]), .ip2(n8167), .op(n8168) );
  nand2_1 U8730 ( .ip1(n8169), .ip2(n8168), .op(n8203) );
  nand2_1 U8731 ( .ip1(m1Inputs[114]), .ip2(n14975), .op(n8205) );
  nor2_1 U8732 ( .ip1(n8203), .ip2(n8205), .op(n8170) );
  nor2_1 U8733 ( .ip1(n8204), .ip2(n8170), .op(n8239) );
  nand2_1 U8734 ( .ip1(n14369), .ip2(m1Inputs[117]), .op(n8173) );
  nor3_1 U8735 ( .ip1(n8172), .ip2(n13835), .ip3(n8171), .op(n8178) );
  or2_1 U8736 ( .ip1(n8173), .ip2(n8178), .op(n8176) );
  or2_1 U8737 ( .ip1(n8174), .ip2(n8178), .op(n8175) );
  nand2_1 U8738 ( .ip1(n8176), .ip2(n8175), .op(n8212) );
  or2_1 U8739 ( .ip1(n8212), .ip2(n8178), .op(n8180) );
  nor2_1 U8740 ( .ip1(n8177), .ip2(n12083), .op(n8211) );
  or2_1 U8741 ( .ip1(n8211), .ip2(n8178), .op(n8179) );
  nand2_1 U8742 ( .ip1(n8180), .ip2(n8179), .op(n8238) );
  xor2_1 U8743 ( .ip1(n8182), .ip2(n8181), .op(n8237) );
  inv_1 U8744 ( .ip(n8183), .op(n8304) );
  fulladder U8745 ( .a(n8186), .b(n8185), .ci(n8184), .co(n8183), .s(n8187) );
  inv_1 U8746 ( .ip(n8187), .op(n8308) );
  fulladder U8747 ( .a(n8190), .b(n8189), .ci(n8188), .co(n8126), .s(n8229) );
  fulladder U8748 ( .a(n8193), .b(n8192), .ci(n8191), .co(n8184), .s(n8228) );
  fulladder U8749 ( .a(n8196), .b(n8195), .ci(n8194), .co(n8128), .s(n8236) );
  fulladder U8750 ( .a(n8199), .b(n8198), .ci(n8197), .co(n8192), .s(n8235) );
  fulladder U8751 ( .a(n8202), .b(n8201), .ci(n8200), .co(n8199), .s(n8259) );
  nor2_1 U8752 ( .ip1(n8204), .ip2(n8203), .op(n8206) );
  xor2_1 U8753 ( .ip1(n8206), .ip2(n8205), .op(n8268) );
  nor2_1 U8754 ( .ip1(n8208), .ip2(n8207), .op(n8209) );
  nor2_1 U8755 ( .ip1(n8210), .ip2(n8209), .op(n8267) );
  xnor2_1 U8756 ( .ip1(n8212), .ip2(n8211), .op(n8266) );
  or2_1 U8757 ( .ip1(n8213), .ip2(n8214), .op(n8217) );
  or2_1 U8758 ( .ip1(n8215), .ip2(n8214), .op(n8216) );
  nand2_1 U8759 ( .ip1(n8217), .ip2(n8216), .op(n8265) );
  or2_1 U8760 ( .ip1(n8218), .ip2(n8220), .op(n8223) );
  inv_1 U8761 ( .ip(n8219), .op(n8221) );
  or2_1 U8762 ( .ip1(n8221), .ip2(n8220), .op(n8222) );
  nand2_1 U8763 ( .ip1(n8223), .ip2(n8222), .op(n8264) );
  xor2_1 U8764 ( .ip1(n8225), .ip2(n8224), .op(n8263) );
  inv_1 U8765 ( .ip(n8226), .op(n8307) );
  fulladder U8766 ( .a(n8229), .b(n8228), .ci(n8227), .co(n8226), .s(n8230) );
  inv_1 U8767 ( .ip(n8230), .op(n8311) );
  fulladder U8768 ( .a(n8233), .b(n8232), .ci(n8231), .co(n8191), .s(n8255) );
  fulladder U8769 ( .a(n8236), .b(n8235), .ci(n8234), .co(n8227), .s(n8254) );
  fulladder U8770 ( .a(n8239), .b(n8238), .ci(n8237), .co(n8231), .s(n8262) );
  fulladder U8771 ( .a(n8242), .b(n8241), .ci(n8240), .co(n8165), .s(n8243) );
  inv_1 U8772 ( .ip(n8243), .op(n8261) );
  xnor2_1 U8773 ( .ip1(n8245), .ip2(n8244), .op(n8279) );
  fulladder U8774 ( .a(n8248), .b(n8247), .ci(n8246), .co(n8278), .s(n7735) );
  fulladder U8775 ( .a(n8251), .b(n8250), .ci(n8249), .co(n8277), .s(n7720) );
  inv_1 U8776 ( .ip(n8252), .op(n8310) );
  fulladder U8777 ( .a(n8255), .b(n8254), .ci(n8253), .co(n8252), .s(n8256) );
  inv_1 U8778 ( .ip(n8256), .op(n8314) );
  fulladder U8779 ( .a(n8259), .b(n8258), .ci(n8257), .co(n8234), .s(n8275) );
  fulladder U8780 ( .a(n8262), .b(n8261), .ci(n8260), .co(n8253), .s(n8274) );
  fulladder U8781 ( .a(n8265), .b(n8264), .ci(n8263), .co(n8257), .s(n8283) );
  fulladder U8782 ( .a(n8268), .b(n8267), .ci(n8266), .co(n8258), .s(n8282) );
  fulladder U8783 ( .a(n8271), .b(n8270), .ci(n8269), .co(n8281), .s(n7714) );
  inv_1 U8784 ( .ip(n8272), .op(n8313) );
  fulladder U8785 ( .a(n8275), .b(n8274), .ci(n8273), .co(n8272), .s(n8276) );
  inv_1 U8786 ( .ip(n8276), .op(n8317) );
  fulladder U8787 ( .a(n8279), .b(n8278), .ci(n8277), .co(n8260), .s(n8280) );
  inv_1 U8788 ( .ip(n8280), .op(n8290) );
  fulladder U8789 ( .a(n8283), .b(n8282), .ci(n8281), .co(n8273), .s(n8284) );
  inv_1 U8790 ( .ip(n8284), .op(n8289) );
  fulladder U8791 ( .a(n8287), .b(n8286), .ci(n8285), .co(n8288), .s(n8295) );
  fulladder U8792 ( .a(n8290), .b(n8289), .ci(n8288), .co(n8316), .s(n8320) );
  fulladder U8793 ( .a(n8293), .b(n8292), .ci(n8291), .co(n8319), .s(
        \STAGE_1/M8/sum [1]) );
  fulladder U8794 ( .a(n8296), .b(n8295), .ci(n8294), .co(n8318), .s(n8293) );
  fulladder U8795 ( .a(n8299), .b(n8298), .ci(n8297), .co(n14336), .s(
        \STAGE_1/M8/sum [9]) );
  fulladder U8796 ( .a(n8302), .b(n8301), .ci(n8300), .co(n8297), .s(
        \STAGE_1/M8/sum [8]) );
  fulladder U8797 ( .a(n8305), .b(n8304), .ci(n8303), .co(n8300), .s(
        \STAGE_1/M8/sum [7]) );
  fulladder U8798 ( .a(n8308), .b(n8307), .ci(n8306), .co(n8303), .s(
        \STAGE_1/M8/sum [6]) );
  fulladder U8799 ( .a(n8311), .b(n8310), .ci(n8309), .co(n8306), .s(
        \STAGE_1/M8/sum [5]) );
  fulladder U8800 ( .a(n8314), .b(n8313), .ci(n8312), .co(n8309), .s(
        \STAGE_1/M8/sum [4]) );
  fulladder U8801 ( .a(n8317), .b(n8316), .ci(n8315), .co(n8312), .s(
        \STAGE_1/M8/sum [3]) );
  fulladder U8802 ( .a(n8320), .b(n8319), .ci(n8318), .co(n8315), .s(
        \STAGE_1/M8/sum [2]) );
  nand2_1 U8803 ( .ip1(m1Inputs[148]), .ip2(\STAGE_1/weightReg [5]), .op(n8322) );
  nor3_1 U8804 ( .ip1(n4624), .ip2(n14852), .ip3(n8321), .op(n8834) );
  or2_1 U8805 ( .ip1(n8322), .ip2(n8834), .op(n8324) );
  nand2_1 U8806 ( .ip1(n11974), .ip2(m1Inputs[149]), .op(n8792) );
  or2_1 U8807 ( .ip1(n8792), .ip2(n8834), .op(n8323) );
  nand2_1 U8808 ( .ip1(n8324), .ip2(n8323), .op(n8833) );
  nor2_1 U8809 ( .ip1(n8797), .ip2(n6503), .op(n8835) );
  xnor2_1 U8810 ( .ip1(n8833), .ip2(n8835), .op(n8891) );
  and3_1 U8811 ( .ip1(n12578), .ip2(m1Inputs[153]), .ip3(n8325), .op(n8830) );
  inv_1 U8812 ( .ip(m1Inputs[153]), .op(n14825) );
  nor2_1 U8813 ( .ip1(n10476), .ip2(n14825), .op(n8326) );
  or2_1 U8814 ( .ip1(m1Inputs[150]), .ip2(n8326), .op(n8328) );
  or2_1 U8815 ( .ip1(n9733), .ip2(n8326), .op(n8327) );
  nand2_1 U8816 ( .ip1(n8328), .ip2(n8327), .op(n8828) );
  nor2_1 U8817 ( .ip1(n8830), .ip2(n8828), .op(n8329) );
  nand2_1 U8818 ( .ip1(m1Inputs[144]), .ip2(n14994), .op(n8827) );
  xor2_1 U8819 ( .ip1(n8329), .ip2(n8827), .op(n8890) );
  fulladder U8820 ( .a(n8332), .b(n8331), .ci(n8330), .co(n8889), .s(n4768) );
  inv_1 U8821 ( .ip(n8333), .op(n8916) );
  inv_1 U8822 ( .ip(n8334), .op(n8338) );
  nor2_1 U8823 ( .ip1(n8336), .ip2(n8335), .op(n8337) );
  nor2_1 U8824 ( .ip1(n8338), .ip2(n8337), .op(n8871) );
  nand2_1 U8825 ( .ip1(m1Inputs[147]), .ip2(\STAGE_1/weightReg [6]), .op(n8870) );
  nand2_1 U8826 ( .ip1(m1Inputs[146]), .ip2(n14835), .op(n8869) );
  inv_1 U8827 ( .ip(n8339), .op(n8907) );
  or2_1 U8828 ( .ip1(n8340), .ip2(n8341), .op(n8344) );
  or2_1 U8829 ( .ip1(n8342), .ip2(n8341), .op(n8343) );
  nand2_1 U8830 ( .ip1(n8344), .ip2(n8343), .op(n8868) );
  or2_1 U8831 ( .ip1(n8345), .ip2(n8346), .op(n8349) );
  or2_1 U8832 ( .ip1(n8347), .ip2(n8346), .op(n8348) );
  nand2_1 U8833 ( .ip1(n8349), .ip2(n8348), .op(n8867) );
  nand2_1 U8834 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[151]), .op(n8351) );
  nor3_1 U8835 ( .ip1(n10555), .ip2(n14882), .ip3(n8350), .op(n8840) );
  or2_1 U8836 ( .ip1(n8351), .ip2(n8840), .op(n8353) );
  nand2_1 U8837 ( .ip1(n10507), .ip2(m1Inputs[152]), .op(n8753) );
  or2_1 U8838 ( .ip1(n8753), .ip2(n8840), .op(n8352) );
  nand2_1 U8839 ( .ip1(n8353), .ip2(n8352), .op(n8838) );
  nand2_1 U8840 ( .ip1(column[145]), .ip2(n13498), .op(n8839) );
  xor2_1 U8841 ( .ip1(n8838), .ip2(n8839), .op(n8866) );
  inv_1 U8842 ( .ip(n8354), .op(n8906) );
  fulladder U8843 ( .a(n8357), .b(n8356), .ci(n8355), .co(n8905), .s(n8361) );
  fulladder U8844 ( .a(n8360), .b(n8359), .ci(n8358), .co(n8914), .s(n8362) );
  fulladder U8845 ( .a(n8363), .b(n8362), .ci(n8361), .co(n8912), .s(n8366) );
  fulladder U8846 ( .a(n8366), .b(n8365), .ci(n8364), .co(n8911), .s(
        \STAGE_1/M10/sum [0]) );
  inv_1 U8847 ( .ip(m1Inputs[158]), .op(n14903) );
  nor2_1 U8848 ( .ip1(n14903), .ip2(n14783), .op(n14774) );
  inv_1 U8849 ( .ip(m1Inputs[155]), .op(n8709) );
  nor2_1 U8850 ( .ip1(n8709), .ip2(n14368), .op(n14773) );
  nand2_1 U8851 ( .ip1(n13614), .ip2(m1Inputs[159]), .op(n14772) );
  nor2_1 U8852 ( .ip1(n12083), .ip2(n14825), .op(n14761) );
  inv_1 U8853 ( .ip(m1Inputs[157]), .op(n14884) );
  nor2_1 U8854 ( .ip1(n14884), .ip2(n13835), .op(n14760) );
  nand2_1 U8855 ( .ip1(m1Inputs[147]), .ip2(\STAGE_1/weightReg [15]), .op(
        n14759) );
  nor2_1 U8856 ( .ip1(n14902), .ip2(n14852), .op(n8393) );
  nor2_1 U8857 ( .ip1(n13594), .ip2(n14841), .op(n8367) );
  or2_1 U8858 ( .ip1(m1Inputs[149]), .ip2(n8367), .op(n8369) );
  or2_1 U8859 ( .ip1(n14847), .ip2(n8367), .op(n8368) );
  nand2_1 U8860 ( .ip1(n8369), .ip2(n8368), .op(n8406) );
  nor3_1 U8861 ( .ip1(n8406), .ip2(n8408), .ip3(n14340), .op(n8370) );
  nor2_1 U8862 ( .ip1(n13594), .ip2(n14852), .op(n8506) );
  and3_1 U8863 ( .ip1(\STAGE_1/weightReg [11]), .ip2(m1Inputs[150]), .ip3(
        n8506), .op(n8407) );
  or2_1 U8864 ( .ip1(n8370), .ip2(n8407), .op(n8392) );
  nor2_1 U8865 ( .ip1(n13854), .ip2(n14903), .op(n8403) );
  nand2_1 U8866 ( .ip1(column[152]), .ip2(n13498), .op(n8402) );
  inv_1 U8867 ( .ip(m1Inputs[151]), .op(n14776) );
  nor2_1 U8868 ( .ip1(n12083), .ip2(n14776), .op(n8401) );
  nor2_1 U8869 ( .ip1(n14340), .ip2(n14852), .op(n14751) );
  nor2_1 U8870 ( .ip1(n14902), .ip2(n14841), .op(n14750) );
  nor2_1 U8871 ( .ip1(n13766), .ip2(n14882), .op(n8379) );
  and2_1 U8872 ( .ip1(column[153]), .ip2(n13498), .op(n8378) );
  inv_1 U8873 ( .ip(n8402), .op(n8377) );
  nor2_1 U8874 ( .ip1(n14825), .ip2(n14836), .op(n8394) );
  and3_1 U8875 ( .ip1(m1Inputs[154]), .ip2(n4627), .ip3(n8394), .op(n8374) );
  inv_1 U8876 ( .ip(m1Inputs[154]), .op(n14901) );
  nor2_1 U8877 ( .ip1(n14901), .ip2(n14836), .op(n8382) );
  or2_1 U8878 ( .ip1(\STAGE_1/weightReg [7]), .ip2(n8382), .op(n8372) );
  or2_1 U8879 ( .ip1(m1Inputs[153]), .ip2(n8382), .op(n8371) );
  nand2_1 U8880 ( .ip1(n8372), .ip2(n8371), .op(n8373) );
  nor2_1 U8881 ( .ip1(n8374), .ip2(n8373), .op(n8412) );
  or2_1 U8882 ( .ip1(n8412), .ip2(n8374), .op(n8376) );
  nor2_1 U8883 ( .ip1(n8709), .ip2(n8942), .op(n8411) );
  or2_1 U8884 ( .ip1(n8411), .ip2(n8374), .op(n8375) );
  nand2_1 U8885 ( .ip1(n8376), .ip2(n8375), .op(n8449) );
  nand2_1 U8886 ( .ip1(n13614), .ip2(m1Inputs[157]), .op(n8527) );
  inv_1 U8887 ( .ip(m1Inputs[159]), .op(n14837) );
  nor2_1 U8888 ( .ip1(n9047), .ip2(n14837), .op(n8455) );
  nand2_1 U8889 ( .ip1(m1Inputs[146]), .ip2(\STAGE_1/weightReg [14]), .op(
        n8454) );
  fulladder U8890 ( .a(n8379), .b(n8378), .ci(n8377), .co(n14749), .s(n8380)
         );
  inv_1 U8891 ( .ip(n8380), .op(n8447) );
  inv_1 U8892 ( .ip(n8381), .op(n14753) );
  nand2_1 U8893 ( .ip1(m1Inputs[155]), .ip2(\STAGE_1/weightReg [6]), .op(n8383) );
  and2_1 U8894 ( .ip1(n8382), .ip2(n14773), .op(n8415) );
  or2_1 U8895 ( .ip1(n8383), .ip2(n8415), .op(n8386) );
  nand2_1 U8896 ( .ip1(m1Inputs[154]), .ip2(n4627), .op(n8384) );
  or2_1 U8897 ( .ip1(n8384), .ip2(n8415), .op(n8385) );
  nand2_1 U8898 ( .ip1(n8386), .ip2(n8385), .op(n8414) );
  inv_1 U8899 ( .ip(m1Inputs[156]), .op(n8568) );
  nor2_1 U8900 ( .ip1(n8568), .ip2(n12746), .op(n8416) );
  xor2_1 U8901 ( .ip1(n8414), .ip2(n8416), .op(n8452) );
  nand2_1 U8902 ( .ip1(n13718), .ip2(m1Inputs[151]), .op(n14839) );
  nor3_1 U8903 ( .ip1(n13594), .ip2(n14841), .ip3(n14839), .op(n8426) );
  nor2_1 U8904 ( .ip1(n14824), .ip2(n14841), .op(n8387) );
  or2_1 U8905 ( .ip1(m1Inputs[151]), .ip2(n8387), .op(n8389) );
  or2_1 U8906 ( .ip1(n14876), .ip2(n8387), .op(n8388) );
  nand2_1 U8907 ( .ip1(n8389), .ip2(n8388), .op(n8390) );
  nor2_1 U8908 ( .ip1(n8426), .ip2(n8390), .op(n8425) );
  nor2_1 U8909 ( .ip1(n14340), .ip2(n14785), .op(n8427) );
  xor2_1 U8910 ( .ip1(n8425), .ip2(n8427), .op(n8451) );
  nor2_1 U8911 ( .ip1(n8568), .ip2(n14783), .op(n8458) );
  nor2_1 U8912 ( .ip1(n6503), .ip2(n14882), .op(n8457) );
  nand2_1 U8913 ( .ip1(m1Inputs[145]), .ip2(\STAGE_1/weightReg [15]), .op(
        n8456) );
  fulladder U8914 ( .a(n8393), .b(n8392), .ci(n8391), .co(n14755), .s(n8515)
         );
  nand2_1 U8915 ( .ip1(m1Inputs[153]), .ip2(n13637), .op(n8556) );
  nor3_1 U8916 ( .ip1(n8709), .ip2(n14836), .ip3(n8556), .op(n8398) );
  or2_1 U8917 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n8394), .op(n8396) );
  or2_1 U8918 ( .ip1(m1Inputs[155]), .ip2(n8394), .op(n8395) );
  nand2_1 U8919 ( .ip1(n8396), .ip2(n8395), .op(n8397) );
  nor2_1 U8920 ( .ip1(n8398), .ip2(n8397), .op(n8477) );
  or2_1 U8921 ( .ip1(n8477), .ip2(n8398), .op(n8400) );
  nor2_1 U8922 ( .ip1(n8797), .ip2(n14842), .op(n8476) );
  or2_1 U8923 ( .ip1(n8476), .ip2(n8398), .op(n8399) );
  nand2_1 U8924 ( .ip1(n8400), .ip2(n8399), .op(n8483) );
  nand2_1 U8925 ( .ip1(n9733), .ip2(m1Inputs[156]), .op(n8633) );
  nor2_1 U8926 ( .ip1(n10476), .ip2(n14837), .op(n8472) );
  nand2_1 U8927 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[150]), .op(n8471) );
  fulladder U8928 ( .a(n8403), .b(n8402), .ci(n8401), .co(n8391), .s(n8404) );
  inv_1 U8929 ( .ip(n8404), .op(n8481) );
  inv_1 U8930 ( .ip(n8405), .op(n8514) );
  nor2_1 U8931 ( .ip1(n8407), .ip2(n8406), .op(n8410) );
  nor2_1 U8932 ( .ip1(n8408), .ip2(n14373), .op(n8409) );
  xor2_1 U8933 ( .ip1(n8410), .ip2(n8409), .op(n8480) );
  xor2_1 U8934 ( .ip1(n8412), .ip2(n8411), .op(n8479) );
  nor2_1 U8935 ( .ip1(n14901), .ip2(n12746), .op(n8475) );
  nand2_1 U8936 ( .ip1(m1Inputs[144]), .ip2(\STAGE_1/weightReg [15]), .op(
        n8474) );
  inv_1 U8937 ( .ip(n8413), .op(n14806) );
  or2_1 U8938 ( .ip1(n8414), .ip2(n8415), .op(n8418) );
  or2_1 U8939 ( .ip1(n8416), .ip2(n8415), .op(n8417) );
  nand2_1 U8940 ( .ip1(n8418), .ip2(n8417), .op(n14747) );
  nand2_1 U8941 ( .ip1(m1Inputs[157]), .ip2(n13637), .op(n8432) );
  nor2_1 U8942 ( .ip1(n8721), .ip2(n14853), .op(n8431) );
  nand2_1 U8943 ( .ip1(n14838), .ip2(m1Inputs[153]), .op(n8430) );
  nand2_1 U8944 ( .ip1(m1Inputs[154]), .ip2(n14975), .op(n8420) );
  nand2_1 U8945 ( .ip1(m1Inputs[152]), .ip2(n14629), .op(n8419) );
  xor2_1 U8946 ( .ip1(n8420), .ip2(n8419), .op(n14736) );
  nand2_1 U8947 ( .ip1(column[154]), .ip2(n15042), .op(n8421) );
  xor2_1 U8948 ( .ip1(n14736), .ip2(n8421), .op(n14745) );
  nand2_1 U8949 ( .ip1(n14847), .ip2(m1Inputs[156]), .op(n15006) );
  nand2_1 U8950 ( .ip1(m1Inputs[151]), .ip2(n12981), .op(n8549) );
  nor2_1 U8951 ( .ip1(n15006), .ip2(n8549), .op(n14740) );
  or2_1 U8952 ( .ip1(n14839), .ip2(n14740), .op(n8424) );
  nand2_1 U8953 ( .ip1(m1Inputs[156]), .ip2(\STAGE_1/weightReg [6]), .op(n8422) );
  or2_1 U8954 ( .ip1(n8422), .ip2(n14740), .op(n8423) );
  nand2_1 U8955 ( .ip1(n8424), .ip2(n8423), .op(n14739) );
  nor2_1 U8956 ( .ip1(n14842), .ip2(n14785), .op(n14741) );
  xnor2_1 U8957 ( .ip1(n14739), .ip2(n14741), .op(n14790) );
  or2_1 U8958 ( .ip1(n8425), .ip2(n8426), .op(n8429) );
  or2_1 U8959 ( .ip1(n8427), .ip2(n8426), .op(n8428) );
  nand2_1 U8960 ( .ip1(n8429), .ip2(n8428), .op(n14789) );
  nor2_1 U8961 ( .ip1(n6745), .ip2(n14837), .op(n8434) );
  nand2_1 U8962 ( .ip1(n13614), .ip2(m1Inputs[158]), .op(n8501) );
  nand2_1 U8963 ( .ip1(m1Inputs[147]), .ip2(\STAGE_1/weightReg [14]), .op(
        n8433) );
  fulladder U8964 ( .a(n8432), .b(n8431), .ci(n8430), .co(n14746), .s(n8470)
         );
  fulladder U8965 ( .a(n8434), .b(n8501), .ci(n8433), .co(n14788), .s(n8469)
         );
  nor2_1 U8966 ( .ip1(n14776), .ip2(n14368), .op(n8493) );
  and2_1 U8967 ( .ip1(n8457), .ip2(n8493), .op(n8498) );
  nor2_1 U8968 ( .ip1(n14882), .ip2(n14384), .op(n8435) );
  or2_1 U8969 ( .ip1(m1Inputs[151]), .ip2(n8435), .op(n8437) );
  or2_1 U8970 ( .ip1(n14838), .ip2(n8435), .op(n8436) );
  nand2_1 U8971 ( .ip1(n8437), .ip2(n8436), .op(n8497) );
  inv_1 U8972 ( .ip(n14373), .op(n15028) );
  nand2_1 U8973 ( .ip1(m1Inputs[146]), .ip2(n15028), .op(n8499) );
  nor2_1 U8974 ( .ip1(n8497), .ip2(n8499), .op(n8438) );
  nor2_1 U8975 ( .ip1(n8498), .ip2(n8438), .op(n8488) );
  nand2_1 U8976 ( .ip1(n4672), .ip2(m1Inputs[157]), .op(n8439) );
  nand2_1 U8977 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[157]), .op(n8461) );
  nor3_1 U8978 ( .ip1(n10555), .ip2(n14903), .ip3(n8461), .op(n8443) );
  or2_1 U8979 ( .ip1(n8439), .ip2(n8443), .op(n8442) );
  nand2_1 U8980 ( .ip1(n13707), .ip2(m1Inputs[158]), .op(n8440) );
  or2_1 U8981 ( .ip1(n8440), .ip2(n8443), .op(n8441) );
  nand2_1 U8982 ( .ip1(n8442), .ip2(n8441), .op(n8512) );
  or2_1 U8983 ( .ip1(n8512), .ip2(n8443), .op(n8446) );
  nand2_1 U8984 ( .ip1(column[151]), .ip2(n13498), .op(n8511) );
  inv_1 U8985 ( .ip(n8511), .op(n8444) );
  or2_1 U8986 ( .ip1(n8444), .ip2(n8443), .op(n8445) );
  nand2_1 U8987 ( .ip1(n8446), .ip2(n8445), .op(n8487) );
  nand2_1 U8988 ( .ip1(n15025), .ip2(m1Inputs[148]), .op(n8486) );
  fulladder U8989 ( .a(n8449), .b(n8448), .ci(n8447), .co(n8381), .s(n8519) );
  fulladder U8990 ( .a(n8452), .b(n8451), .ci(n8450), .co(n14752), .s(n8453)
         );
  inv_1 U8991 ( .ip(n8453), .op(n8518) );
  fulladder U8992 ( .a(n8527), .b(n8455), .ci(n8454), .co(n8448), .s(n8522) );
  fulladder U8993 ( .a(n8458), .b(n8457), .ci(n8456), .co(n8450), .s(n8459) );
  inv_1 U8994 ( .ip(n8459), .op(n8521) );
  nand2_1 U8995 ( .ip1(n4619), .ip2(m1Inputs[156]), .op(n8460) );
  nand2_1 U8996 ( .ip1(n10507), .ip2(m1Inputs[156]), .op(n8570) );
  nor3_1 U8997 ( .ip1(n10555), .ip2(n14884), .ip3(n8570), .op(n8464) );
  or2_1 U8998 ( .ip1(n8460), .ip2(n8464), .op(n8463) );
  or2_1 U8999 ( .ip1(n8461), .ip2(n8464), .op(n8462) );
  nand2_1 U9000 ( .ip1(n8463), .ip2(n8462), .op(n8563) );
  or2_1 U9001 ( .ip1(n8563), .ip2(n8464), .op(n8467) );
  nand2_1 U9002 ( .ip1(column[150]), .ip2(n13498), .op(n8562) );
  inv_1 U9003 ( .ip(n8562), .op(n8465) );
  or2_1 U9004 ( .ip1(n8465), .ip2(n8464), .op(n8466) );
  nand2_1 U9005 ( .ip1(n8467), .ip2(n8466), .op(n8547) );
  nand2_1 U9006 ( .ip1(m1Inputs[147]), .ip2(\STAGE_1/weightReg [12]), .op(
        n8546) );
  nand2_1 U9007 ( .ip1(n14847), .ip2(m1Inputs[148]), .op(n8545) );
  fulladder U9008 ( .a(n8470), .b(n8469), .ci(n8468), .co(n14792), .s(n8580)
         );
  fulladder U9009 ( .a(n8633), .b(n8472), .ci(n8471), .co(n8482), .s(n8473) );
  inv_1 U9010 ( .ip(n8473), .op(n8593) );
  fulladder U9011 ( .a(n8475), .b(n8506), .ci(n8474), .co(n8478), .s(n8592) );
  xor2_1 U9012 ( .ip1(n8477), .ip2(n8476), .op(n8591) );
  fulladder U9013 ( .a(n8480), .b(n8479), .ci(n8478), .co(n8513), .s(n8588) );
  fulladder U9014 ( .a(n8483), .b(n8482), .ci(n8481), .co(n8405), .s(n8484) );
  inv_1 U9015 ( .ip(n8484), .op(n8587) );
  inv_1 U9016 ( .ip(n8485), .op(n8579) );
  fulladder U9017 ( .a(n8488), .b(n8487), .ci(n8486), .co(n8468), .s(n8586) );
  nor3_1 U9018 ( .ip1(n14901), .ip2(n4624), .ip3(n8556), .op(n8613) );
  nor2_1 U9019 ( .ip1(n14825), .ip2(n13835), .op(n8489) );
  or2_1 U9020 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n8489), .op(n8491) );
  or2_1 U9021 ( .ip1(m1Inputs[154]), .ip2(n8489), .op(n8490) );
  nand2_1 U9022 ( .ip1(n8491), .ip2(n8490), .op(n8612) );
  nand2_1 U9023 ( .ip1(n14838), .ip2(m1Inputs[150]), .op(n8614) );
  nor2_1 U9024 ( .ip1(n8612), .ip2(n8614), .op(n8492) );
  nor2_1 U9025 ( .ip1(n8613), .ip2(n8492), .op(n8541) );
  nor3_1 U9026 ( .ip1(n14882), .ip2(n14384), .ip3(n8549), .op(n8524) );
  or2_1 U9027 ( .ip1(n13749), .ip2(n8493), .op(n8495) );
  or2_1 U9028 ( .ip1(m1Inputs[152]), .ip2(n8493), .op(n8494) );
  nand2_1 U9029 ( .ip1(n8495), .ip2(n8494), .op(n8523) );
  nand2_1 U9030 ( .ip1(m1Inputs[145]), .ip2(n15028), .op(n8525) );
  nor2_1 U9031 ( .ip1(n8523), .ip2(n8525), .op(n8496) );
  nor2_1 U9032 ( .ip1(n8524), .ip2(n8496), .op(n8540) );
  nor2_1 U9033 ( .ip1(n8498), .ip2(n8497), .op(n8500) );
  xor2_1 U9034 ( .ip1(n8500), .ip2(n8499), .op(n8539) );
  nand2_1 U9035 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[155]), .op(n8711) );
  nor2_1 U9036 ( .ip1(n8711), .ip2(n8501), .op(n8617) );
  nor2_1 U9037 ( .ip1(n13082), .ip2(n8709), .op(n8502) );
  or2_1 U9038 ( .ip1(m1Inputs[158]), .ip2(n8502), .op(n8504) );
  or2_1 U9039 ( .ip1(n13803), .ip2(n8502), .op(n8503) );
  nand2_1 U9040 ( .ip1(n8504), .ip2(n8503), .op(n8616) );
  nand2_1 U9041 ( .ip1(m1Inputs[144]), .ip2(\STAGE_1/weightReg [14]), .op(
        n8618) );
  nor2_1 U9042 ( .ip1(n8616), .ip2(n8618), .op(n8505) );
  nor2_1 U9043 ( .ip1(n8617), .ip2(n8505), .op(n8544) );
  nor2_1 U9044 ( .ip1(n12083), .ip2(n14785), .op(n8564) );
  and2_1 U9045 ( .ip1(n8564), .ip2(n8506), .op(n8536) );
  nor2_1 U9046 ( .ip1(n13766), .ip2(n14852), .op(n8507) );
  or2_1 U9047 ( .ip1(m1Inputs[148]), .ip2(n8507), .op(n8509) );
  or2_1 U9048 ( .ip1(n14876), .ip2(n8507), .op(n8508) );
  nand2_1 U9049 ( .ip1(n8509), .ip2(n8508), .op(n8535) );
  nand2_1 U9050 ( .ip1(m1Inputs[146]), .ip2(\STAGE_1/weightReg [12]), .op(
        n8537) );
  nor2_1 U9051 ( .ip1(n8535), .ip2(n8537), .op(n8510) );
  nor2_1 U9052 ( .ip1(n8536), .ip2(n8510), .op(n8543) );
  xor2_1 U9053 ( .ip1(n8512), .ip2(n8511), .op(n8542) );
  fulladder U9054 ( .a(n8515), .b(n8514), .ci(n8513), .co(n14796), .s(n8516)
         );
  inv_1 U9055 ( .ip(n8516), .op(n8583) );
  fulladder U9056 ( .a(n8519), .b(n8518), .ci(n8517), .co(n14801), .s(n8582)
         );
  fulladder U9057 ( .a(n8522), .b(n8521), .ci(n8520), .co(n8517), .s(n8649) );
  nor2_1 U9058 ( .ip1(n8524), .ip2(n8523), .op(n8526) );
  xor2_1 U9059 ( .ip1(n8526), .ip2(n8525), .op(n8665) );
  nand2_1 U9060 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[154]), .op(n8764) );
  nor2_1 U9061 ( .ip1(n8764), .ip2(n8527), .op(n8532) );
  nor2_1 U9062 ( .ip1(n13082), .ip2(n14901), .op(n8528) );
  or2_1 U9063 ( .ip1(m1Inputs[157]), .ip2(n8528), .op(n8530) );
  or2_1 U9064 ( .ip1(n13803), .ip2(n8528), .op(n8529) );
  nand2_1 U9065 ( .ip1(n8530), .ip2(n8529), .op(n8531) );
  nor2_1 U9066 ( .ip1(n8532), .ip2(n8531), .op(n8672) );
  or2_1 U9067 ( .ip1(n8672), .ip2(n8532), .op(n8534) );
  nor2_1 U9068 ( .ip1(n8767), .ip2(n14340), .op(n8671) );
  or2_1 U9069 ( .ip1(n8671), .ip2(n8532), .op(n8533) );
  nand2_1 U9070 ( .ip1(n8534), .ip2(n8533), .op(n8664) );
  nor2_1 U9071 ( .ip1(n8536), .ip2(n8535), .op(n8538) );
  xor2_1 U9072 ( .ip1(n8538), .ip2(n8537), .op(n8663) );
  fulladder U9073 ( .a(n8541), .b(n8540), .ci(n8539), .co(n8585), .s(n8660) );
  fulladder U9074 ( .a(n8544), .b(n8543), .ci(n8542), .co(n8584), .s(n8659) );
  fulladder U9075 ( .a(n8547), .b(n8546), .ci(n8545), .co(n8520), .s(n8657) );
  nand2_1 U9076 ( .ip1(m1Inputs[150]), .ip2(n14835), .op(n8548) );
  nand2_1 U9077 ( .ip1(m1Inputs[150]), .ip2(\STAGE_1/weightReg [6]), .op(n8604) );
  nor3_1 U9078 ( .ip1(n14776), .ip2(n14368), .ip3(n8604), .op(n8552) );
  or2_1 U9079 ( .ip1(n8548), .ip2(n8552), .op(n8551) );
  or2_1 U9080 ( .ip1(n8549), .ip2(n8552), .op(n8550) );
  nand2_1 U9081 ( .ip1(n8551), .ip2(n8550), .op(n8676) );
  or2_1 U9082 ( .ip1(n8676), .ip2(n8552), .op(n8554) );
  nor2_1 U9083 ( .ip1(n8721), .ip2(n14824), .op(n8675) );
  or2_1 U9084 ( .ip1(n8675), .ip2(n8552), .op(n8553) );
  nand2_1 U9085 ( .ip1(n8554), .ip2(n8553), .op(n8625) );
  nand2_1 U9086 ( .ip1(m1Inputs[152]), .ip2(\STAGE_1/weightReg [5]), .op(n8555) );
  nand2_1 U9087 ( .ip1(m1Inputs[152]), .ip2(n13637), .op(n8627) );
  nor3_1 U9088 ( .ip1(n14825), .ip2(n4624), .ip3(n8627), .op(n8559) );
  or2_1 U9089 ( .ip1(n8555), .ip2(n8559), .op(n8558) );
  or2_1 U9090 ( .ip1(n8556), .ip2(n8559), .op(n8557) );
  nand2_1 U9091 ( .ip1(n8558), .ip2(n8557), .op(n8674) );
  or2_1 U9092 ( .ip1(n8674), .ip2(n8559), .op(n8561) );
  nor2_1 U9093 ( .ip1(n8797), .ip2(n14188), .op(n8673) );
  or2_1 U9094 ( .ip1(n8673), .ip2(n8559), .op(n8560) );
  nand2_1 U9095 ( .ip1(n8561), .ip2(n8560), .op(n8624) );
  xor2_1 U9096 ( .ip1(n8563), .ip2(n8562), .op(n8623) );
  nand2_1 U9097 ( .ip1(n14838), .ip2(m1Inputs[148]), .op(n8773) );
  nor3_1 U9098 ( .ip1(n12083), .ip2(n14852), .ip3(n8773), .op(n8639) );
  or2_1 U9099 ( .ip1(m1Inputs[149]), .ip2(n8564), .op(n8566) );
  or2_1 U9100 ( .ip1(n14838), .ip2(n8564), .op(n8565) );
  nand2_1 U9101 ( .ip1(n8566), .ip2(n8565), .op(n8638) );
  nand2_1 U9102 ( .ip1(m1Inputs[147]), .ip2(\STAGE_1/weightReg [10]), .op(
        n8640) );
  nor2_1 U9103 ( .ip1(n8638), .ip2(n8640), .op(n8567) );
  nor2_1 U9104 ( .ip1(n8639), .ip2(n8567), .op(n8622) );
  nand2_1 U9105 ( .ip1(n4672), .ip2(m1Inputs[155]), .op(n8569) );
  nand2_1 U9106 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[155]), .op(n8596) );
  nor3_1 U9107 ( .ip1(n10555), .ip2(n8568), .ip3(n8596), .op(n8573) );
  or2_1 U9108 ( .ip1(n8569), .ip2(n8573), .op(n8572) );
  or2_1 U9109 ( .ip1(n8570), .ip2(n8573), .op(n8571) );
  nand2_1 U9110 ( .ip1(n8572), .ip2(n8571), .op(n8611) );
  or2_1 U9111 ( .ip1(n8611), .ip2(n8573), .op(n8576) );
  nand2_1 U9112 ( .ip1(column[149]), .ip2(n13498), .op(n8610) );
  inv_1 U9113 ( .ip(n8610), .op(n8574) );
  or2_1 U9114 ( .ip1(n8574), .ip2(n8573), .op(n8575) );
  nand2_1 U9115 ( .ip1(n8576), .ip2(n8575), .op(n8621) );
  nand2_1 U9116 ( .ip1(m1Inputs[147]), .ip2(\STAGE_1/weightReg [11]), .op(
        n8620) );
  inv_1 U9117 ( .ip(n8577), .op(n14810) );
  fulladder U9118 ( .a(n8580), .b(n8579), .ci(n8578), .co(n14800), .s(n8645)
         );
  fulladder U9119 ( .a(n8583), .b(n8582), .ci(n8581), .co(n14804), .s(n8644)
         );
  fulladder U9120 ( .a(n8586), .b(n8585), .ci(n8584), .co(n8578), .s(n8653) );
  fulladder U9121 ( .a(n8589), .b(n8588), .ci(n8587), .co(n8485), .s(n8590) );
  inv_1 U9122 ( .ip(n8590), .op(n8652) );
  fulladder U9123 ( .a(n8593), .b(n8592), .ci(n8591), .co(n8589), .s(n8594) );
  inv_1 U9124 ( .ip(n8594), .op(n8682) );
  nand2_1 U9125 ( .ip1(n4619), .ip2(m1Inputs[154]), .op(n8595) );
  nand2_1 U9126 ( .ip1(n10507), .ip2(m1Inputs[154]), .op(n8701) );
  nor3_1 U9127 ( .ip1(n10555), .ip2(n8709), .ip3(n8701), .op(n8599) );
  or2_1 U9128 ( .ip1(n8595), .ip2(n8599), .op(n8598) );
  or2_1 U9129 ( .ip1(n8596), .ip2(n8599), .op(n8597) );
  nand2_1 U9130 ( .ip1(n8598), .ip2(n8597), .op(n8726) );
  or2_1 U9131 ( .ip1(n8726), .ip2(n8599), .op(n8602) );
  nand2_1 U9132 ( .ip1(column[148]), .ip2(n14768), .op(n8725) );
  inv_1 U9133 ( .ip(n8725), .op(n8600) );
  or2_1 U9134 ( .ip1(n8600), .ip2(n8599), .op(n8601) );
  nand2_1 U9135 ( .ip1(n8602), .ip2(n8601), .op(n8699) );
  nand2_1 U9136 ( .ip1(n4627), .ip2(m1Inputs[149]), .op(n8603) );
  nand2_1 U9137 ( .ip1(n13749), .ip2(m1Inputs[149]), .op(n8718) );
  nor3_1 U9138 ( .ip1(n14841), .ip2(n14384), .ip3(n8718), .op(n8607) );
  or2_1 U9139 ( .ip1(n8603), .ip2(n8607), .op(n8606) );
  or2_1 U9140 ( .ip1(n8604), .ip2(n8607), .op(n8605) );
  nand2_1 U9141 ( .ip1(n8606), .ip2(n8605), .op(n8737) );
  or2_1 U9142 ( .ip1(n8737), .ip2(n8607), .op(n8609) );
  nor2_1 U9143 ( .ip1(n8721), .ip2(n13594), .op(n8736) );
  or2_1 U9144 ( .ip1(n8736), .ip2(n8607), .op(n8608) );
  nand2_1 U9145 ( .ip1(n8609), .ip2(n8608), .op(n8698) );
  xor2_1 U9146 ( .ip1(n8611), .ip2(n8610), .op(n8697) );
  nor2_1 U9147 ( .ip1(n8613), .ip2(n8612), .op(n8615) );
  xor2_1 U9148 ( .ip1(n8615), .ip2(n8614), .op(n8668) );
  nor2_1 U9149 ( .ip1(n8617), .ip2(n8616), .op(n8619) );
  xor2_1 U9150 ( .ip1(n8619), .ip2(n8618), .op(n8667) );
  fulladder U9151 ( .a(n8622), .b(n8621), .ci(n8620), .co(n8655), .s(n8689) );
  fulladder U9152 ( .a(n8625), .b(n8624), .ci(n8623), .co(n8656), .s(n8688) );
  nand2_1 U9153 ( .ip1(m1Inputs[151]), .ip2(\STAGE_1/weightReg [5]), .op(n8626) );
  nand2_1 U9154 ( .ip1(m1Inputs[151]), .ip2(n13637), .op(n8728) );
  nor3_1 U9155 ( .ip1(n14882), .ip2(n4624), .ip3(n8728), .op(n8630) );
  or2_1 U9156 ( .ip1(n8626), .ip2(n8630), .op(n8629) );
  or2_1 U9157 ( .ip1(n8627), .ip2(n8630), .op(n8628) );
  nand2_1 U9158 ( .ip1(n8629), .ip2(n8628), .op(n8735) );
  or2_1 U9159 ( .ip1(n8735), .ip2(n8630), .op(n8632) );
  nor2_1 U9160 ( .ip1(n8797), .ip2(n14824), .op(n8734) );
  or2_1 U9161 ( .ip1(n8734), .ip2(n8630), .op(n8631) );
  nand2_1 U9162 ( .ip1(n8632), .ip2(n8631), .op(n8692) );
  nor3_1 U9163 ( .ip1(n10476), .ip2(n14825), .ip3(n8633), .op(n8775) );
  nor2_1 U9164 ( .ip1(n13487), .ip2(n14825), .op(n8634) );
  or2_1 U9165 ( .ip1(m1Inputs[156]), .ip2(n8634), .op(n8636) );
  or2_1 U9166 ( .ip1(n13803), .ip2(n8634), .op(n8635) );
  nand2_1 U9167 ( .ip1(n8636), .ip2(n8635), .op(n8774) );
  nand2_1 U9168 ( .ip1(m1Inputs[144]), .ip2(\STAGE_1/weightReg [12]), .op(
        n8776) );
  nor2_1 U9169 ( .ip1(n8774), .ip2(n8776), .op(n8637) );
  nor2_1 U9170 ( .ip1(n8775), .ip2(n8637), .op(n8691) );
  nor2_1 U9171 ( .ip1(n8639), .ip2(n8638), .op(n8641) );
  xor2_1 U9172 ( .ip1(n8641), .ip2(n8640), .op(n8690) );
  inv_1 U9173 ( .ip(n8642), .op(n14809) );
  fulladder U9174 ( .a(n8645), .b(n8644), .ci(n8643), .co(n8642), .s(n8646) );
  inv_1 U9175 ( .ip(n8646), .op(n8919) );
  fulladder U9176 ( .a(n8649), .b(n8648), .ci(n8647), .co(n8581), .s(n8650) );
  inv_1 U9177 ( .ip(n8650), .op(n8679) );
  fulladder U9178 ( .a(n8653), .b(n8652), .ci(n8651), .co(n8643), .s(n8654) );
  inv_1 U9179 ( .ip(n8654), .op(n8678) );
  fulladder U9180 ( .a(n8657), .b(n8656), .ci(n8655), .co(n8647), .s(n8658) );
  inv_1 U9181 ( .ip(n8658), .op(n8685) );
  fulladder U9182 ( .a(n8661), .b(n8660), .ci(n8659), .co(n8648), .s(n8662) );
  inv_1 U9183 ( .ip(n8662), .op(n8684) );
  fulladder U9184 ( .a(n8665), .b(n8664), .ci(n8663), .co(n8661), .s(n8666) );
  inv_1 U9185 ( .ip(n8666), .op(n8745) );
  fulladder U9186 ( .a(n8669), .b(n8668), .ci(n8667), .co(n8681), .s(n8670) );
  inv_1 U9187 ( .ip(n8670), .op(n8744) );
  xor2_1 U9188 ( .ip1(n8672), .ip2(n8671), .op(n8695) );
  xor2_1 U9189 ( .ip1(n8674), .ip2(n8673), .op(n8694) );
  xor2_1 U9190 ( .ip1(n8676), .ip2(n8675), .op(n8693) );
  fulladder U9191 ( .a(n8679), .b(n8678), .ci(n8677), .co(n8918), .s(n8922) );
  fulladder U9192 ( .a(n8682), .b(n8681), .ci(n8680), .co(n8651), .s(n8741) );
  fulladder U9193 ( .a(n8685), .b(n8684), .ci(n8683), .co(n8677), .s(n8686) );
  inv_1 U9194 ( .ip(n8686), .op(n8740) );
  fulladder U9195 ( .a(n8689), .b(n8688), .ci(n8687), .co(n8680), .s(n8749) );
  fulladder U9196 ( .a(n8692), .b(n8691), .ci(n8690), .co(n8687), .s(n8810) );
  fulladder U9197 ( .a(n8695), .b(n8694), .ci(n8693), .co(n8743), .s(n8696) );
  inv_1 U9198 ( .ip(n8696), .op(n8809) );
  fulladder U9199 ( .a(n8699), .b(n8698), .ci(n8697), .co(n8669), .s(n8808) );
  nand2_1 U9200 ( .ip1(n4672), .ip2(m1Inputs[153]), .op(n8700) );
  nand2_1 U9201 ( .ip1(n10507), .ip2(m1Inputs[153]), .op(n8755) );
  nor3_1 U9202 ( .ip1(n10555), .ip2(n14901), .ip3(n8755), .op(n8704) );
  or2_1 U9203 ( .ip1(n8700), .ip2(n8704), .op(n8703) );
  or2_1 U9204 ( .ip1(n8701), .ip2(n8704), .op(n8702) );
  nand2_1 U9205 ( .ip1(n8703), .ip2(n8702), .op(n8802) );
  or2_1 U9206 ( .ip1(n8802), .ip2(n8704), .op(n8707) );
  nand2_1 U9207 ( .ip1(column[147]), .ip2(n13498), .op(n8801) );
  inv_1 U9208 ( .ip(n8801), .op(n8705) );
  or2_1 U9209 ( .ip1(n8705), .ip2(n8704), .op(n8706) );
  nand2_1 U9210 ( .ip1(n8707), .ip2(n8706), .op(n8772) );
  nand2_1 U9211 ( .ip1(m1Inputs[147]), .ip2(n14994), .op(n8771) );
  nand2_1 U9212 ( .ip1(n13614), .ip2(m1Inputs[152]), .op(n8710) );
  nor3_1 U9213 ( .ip1(n13801), .ip2(n8709), .ip3(n8708), .op(n8714) );
  or2_1 U9214 ( .ip1(n8710), .ip2(n8714), .op(n8713) );
  or2_1 U9215 ( .ip1(n8711), .ip2(n8714), .op(n8712) );
  nand2_1 U9216 ( .ip1(n8713), .ip2(n8712), .op(n8786) );
  or2_1 U9217 ( .ip1(n8786), .ip2(n8714), .op(n8716) );
  nor2_1 U9218 ( .ip1(n8767), .ip2(n13579), .op(n8785) );
  or2_1 U9219 ( .ip1(n8785), .ip2(n8714), .op(n8715) );
  nand2_1 U9220 ( .ip1(n8716), .ip2(n8715), .op(n8780) );
  nand2_1 U9221 ( .ip1(m1Inputs[148]), .ip2(n14835), .op(n8717) );
  nor2_1 U9222 ( .ip1(n14785), .ip2(n14836), .op(n8788) );
  and3_1 U9223 ( .ip1(n4627), .ip2(m1Inputs[149]), .ip3(n8788), .op(n8722) );
  or2_1 U9224 ( .ip1(n8717), .ip2(n8722), .op(n8720) );
  or2_1 U9225 ( .ip1(n8718), .ip2(n8722), .op(n8719) );
  nand2_1 U9226 ( .ip1(n8720), .ip2(n8719), .op(n8782) );
  or2_1 U9227 ( .ip1(n8782), .ip2(n8722), .op(n8724) );
  nor2_1 U9228 ( .ip1(n8721), .ip2(n12083), .op(n8781) );
  or2_1 U9229 ( .ip1(n8781), .ip2(n8722), .op(n8723) );
  nand2_1 U9230 ( .ip1(n8724), .ip2(n8723), .op(n8779) );
  xor2_1 U9231 ( .ip1(n8726), .ip2(n8725), .op(n8778) );
  nand2_1 U9232 ( .ip1(m1Inputs[150]), .ip2(\STAGE_1/weightReg [5]), .op(n8727) );
  nand2_1 U9233 ( .ip1(m1Inputs[150]), .ip2(n13637), .op(n8794) );
  nor3_1 U9234 ( .ip1(n14776), .ip2(n13835), .ip3(n8794), .op(n8731) );
  or2_1 U9235 ( .ip1(n8727), .ip2(n8731), .op(n8730) );
  or2_1 U9236 ( .ip1(n8728), .ip2(n8731), .op(n8729) );
  nand2_1 U9237 ( .ip1(n8730), .ip2(n8729), .op(n8784) );
  or2_1 U9238 ( .ip1(n8784), .ip2(n8731), .op(n8733) );
  nor2_1 U9239 ( .ip1(n8797), .ip2(n13594), .op(n8783) );
  or2_1 U9240 ( .ip1(n8783), .ip2(n8731), .op(n8732) );
  nand2_1 U9241 ( .ip1(n8733), .ip2(n8732), .op(n8816) );
  xnor2_1 U9242 ( .ip1(n8735), .ip2(n8734), .op(n8815) );
  xnor2_1 U9243 ( .ip1(n8737), .ip2(n8736), .op(n8814) );
  inv_1 U9244 ( .ip(n8738), .op(n8921) );
  fulladder U9245 ( .a(n8741), .b(n8740), .ci(n8739), .co(n8738), .s(n8742) );
  inv_1 U9246 ( .ip(n8742), .op(n8925) );
  fulladder U9247 ( .a(n8745), .b(n8744), .ci(n8743), .co(n8683), .s(n8746) );
  inv_1 U9248 ( .ip(n8746), .op(n8806) );
  fulladder U9249 ( .a(n8749), .b(n8748), .ci(n8747), .co(n8739), .s(n8805) );
  fulladder U9250 ( .a(n8752), .b(n8751), .ci(n8750), .co(n8747), .s(n8813) );
  nand2_1 U9251 ( .ip1(n4672), .ip2(m1Inputs[152]), .op(n8754) );
  nor3_1 U9252 ( .ip1(n10555), .ip2(n14825), .ip3(n8753), .op(n8758) );
  or2_1 U9253 ( .ip1(n8754), .ip2(n8758), .op(n8757) );
  or2_1 U9254 ( .ip1(n8755), .ip2(n8758), .op(n8756) );
  nand2_1 U9255 ( .ip1(n8757), .ip2(n8756), .op(n8845) );
  or2_1 U9256 ( .ip1(n8845), .ip2(n8758), .op(n8761) );
  nand2_1 U9257 ( .ip1(column[146]), .ip2(n13498), .op(n8844) );
  inv_1 U9258 ( .ip(n8844), .op(n8759) );
  or2_1 U9259 ( .ip1(n8759), .ip2(n8758), .op(n8760) );
  nand2_1 U9260 ( .ip1(n8761), .ip2(n8760), .op(n8822) );
  nand2_1 U9261 ( .ip1(n9733), .ip2(m1Inputs[151]), .op(n8763) );
  nor3_1 U9262 ( .ip1(n13487), .ip2(n14901), .ip3(n8762), .op(n8768) );
  or2_1 U9263 ( .ip1(n8763), .ip2(n8768), .op(n8766) );
  or2_1 U9264 ( .ip1(n8764), .ip2(n8768), .op(n8765) );
  nand2_1 U9265 ( .ip1(n8766), .ip2(n8765), .op(n8865) );
  or2_1 U9266 ( .ip1(n8865), .ip2(n8768), .op(n8770) );
  nor2_1 U9267 ( .ip1(n8767), .ip2(n13594), .op(n8864) );
  or2_1 U9268 ( .ip1(n8864), .ip2(n8768), .op(n8769) );
  nand2_1 U9269 ( .ip1(n8770), .ip2(n8769), .op(n8821) );
  nand2_1 U9270 ( .ip1(m1Inputs[147]), .ip2(n14975), .op(n8820) );
  fulladder U9271 ( .a(n8773), .b(n8772), .ci(n8771), .co(n8752), .s(n8818) );
  nor2_1 U9272 ( .ip1(n8775), .ip2(n8774), .op(n8777) );
  xor2_1 U9273 ( .ip1(n8777), .ip2(n8776), .op(n8817) );
  fulladder U9274 ( .a(n8780), .b(n8779), .ci(n8778), .co(n8751), .s(n8853) );
  xor2_1 U9275 ( .ip1(n8782), .ip2(n8781), .op(n8862) );
  xor2_1 U9276 ( .ip1(n8784), .ip2(n8783), .op(n8861) );
  xor2_1 U9277 ( .ip1(n8786), .ip2(n8785), .op(n8860) );
  inv_1 U9278 ( .ip(n8787), .op(n8852) );
  nor3_1 U9279 ( .ip1(n14785), .ip2(n14368), .ip3(n8870), .op(n8824) );
  or2_1 U9280 ( .ip1(\STAGE_1/weightReg [7]), .ip2(n8788), .op(n8790) );
  or2_1 U9281 ( .ip1(m1Inputs[147]), .ip2(n8788), .op(n8789) );
  nand2_1 U9282 ( .ip1(n8790), .ip2(n8789), .op(n8823) );
  nand2_1 U9283 ( .ip1(m1Inputs[146]), .ip2(n14975), .op(n8825) );
  nor2_1 U9284 ( .ip1(n8823), .ip2(n8825), .op(n8791) );
  nor2_1 U9285 ( .ip1(n8824), .ip2(n8791), .op(n8859) );
  nand2_1 U9286 ( .ip1(n14369), .ip2(m1Inputs[149]), .op(n8793) );
  nor3_1 U9287 ( .ip1(n14841), .ip2(n4624), .ip3(n8792), .op(n8798) );
  or2_1 U9288 ( .ip1(n8793), .ip2(n8798), .op(n8796) );
  or2_1 U9289 ( .ip1(n8794), .ip2(n8798), .op(n8795) );
  nand2_1 U9290 ( .ip1(n8796), .ip2(n8795), .op(n8832) );
  or2_1 U9291 ( .ip1(n8832), .ip2(n8798), .op(n8800) );
  nor2_1 U9292 ( .ip1(n8797), .ip2(n12083), .op(n8831) );
  or2_1 U9293 ( .ip1(n8831), .ip2(n8798), .op(n8799) );
  nand2_1 U9294 ( .ip1(n8800), .ip2(n8799), .op(n8858) );
  xor2_1 U9295 ( .ip1(n8802), .ip2(n8801), .op(n8857) );
  inv_1 U9296 ( .ip(n8803), .op(n8924) );
  fulladder U9297 ( .a(n8806), .b(n8805), .ci(n8804), .co(n8803), .s(n8807) );
  inv_1 U9298 ( .ip(n8807), .op(n8928) );
  fulladder U9299 ( .a(n8810), .b(n8809), .ci(n8808), .co(n8748), .s(n8849) );
  fulladder U9300 ( .a(n8813), .b(n8812), .ci(n8811), .co(n8804), .s(n8848) );
  fulladder U9301 ( .a(n8816), .b(n8815), .ci(n8814), .co(n8750), .s(n8856) );
  fulladder U9302 ( .a(n8819), .b(n8818), .ci(n8817), .co(n8812), .s(n8855) );
  fulladder U9303 ( .a(n8822), .b(n8821), .ci(n8820), .co(n8819), .s(n8879) );
  nor2_1 U9304 ( .ip1(n8824), .ip2(n8823), .op(n8826) );
  xor2_1 U9305 ( .ip1(n8826), .ip2(n8825), .op(n8888) );
  nor2_1 U9306 ( .ip1(n8828), .ip2(n8827), .op(n8829) );
  nor2_1 U9307 ( .ip1(n8830), .ip2(n8829), .op(n8887) );
  xnor2_1 U9308 ( .ip1(n8832), .ip2(n8831), .op(n8886) );
  or2_1 U9309 ( .ip1(n8833), .ip2(n8834), .op(n8837) );
  or2_1 U9310 ( .ip1(n8835), .ip2(n8834), .op(n8836) );
  nand2_1 U9311 ( .ip1(n8837), .ip2(n8836), .op(n8885) );
  or2_1 U9312 ( .ip1(n8838), .ip2(n8840), .op(n8843) );
  inv_1 U9313 ( .ip(n8839), .op(n8841) );
  or2_1 U9314 ( .ip1(n8841), .ip2(n8840), .op(n8842) );
  nand2_1 U9315 ( .ip1(n8843), .ip2(n8842), .op(n8884) );
  xor2_1 U9316 ( .ip1(n8845), .ip2(n8844), .op(n8883) );
  inv_1 U9317 ( .ip(n8846), .op(n8927) );
  fulladder U9318 ( .a(n8849), .b(n8848), .ci(n8847), .co(n8846), .s(n8850) );
  inv_1 U9319 ( .ip(n8850), .op(n8931) );
  fulladder U9320 ( .a(n8853), .b(n8852), .ci(n8851), .co(n8811), .s(n8875) );
  fulladder U9321 ( .a(n8856), .b(n8855), .ci(n8854), .co(n8847), .s(n8874) );
  fulladder U9322 ( .a(n8859), .b(n8858), .ci(n8857), .co(n8851), .s(n8882) );
  fulladder U9323 ( .a(n8862), .b(n8861), .ci(n8860), .co(n8787), .s(n8863) );
  inv_1 U9324 ( .ip(n8863), .op(n8881) );
  xnor2_1 U9325 ( .ip1(n8865), .ip2(n8864), .op(n8899) );
  fulladder U9326 ( .a(n8868), .b(n8867), .ci(n8866), .co(n8898), .s(n8354) );
  fulladder U9327 ( .a(n8871), .b(n8870), .ci(n8869), .co(n8897), .s(n8339) );
  inv_1 U9328 ( .ip(n8872), .op(n8930) );
  fulladder U9329 ( .a(n8875), .b(n8874), .ci(n8873), .co(n8872), .s(n8876) );
  inv_1 U9330 ( .ip(n8876), .op(n8934) );
  fulladder U9331 ( .a(n8879), .b(n8878), .ci(n8877), .co(n8854), .s(n8895) );
  fulladder U9332 ( .a(n8882), .b(n8881), .ci(n8880), .co(n8873), .s(n8894) );
  fulladder U9333 ( .a(n8885), .b(n8884), .ci(n8883), .co(n8877), .s(n8903) );
  fulladder U9334 ( .a(n8888), .b(n8887), .ci(n8886), .co(n8878), .s(n8902) );
  fulladder U9335 ( .a(n8891), .b(n8890), .ci(n8889), .co(n8901), .s(n8333) );
  inv_1 U9336 ( .ip(n8892), .op(n8933) );
  fulladder U9337 ( .a(n8895), .b(n8894), .ci(n8893), .co(n8892), .s(n8896) );
  inv_1 U9338 ( .ip(n8896), .op(n8937) );
  fulladder U9339 ( .a(n8899), .b(n8898), .ci(n8897), .co(n8880), .s(n8900) );
  inv_1 U9340 ( .ip(n8900), .op(n8910) );
  fulladder U9341 ( .a(n8903), .b(n8902), .ci(n8901), .co(n8893), .s(n8904) );
  inv_1 U9342 ( .ip(n8904), .op(n8909) );
  fulladder U9343 ( .a(n8907), .b(n8906), .ci(n8905), .co(n8908), .s(n8915) );
  fulladder U9344 ( .a(n8910), .b(n8909), .ci(n8908), .co(n8936), .s(n8940) );
  fulladder U9345 ( .a(n8913), .b(n8912), .ci(n8911), .co(n8939), .s(
        \STAGE_1/M10/sum [1]) );
  fulladder U9346 ( .a(n8916), .b(n8915), .ci(n8914), .co(n8938), .s(n8913) );
  fulladder U9347 ( .a(n8919), .b(n8918), .ci(n8917), .co(n14808), .s(
        \STAGE_1/M10/sum [9]) );
  fulladder U9348 ( .a(n8922), .b(n8921), .ci(n8920), .co(n8917), .s(
        \STAGE_1/M10/sum [8]) );
  fulladder U9349 ( .a(n8925), .b(n8924), .ci(n8923), .co(n8920), .s(
        \STAGE_1/M10/sum [7]) );
  fulladder U9350 ( .a(n8928), .b(n8927), .ci(n8926), .co(n8923), .s(
        \STAGE_1/M10/sum [6]) );
  fulladder U9351 ( .a(n8931), .b(n8930), .ci(n8929), .co(n8926), .s(
        \STAGE_1/M10/sum [5]) );
  fulladder U9352 ( .a(n8934), .b(n8933), .ci(n8932), .co(n8929), .s(
        \STAGE_1/M10/sum [4]) );
  fulladder U9353 ( .a(n8937), .b(n8936), .ci(n8935), .co(n8932), .s(
        \STAGE_1/M10/sum [3]) );
  fulladder U9354 ( .a(n8940), .b(n8939), .ci(n8938), .co(n8935), .s(
        \STAGE_1/M10/sum [2]) );
  nand2_1 U9355 ( .ip1(m1Inputs[132]), .ip2(\STAGE_1/weightReg [5]), .op(n8943) );
  nor3_1 U9356 ( .ip1(n8942), .ip2(n9299), .ip3(n8941), .op(n9577) );
  or2_1 U9357 ( .ip1(n8943), .ip2(n9577), .op(n8945) );
  nand2_1 U9358 ( .ip1(n13637), .ip2(m1Inputs[133]), .op(n9535) );
  or2_1 U9359 ( .ip1(n9535), .ip2(n9577), .op(n8944) );
  nand2_1 U9360 ( .ip1(n8945), .ip2(n8944), .op(n9576) );
  nor2_1 U9361 ( .ip1(n9540), .ip2(n6503), .op(n9578) );
  xnor2_1 U9362 ( .ip1(n9576), .ip2(n9578), .op(n9634) );
  and3_1 U9363 ( .ip1(n12578), .ip2(m1Inputs[137]), .ip3(n8946), .op(n9573) );
  inv_1 U9364 ( .ip(m1Inputs[137]), .op(n9495) );
  nor2_1 U9365 ( .ip1(n10476), .ip2(n9495), .op(n8947) );
  or2_1 U9366 ( .ip1(m1Inputs[134]), .ip2(n8947), .op(n8949) );
  or2_1 U9367 ( .ip1(n9733), .ip2(n8947), .op(n8948) );
  nand2_1 U9368 ( .ip1(n8949), .ip2(n8948), .op(n9571) );
  nor2_1 U9369 ( .ip1(n9573), .ip2(n9571), .op(n8950) );
  nand2_1 U9370 ( .ip1(m1Inputs[128]), .ip2(n14994), .op(n9570) );
  xor2_1 U9371 ( .ip1(n8950), .ip2(n9570), .op(n9633) );
  fulladder U9372 ( .a(n8953), .b(n8952), .ci(n8951), .co(n9632), .s(n4635) );
  inv_1 U9373 ( .ip(n8954), .op(n9659) );
  inv_1 U9374 ( .ip(n8955), .op(n8959) );
  nor2_1 U9375 ( .ip1(n8957), .ip2(n8956), .op(n8958) );
  nor2_1 U9376 ( .ip1(n8959), .ip2(n8958), .op(n9614) );
  nand2_1 U9377 ( .ip1(m1Inputs[131]), .ip2(\STAGE_1/weightReg [6]), .op(n9613) );
  nand2_1 U9378 ( .ip1(m1Inputs[130]), .ip2(n14835), .op(n9612) );
  inv_1 U9379 ( .ip(n8960), .op(n9650) );
  or2_1 U9380 ( .ip1(n8961), .ip2(n8962), .op(n8965) );
  or2_1 U9381 ( .ip1(n8963), .ip2(n8962), .op(n8964) );
  nand2_1 U9382 ( .ip1(n8965), .ip2(n8964), .op(n9611) );
  or2_1 U9383 ( .ip1(n8966), .ip2(n8967), .op(n8970) );
  or2_1 U9384 ( .ip1(n8968), .ip2(n8967), .op(n8969) );
  nand2_1 U9385 ( .ip1(n8970), .ip2(n8969), .op(n9610) );
  nand2_1 U9386 ( .ip1(n4672), .ip2(m1Inputs[135]), .op(n8972) );
  nor3_1 U9387 ( .ip1(n10555), .ip2(n14635), .ip3(n8971), .op(n9583) );
  or2_1 U9388 ( .ip1(n8972), .ip2(n9583), .op(n8974) );
  nand2_1 U9389 ( .ip1(n10507), .ip2(m1Inputs[136]), .op(n9494) );
  or2_1 U9390 ( .ip1(n9494), .ip2(n9583), .op(n8973) );
  nand2_1 U9391 ( .ip1(n8974), .ip2(n8973), .op(n9581) );
  nand2_1 U9392 ( .ip1(column[129]), .ip2(n13498), .op(n9582) );
  xor2_1 U9393 ( .ip1(n9581), .ip2(n9582), .op(n9609) );
  inv_1 U9394 ( .ip(n8975), .op(n9649) );
  fulladder U9395 ( .a(n8978), .b(n8977), .ci(n8976), .co(n9648), .s(n8982) );
  fulladder U9396 ( .a(n8981), .b(n8980), .ci(n8979), .co(n9657), .s(n8983) );
  fulladder U9397 ( .a(n8984), .b(n8983), .ci(n8982), .co(n9655), .s(n8987) );
  fulladder U9398 ( .a(n8987), .b(n8986), .ci(n8985), .co(n9654), .s(
        \STAGE_1/M9/sum [0]) );
  nand2_1 U9399 ( .ip1(n14629), .ip2(m1Inputs[138]), .op(n14590) );
  nor3_1 U9400 ( .ip1(n13766), .ip2(n9495), .ip3(n14590), .op(n8992) );
  nand2_1 U9401 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[138]), .op(n8988) );
  or2_1 U9402 ( .ip1(n8988), .ip2(n8992), .op(n8991) );
  nand2_1 U9403 ( .ip1(n14629), .ip2(m1Inputs[137]), .op(n8989) );
  or2_1 U9404 ( .ip1(n8989), .ip2(n8992), .op(n8990) );
  nand2_1 U9405 ( .ip1(n8991), .ip2(n8990), .op(n9009) );
  and3_1 U9406 ( .ip1(column[139]), .ip2(n15042), .ip3(n9009), .op(n9011) );
  nor2_1 U9407 ( .ip1(n8992), .ip2(n9011), .op(n14576) );
  nand2_1 U9408 ( .ip1(m1Inputs[141]), .ip2(n12981), .op(n9007) );
  nor2_1 U9409 ( .ip1(n14853), .ip2(n9530), .op(n9006) );
  nand2_1 U9410 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[139]), .op(n9005) );
  nand2_1 U9411 ( .ip1(n14876), .ip2(m1Inputs[139]), .op(n14591) );
  inv_1 U9412 ( .ip(m1Inputs[138]), .op(n14650) );
  nor3_1 U9413 ( .ip1(n13766), .ip2(n14591), .ip3(n14650), .op(n14573) );
  or2_1 U9414 ( .ip1(n14590), .ip2(n14573), .op(n8995) );
  nand2_1 U9415 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[139]), .op(n8993) );
  or2_1 U9416 ( .ip1(n8993), .ip2(n14573), .op(n8994) );
  nand2_1 U9417 ( .ip1(n8995), .ip2(n8994), .op(n14571) );
  nand2_1 U9418 ( .ip1(column[140]), .ip2(n13498), .op(n8996) );
  xor2_1 U9419 ( .ip1(n14571), .ip2(n8996), .op(n14574) );
  inv_1 U9420 ( .ip(n8997), .op(n14605) );
  nand2_1 U9421 ( .ip1(m1Inputs[136]), .ip2(n14847), .op(n8999) );
  inv_1 U9422 ( .ip(m1Inputs[135]), .op(n9467) );
  nor2_1 U9423 ( .ip1(n14902), .ip2(n9467), .op(n8998) );
  xor2_1 U9424 ( .ip1(n8999), .ip2(n8998), .op(n9000) );
  nor3_1 U9425 ( .ip1(n14842), .ip2(n9299), .ip3(n9000), .op(n9094) );
  or2_1 U9426 ( .ip1(n9000), .ip2(n9094), .op(n9003) );
  nand2_1 U9427 ( .ip1(n14816), .ip2(m1Inputs[133]), .op(n9001) );
  or2_1 U9428 ( .ip1(n9001), .ip2(n9094), .op(n9002) );
  nand2_1 U9429 ( .ip1(n9003), .ip2(n9002), .op(n9080) );
  inv_1 U9430 ( .ip(m1Inputs[143]), .op(n14581) );
  nor2_1 U9431 ( .ip1(n14581), .ip2(n14783), .op(n9098) );
  nand2_1 U9432 ( .ip1(m1Inputs[140]), .ip2(n14835), .op(n9097) );
  nand2_1 U9433 ( .ip1(m1Inputs[142]), .ip2(\STAGE_1/weightReg [5]), .op(n9096) );
  inv_1 U9434 ( .ip(n9004), .op(n9079) );
  fulladder U9435 ( .a(n9007), .b(n9006), .ci(n9005), .co(n14575), .s(n9008)
         );
  inv_1 U9436 ( .ip(n9008), .op(n9078) );
  inv_1 U9437 ( .ip(n9009), .op(n9010) );
  or2_1 U9438 ( .ip1(n9010), .ip2(n9011), .op(n9014) );
  nand2_1 U9439 ( .ip1(column[139]), .ip2(n14768), .op(n9012) );
  or2_1 U9440 ( .ip1(n9012), .ip2(n9011), .op(n9013) );
  nand2_1 U9441 ( .ip1(n9014), .ip2(n9013), .op(n9076) );
  inv_1 U9442 ( .ip(m1Inputs[139]), .op(n9449) );
  nor2_1 U9443 ( .ip1(n9449), .ip2(n14384), .op(n9065) );
  inv_1 U9444 ( .ip(m1Inputs[142]), .op(n14651) );
  nor2_1 U9445 ( .ip1(n14651), .ip2(n14783), .op(n9064) );
  nand2_1 U9446 ( .ip1(n13614), .ip2(m1Inputs[143]), .op(n9063) );
  inv_1 U9447 ( .ip(m1Inputs[141]), .op(n14636) );
  nor2_1 U9448 ( .ip1(n14636), .ip2(n4624), .op(n9068) );
  nor2_1 U9449 ( .ip1(n13766), .ip2(n9495), .op(n9067) );
  nand2_1 U9450 ( .ip1(m1Inputs[131]), .ip2(\STAGE_1/weightReg [15]), .op(
        n9066) );
  inv_1 U9451 ( .ip(n9015), .op(n14613) );
  nor3_1 U9452 ( .ip1(n6503), .ip2(n14635), .ip3(n14590), .op(n9019) );
  nand2_1 U9453 ( .ip1(m1Inputs[138]), .ip2(n14975), .op(n9017) );
  nand2_1 U9454 ( .ip1(m1Inputs[136]), .ip2(n14629), .op(n9016) );
  xor2_1 U9455 ( .ip1(n9017), .ip2(n9016), .op(n9035) );
  and3_1 U9456 ( .ip1(column[138]), .ip2(n15042), .ip3(n9035), .op(n9018) );
  nor2_1 U9457 ( .ip1(n9019), .ip2(n9018), .op(n9089) );
  nand2_1 U9458 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[134]), .op(
        n9088) );
  nand2_1 U9459 ( .ip1(n13718), .ip2(m1Inputs[135]), .op(n14585) );
  nand2_1 U9460 ( .ip1(n14847), .ip2(m1Inputs[140]), .op(n14698) );
  nand2_1 U9461 ( .ip1(m1Inputs[135]), .ip2(n13749), .op(n9284) );
  nor2_1 U9462 ( .ip1(n14698), .ip2(n9284), .op(n9023) );
  or2_1 U9463 ( .ip1(n14585), .ip2(n9023), .op(n9022) );
  nand2_1 U9464 ( .ip1(m1Inputs[140]), .ip2(\STAGE_1/weightReg [6]), .op(n9020) );
  or2_1 U9465 ( .ip1(n9020), .ip2(n9023), .op(n9021) );
  nand2_1 U9466 ( .ip1(n9022), .ip2(n9021), .op(n9083) );
  or2_1 U9467 ( .ip1(n9083), .ip2(n9023), .op(n9025) );
  nor2_1 U9468 ( .ip1(n14842), .ip2(n9530), .op(n9082) );
  or2_1 U9469 ( .ip1(n9082), .ip2(n9023), .op(n9024) );
  nand2_1 U9470 ( .ip1(n9025), .ip2(n9024), .op(n9087) );
  inv_1 U9471 ( .ip(n9026), .op(n9102) );
  nand2_1 U9472 ( .ip1(m1Inputs[139]), .ip2(\STAGE_1/weightReg [6]), .op(n9027) );
  nor2_1 U9473 ( .ip1(n14650), .ip2(n14289), .op(n9040) );
  and2_1 U9474 ( .ip1(n9040), .ip2(n9065), .op(n9031) );
  or2_1 U9475 ( .ip1(n9027), .ip2(n9031), .op(n9030) );
  nand2_1 U9476 ( .ip1(m1Inputs[138]), .ip2(n4627), .op(n9028) );
  or2_1 U9477 ( .ip1(n9028), .ip2(n9031), .op(n9029) );
  nand2_1 U9478 ( .ip1(n9030), .ip2(n9029), .op(n9054) );
  or2_1 U9479 ( .ip1(n9054), .ip2(n9031), .op(n9033) );
  inv_1 U9480 ( .ip(m1Inputs[140]), .op(n9304) );
  nor2_1 U9481 ( .ip1(n9304), .ip2(n13835), .op(n9053) );
  or2_1 U9482 ( .ip1(n9053), .ip2(n9031), .op(n9032) );
  nand2_1 U9483 ( .ip1(n9033), .ip2(n9032), .op(n9109) );
  nand2_1 U9484 ( .ip1(m1Inputs[141]), .ip2(n13637), .op(n9115) );
  nor2_1 U9485 ( .ip1(n9461), .ip2(n14853), .op(n9114) );
  nand2_1 U9486 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[137]), .op(n9113) );
  nand2_1 U9487 ( .ip1(column[138]), .ip2(n13498), .op(n9034) );
  xor2_1 U9488 ( .ip1(n9035), .ip2(n9034), .op(n9107) );
  inv_1 U9489 ( .ip(n9036), .op(n9101) );
  nor2_1 U9490 ( .ip1(n14340), .ip2(n9299), .op(n9039) );
  nor2_1 U9491 ( .ip1(n14902), .ip2(n14587), .op(n9038) );
  nor2_1 U9492 ( .ip1(n12083), .ip2(n14635), .op(n9050) );
  and2_1 U9493 ( .ip1(column[137]), .ip2(n13498), .op(n9049) );
  nand2_1 U9494 ( .ip1(column[136]), .ip2(n14768), .op(n9148) );
  inv_1 U9495 ( .ip(n9148), .op(n9048) );
  fulladder U9496 ( .a(n9039), .b(n9038), .ci(n9037), .co(n9100), .s(n9136) );
  nor2_1 U9497 ( .ip1(n9495), .ip2(n14836), .op(n9140) );
  and3_1 U9498 ( .ip1(m1Inputs[138]), .ip2(n14835), .ip3(n9140), .op(n9044) );
  or2_1 U9499 ( .ip1(n4627), .ip2(n9040), .op(n9042) );
  or2_1 U9500 ( .ip1(m1Inputs[137]), .ip2(n9040), .op(n9041) );
  nand2_1 U9501 ( .ip1(n9042), .ip2(n9041), .op(n9043) );
  nor2_1 U9502 ( .ip1(n9044), .ip2(n9043), .op(n9158) );
  or2_1 U9503 ( .ip1(n9158), .ip2(n9044), .op(n9046) );
  nor2_1 U9504 ( .ip1(n9449), .ip2(n13835), .op(n9157) );
  or2_1 U9505 ( .ip1(n9157), .ip2(n9044), .op(n9045) );
  nand2_1 U9506 ( .ip1(n9046), .ip2(n9045), .op(n9172) );
  nand2_1 U9507 ( .ip1(n13614), .ip2(m1Inputs[141]), .op(n9262) );
  nor2_1 U9508 ( .ip1(n9047), .ip2(n14581), .op(n9178) );
  nand2_1 U9509 ( .ip1(m1Inputs[130]), .ip2(\STAGE_1/weightReg [14]), .op(
        n9177) );
  fulladder U9510 ( .a(n9050), .b(n9049), .ci(n9048), .co(n9037), .s(n9051) );
  inv_1 U9511 ( .ip(n9051), .op(n9170) );
  inv_1 U9512 ( .ip(n9052), .op(n9135) );
  xor2_1 U9513 ( .ip1(n9054), .ip2(n9053), .op(n9175) );
  nand2_1 U9514 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[132]), .op(
        n9059) );
  nand2_1 U9515 ( .ip1(m1Inputs[135]), .ip2(\STAGE_1/weightReg [10]), .op(
        n9056) );
  nand2_1 U9516 ( .ip1(n14847), .ip2(m1Inputs[134]), .op(n9055) );
  nand2_1 U9517 ( .ip1(n9056), .ip2(n9055), .op(n9058) );
  nor3_1 U9518 ( .ip1(n13594), .ip2(n14587), .ip3(n14585), .op(n9085) );
  inv_1 U9519 ( .ip(n9085), .op(n9057) );
  nand2_1 U9520 ( .ip1(n9058), .ip2(n9057), .op(n9060) );
  nor3_1 U9521 ( .ip1(n14340), .ip2(n9530), .ip3(n9060), .op(n9084) );
  or2_1 U9522 ( .ip1(n9059), .ip2(n9084), .op(n9062) );
  or2_1 U9523 ( .ip1(n9060), .ip2(n9084), .op(n9061) );
  nand2_1 U9524 ( .ip1(n9062), .ip2(n9061), .op(n9174) );
  nor2_1 U9525 ( .ip1(n9304), .ip2(n14783), .op(n9181) );
  nor2_1 U9526 ( .ip1(n6503), .ip2(n14635), .op(n9180) );
  nand2_1 U9527 ( .ip1(m1Inputs[129]), .ip2(\STAGE_1/weightReg [15]), .op(
        n9179) );
  fulladder U9528 ( .a(n9065), .b(n9064), .ci(n9063), .co(n9075), .s(n9133) );
  fulladder U9529 ( .a(n9068), .b(n9067), .ci(n9066), .co(n9074), .s(n9132) );
  nor2_1 U9530 ( .ip1(n14902), .ip2(n9299), .op(n9139) );
  nor2_1 U9531 ( .ip1(n13594), .ip2(n14587), .op(n9069) );
  or2_1 U9532 ( .ip1(m1Inputs[133]), .ip2(n9069), .op(n9071) );
  or2_1 U9533 ( .ip1(n14847), .ip2(n9069), .op(n9070) );
  nand2_1 U9534 ( .ip1(n9071), .ip2(n9070), .op(n9152) );
  nor3_1 U9535 ( .ip1(n9152), .ip2(n9154), .ip3(n14340), .op(n9072) );
  nor2_1 U9536 ( .ip1(n13594), .ip2(n9299), .op(n9229) );
  and3_1 U9537 ( .ip1(\STAGE_1/weightReg [11]), .ip2(m1Inputs[134]), .ip3(
        n9229), .op(n9153) );
  or2_1 U9538 ( .ip1(n9072), .ip2(n9153), .op(n9138) );
  nor2_1 U9539 ( .ip1(n13854), .ip2(n14651), .op(n9149) );
  nor2_1 U9540 ( .ip1(n12083), .ip2(n9467), .op(n9147) );
  inv_1 U9541 ( .ip(n9073), .op(n14612) );
  fulladder U9542 ( .a(n9076), .b(n9075), .ci(n9074), .co(n14603), .s(n9077)
         );
  inv_1 U9543 ( .ip(n9077), .op(n9105) );
  fulladder U9544 ( .a(n9080), .b(n9079), .ci(n9078), .co(n14604), .s(n9081)
         );
  inv_1 U9545 ( .ip(n9081), .op(n9104) );
  xnor2_1 U9546 ( .ip1(n9083), .ip2(n9082), .op(n9112) );
  nor2_1 U9547 ( .ip1(n9085), .ip2(n9084), .op(n9111) );
  nor2_1 U9548 ( .ip1(n13854), .ip2(n14581), .op(n9117) );
  nand2_1 U9549 ( .ip1(n13614), .ip2(m1Inputs[142]), .op(n9224) );
  nand2_1 U9550 ( .ip1(m1Inputs[131]), .ip2(\STAGE_1/weightReg [14]), .op(
        n9116) );
  inv_1 U9551 ( .ip(n9086), .op(n14617) );
  nor2_1 U9552 ( .ip1(n14853), .ip2(n9299), .op(n14598) );
  nand2_1 U9553 ( .ip1(n15025), .ip2(m1Inputs[136]), .op(n14597) );
  nand2_1 U9554 ( .ip1(m1Inputs[141]), .ip2(n14835), .op(n14596) );
  nor2_1 U9555 ( .ip1(n14581), .ip2(n8942), .op(n14584) );
  nand2_1 U9556 ( .ip1(m1Inputs[142]), .ip2(n12981), .op(n14583) );
  nand2_1 U9557 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[140]), .op(
        n14582) );
  fulladder U9558 ( .a(n9089), .b(n9088), .ci(n9087), .co(n14599), .s(n9026)
         );
  inv_1 U9559 ( .ip(n9090), .op(n14609) );
  nor2_1 U9560 ( .ip1(n14842), .ip2(n14587), .op(n9093) );
  nor2_1 U9561 ( .ip1(n9495), .ip2(n14824), .op(n9092) );
  nand2_1 U9562 ( .ip1(m1Inputs[135]), .ip2(\STAGE_1/weightReg [13]), .op(
        n9091) );
  xor2_1 U9563 ( .ip1(n9092), .ip2(n9091), .op(n14586) );
  xor2_1 U9564 ( .ip1(n9093), .ip2(n14586), .op(n14579) );
  nor2_1 U9565 ( .ip1(n14585), .ip2(n14597), .op(n9095) );
  nor2_1 U9566 ( .ip1(n9095), .ip2(n9094), .op(n14578) );
  fulladder U9567 ( .a(n9098), .b(n9097), .ci(n9096), .co(n14577), .s(n9004)
         );
  inv_1 U9568 ( .ip(n9099), .op(n14608) );
  fulladder U9569 ( .a(n9102), .b(n9101), .ci(n9100), .co(n14607), .s(n9161)
         );
  fulladder U9570 ( .a(n9105), .b(n9104), .ci(n9103), .co(n14611), .s(n9106)
         );
  inv_1 U9571 ( .ip(n9106), .op(n9165) );
  fulladder U9572 ( .a(n9109), .b(n9108), .ci(n9107), .co(n9036), .s(n9169) );
  fulladder U9573 ( .a(n9112), .b(n9111), .ci(n9110), .co(n9103), .s(n9168) );
  fulladder U9574 ( .a(n9115), .b(n9114), .ci(n9113), .co(n9108), .s(n9193) );
  fulladder U9575 ( .a(n9117), .b(n9224), .ci(n9116), .co(n9110), .s(n9192) );
  nor2_1 U9576 ( .ip1(n9467), .ip2(n14384), .op(n9216) );
  and2_1 U9577 ( .ip1(n9180), .ip2(n9216), .op(n9221) );
  nor2_1 U9578 ( .ip1(n14635), .ip2(n14368), .op(n9118) );
  or2_1 U9579 ( .ip1(m1Inputs[135]), .ip2(n9118), .op(n9120) );
  or2_1 U9580 ( .ip1(n14838), .ip2(n9118), .op(n9119) );
  nand2_1 U9581 ( .ip1(n9120), .ip2(n9119), .op(n9220) );
  nand2_1 U9582 ( .ip1(m1Inputs[130]), .ip2(n15028), .op(n9222) );
  nor2_1 U9583 ( .ip1(n9220), .ip2(n9222), .op(n9121) );
  nor2_1 U9584 ( .ip1(n9221), .ip2(n9121), .op(n9211) );
  nand2_1 U9585 ( .ip1(n4619), .ip2(m1Inputs[141]), .op(n9122) );
  nand2_1 U9586 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[141]), .op(n9184) );
  nor3_1 U9587 ( .ip1(n13709), .ip2(n14651), .ip3(n9184), .op(n9126) );
  or2_1 U9588 ( .ip1(n9122), .ip2(n9126), .op(n9125) );
  nand2_1 U9589 ( .ip1(n13707), .ip2(m1Inputs[142]), .op(n9123) );
  or2_1 U9590 ( .ip1(n9123), .ip2(n9126), .op(n9124) );
  nand2_1 U9591 ( .ip1(n9125), .ip2(n9124), .op(n9235) );
  or2_1 U9592 ( .ip1(n9235), .ip2(n9126), .op(n9129) );
  nand2_1 U9593 ( .ip1(column[135]), .ip2(n14768), .op(n9234) );
  inv_1 U9594 ( .ip(n9234), .op(n9127) );
  or2_1 U9595 ( .ip1(n9127), .ip2(n9126), .op(n9128) );
  nand2_1 U9596 ( .ip1(n9129), .ip2(n9128), .op(n9210) );
  nand2_1 U9597 ( .ip1(n15025), .ip2(m1Inputs[132]), .op(n9209) );
  inv_1 U9598 ( .ip(n9130), .op(n9164) );
  fulladder U9599 ( .a(n9133), .b(n9132), .ci(n9131), .co(n9159), .s(n9243) );
  fulladder U9600 ( .a(n9136), .b(n9135), .ci(n9134), .co(n9160), .s(n9242) );
  fulladder U9601 ( .a(n9139), .b(n9138), .ci(n9137), .co(n9131), .s(n9250) );
  nand2_1 U9602 ( .ip1(m1Inputs[137]), .ip2(n13637), .op(n9291) );
  nor3_1 U9603 ( .ip1(n9449), .ip2(n14289), .ip3(n9291), .op(n9144) );
  or2_1 U9604 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n9140), .op(n9142) );
  or2_1 U9605 ( .ip1(m1Inputs[139]), .ip2(n9140), .op(n9141) );
  nand2_1 U9606 ( .ip1(n9142), .ip2(n9141), .op(n9143) );
  nor2_1 U9607 ( .ip1(n9144), .ip2(n9143), .op(n9200) );
  or2_1 U9608 ( .ip1(n9200), .ip2(n9144), .op(n9146) );
  nor2_1 U9609 ( .ip1(n9540), .ip2(n14842), .op(n9199) );
  or2_1 U9610 ( .ip1(n9199), .ip2(n9144), .op(n9145) );
  nand2_1 U9611 ( .ip1(n9146), .ip2(n9145), .op(n9206) );
  nand2_1 U9612 ( .ip1(n13614), .ip2(m1Inputs[140]), .op(n9373) );
  nor2_1 U9613 ( .ip1(n10476), .ip2(n14581), .op(n9195) );
  nand2_1 U9614 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[134]), .op(n9194) );
  fulladder U9615 ( .a(n9149), .b(n9148), .ci(n9147), .co(n9137), .s(n9150) );
  inv_1 U9616 ( .ip(n9150), .op(n9204) );
  inv_1 U9617 ( .ip(n9151), .op(n9249) );
  nor2_1 U9618 ( .ip1(n9153), .ip2(n9152), .op(n9156) );
  nor2_1 U9619 ( .ip1(n9154), .ip2(n14373), .op(n9155) );
  xor2_1 U9620 ( .ip1(n9156), .ip2(n9155), .op(n9203) );
  xor2_1 U9621 ( .ip1(n9158), .ip2(n9157), .op(n9202) );
  nor2_1 U9622 ( .ip1(n14650), .ip2(n13835), .op(n9198) );
  nand2_1 U9623 ( .ip1(m1Inputs[128]), .ip2(\STAGE_1/weightReg [15]), .op(
        n9197) );
  fulladder U9624 ( .a(n9161), .b(n9160), .ci(n9159), .co(n9073), .s(n9162) );
  inv_1 U9625 ( .ip(n9162), .op(n9239) );
  fulladder U9626 ( .a(n9165), .b(n9164), .ci(n9163), .co(n14615), .s(n9166)
         );
  inv_1 U9627 ( .ip(n9166), .op(n9238) );
  fulladder U9628 ( .a(n9169), .b(n9168), .ci(n9167), .co(n9130), .s(n9247) );
  fulladder U9629 ( .a(n9172), .b(n9171), .ci(n9170), .co(n9052), .s(n9254) );
  fulladder U9630 ( .a(n9175), .b(n9174), .ci(n9173), .co(n9134), .s(n9176) );
  inv_1 U9631 ( .ip(n9176), .op(n9253) );
  fulladder U9632 ( .a(n9262), .b(n9178), .ci(n9177), .co(n9171), .s(n9257) );
  fulladder U9633 ( .a(n9181), .b(n9180), .ci(n9179), .co(n9173), .s(n9182) );
  inv_1 U9634 ( .ip(n9182), .op(n9256) );
  nand2_1 U9635 ( .ip1(n4672), .ip2(m1Inputs[140]), .op(n9183) );
  nand2_1 U9636 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[140]), .op(n9306) );
  nor3_1 U9637 ( .ip1(n10555), .ip2(n14636), .ip3(n9306), .op(n9187) );
  or2_1 U9638 ( .ip1(n9183), .ip2(n9187), .op(n9186) );
  or2_1 U9639 ( .ip1(n9184), .ip2(n9187), .op(n9185) );
  nand2_1 U9640 ( .ip1(n9186), .ip2(n9185), .op(n9298) );
  or2_1 U9641 ( .ip1(n9298), .ip2(n9187), .op(n9190) );
  nand2_1 U9642 ( .ip1(column[134]), .ip2(n14768), .op(n9297) );
  inv_1 U9643 ( .ip(n9297), .op(n9188) );
  or2_1 U9644 ( .ip1(n9188), .ip2(n9187), .op(n9189) );
  nand2_1 U9645 ( .ip1(n9190), .ip2(n9189), .op(n9282) );
  nand2_1 U9646 ( .ip1(m1Inputs[131]), .ip2(\STAGE_1/weightReg [12]), .op(
        n9281) );
  nand2_1 U9647 ( .ip1(n14847), .ip2(m1Inputs[132]), .op(n9280) );
  fulladder U9648 ( .a(n9193), .b(n9192), .ci(n9191), .co(n9167), .s(n9320) );
  fulladder U9649 ( .a(n9373), .b(n9195), .ci(n9194), .co(n9205), .s(n9196) );
  inv_1 U9650 ( .ip(n9196), .op(n9333) );
  fulladder U9651 ( .a(n9198), .b(n9229), .ci(n9197), .co(n9201), .s(n9332) );
  xor2_1 U9652 ( .ip1(n9200), .ip2(n9199), .op(n9331) );
  fulladder U9653 ( .a(n9203), .b(n9202), .ci(n9201), .co(n9248), .s(n9328) );
  fulladder U9654 ( .a(n9206), .b(n9205), .ci(n9204), .co(n9151), .s(n9207) );
  inv_1 U9655 ( .ip(n9207), .op(n9327) );
  inv_1 U9656 ( .ip(n9208), .op(n9319) );
  fulladder U9657 ( .a(n9211), .b(n9210), .ci(n9209), .co(n9191), .s(n9326) );
  nor3_1 U9658 ( .ip1(n14650), .ip2(n4624), .ip3(n9291), .op(n9353) );
  nor2_1 U9659 ( .ip1(n9495), .ip2(n12746), .op(n9212) );
  or2_1 U9660 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n9212), .op(n9214) );
  or2_1 U9661 ( .ip1(m1Inputs[138]), .ip2(n9212), .op(n9213) );
  nand2_1 U9662 ( .ip1(n9214), .ip2(n9213), .op(n9352) );
  nand2_1 U9663 ( .ip1(n14838), .ip2(m1Inputs[134]), .op(n9354) );
  nor2_1 U9664 ( .ip1(n9352), .ip2(n9354), .op(n9215) );
  nor2_1 U9665 ( .ip1(n9353), .ip2(n9215), .op(n9276) );
  nor3_1 U9666 ( .ip1(n14635), .ip2(n14368), .ip3(n9284), .op(n9259) );
  or2_1 U9667 ( .ip1(n13749), .ip2(n9216), .op(n9218) );
  or2_1 U9668 ( .ip1(m1Inputs[136]), .ip2(n9216), .op(n9217) );
  nand2_1 U9669 ( .ip1(n9218), .ip2(n9217), .op(n9258) );
  nand2_1 U9670 ( .ip1(m1Inputs[129]), .ip2(\STAGE_1/weightReg [13]), .op(
        n9260) );
  nor2_1 U9671 ( .ip1(n9258), .ip2(n9260), .op(n9219) );
  nor2_1 U9672 ( .ip1(n9259), .ip2(n9219), .op(n9275) );
  nor2_1 U9673 ( .ip1(n9221), .ip2(n9220), .op(n9223) );
  xor2_1 U9674 ( .ip1(n9223), .ip2(n9222), .op(n9274) );
  nand2_1 U9675 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[139]), .op(n9451) );
  nor2_1 U9676 ( .ip1(n9451), .ip2(n9224), .op(n9357) );
  nor2_1 U9677 ( .ip1(n13801), .ip2(n9449), .op(n9225) );
  or2_1 U9678 ( .ip1(m1Inputs[142]), .ip2(n9225), .op(n9227) );
  or2_1 U9679 ( .ip1(n13803), .ip2(n9225), .op(n9226) );
  nand2_1 U9680 ( .ip1(n9227), .ip2(n9226), .op(n9356) );
  nand2_1 U9681 ( .ip1(m1Inputs[128]), .ip2(\STAGE_1/weightReg [14]), .op(
        n9358) );
  nor2_1 U9682 ( .ip1(n9356), .ip2(n9358), .op(n9228) );
  nor2_1 U9683 ( .ip1(n9357), .ip2(n9228), .op(n9279) );
  nor2_1 U9684 ( .ip1(n12083), .ip2(n9530), .op(n9300) );
  and2_1 U9685 ( .ip1(n9300), .ip2(n9229), .op(n9271) );
  nor2_1 U9686 ( .ip1(n13766), .ip2(n9299), .op(n9230) );
  or2_1 U9687 ( .ip1(m1Inputs[132]), .ip2(n9230), .op(n9232) );
  or2_1 U9688 ( .ip1(n14876), .ip2(n9230), .op(n9231) );
  nand2_1 U9689 ( .ip1(n9232), .ip2(n9231), .op(n9270) );
  nand2_1 U9690 ( .ip1(m1Inputs[130]), .ip2(\STAGE_1/weightReg [12]), .op(
        n9272) );
  nor2_1 U9691 ( .ip1(n9270), .ip2(n9272), .op(n9233) );
  nor2_1 U9692 ( .ip1(n9271), .ip2(n9233), .op(n9278) );
  xor2_1 U9693 ( .ip1(n9235), .ip2(n9234), .op(n9277) );
  inv_1 U9694 ( .ip(n9236), .op(n14619) );
  fulladder U9695 ( .a(n9239), .b(n9238), .ci(n9237), .co(n9236), .s(n9240) );
  inv_1 U9696 ( .ip(n9240), .op(n9662) );
  fulladder U9697 ( .a(n9243), .b(n9242), .ci(n9241), .co(n9163), .s(n9244) );
  inv_1 U9698 ( .ip(n9244), .op(n9316) );
  fulladder U9699 ( .a(n9247), .b(n9246), .ci(n9245), .co(n9237), .s(n9315) );
  fulladder U9700 ( .a(n9250), .b(n9249), .ci(n9248), .co(n9241), .s(n9251) );
  inv_1 U9701 ( .ip(n9251), .op(n9323) );
  fulladder U9702 ( .a(n9254), .b(n9253), .ci(n9252), .co(n9246), .s(n9322) );
  fulladder U9703 ( .a(n9257), .b(n9256), .ci(n9255), .co(n9252), .s(n9389) );
  nor2_1 U9704 ( .ip1(n9259), .ip2(n9258), .op(n9261) );
  xor2_1 U9705 ( .ip1(n9261), .ip2(n9260), .op(n9405) );
  nand2_1 U9706 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[138]), .op(n9506) );
  nor2_1 U9707 ( .ip1(n9506), .ip2(n9262), .op(n9267) );
  nor2_1 U9708 ( .ip1(n13082), .ip2(n14650), .op(n9263) );
  or2_1 U9709 ( .ip1(m1Inputs[141]), .ip2(n9263), .op(n9265) );
  or2_1 U9710 ( .ip1(n13803), .ip2(n9263), .op(n9264) );
  nand2_1 U9711 ( .ip1(n9265), .ip2(n9264), .op(n9266) );
  nor2_1 U9712 ( .ip1(n9267), .ip2(n9266), .op(n9412) );
  or2_1 U9713 ( .ip1(n9412), .ip2(n9267), .op(n9269) );
  nor2_1 U9714 ( .ip1(n9509), .ip2(n14373), .op(n9411) );
  or2_1 U9715 ( .ip1(n9411), .ip2(n9267), .op(n9268) );
  nand2_1 U9716 ( .ip1(n9269), .ip2(n9268), .op(n9404) );
  nor2_1 U9717 ( .ip1(n9271), .ip2(n9270), .op(n9273) );
  xor2_1 U9718 ( .ip1(n9273), .ip2(n9272), .op(n9403) );
  fulladder U9719 ( .a(n9276), .b(n9275), .ci(n9274), .co(n9325), .s(n9400) );
  fulladder U9720 ( .a(n9279), .b(n9278), .ci(n9277), .co(n9324), .s(n9399) );
  fulladder U9721 ( .a(n9282), .b(n9281), .ci(n9280), .co(n9255), .s(n9397) );
  nand2_1 U9722 ( .ip1(m1Inputs[134]), .ip2(n14835), .op(n9283) );
  nand2_1 U9723 ( .ip1(m1Inputs[134]), .ip2(\STAGE_1/weightReg [6]), .op(n9344) );
  nor3_1 U9724 ( .ip1(n9467), .ip2(n14368), .ip3(n9344), .op(n9287) );
  or2_1 U9725 ( .ip1(n9283), .ip2(n9287), .op(n9286) );
  or2_1 U9726 ( .ip1(n9284), .ip2(n9287), .op(n9285) );
  nand2_1 U9727 ( .ip1(n9286), .ip2(n9285), .op(n9416) );
  or2_1 U9728 ( .ip1(n9416), .ip2(n9287), .op(n9289) );
  nor2_1 U9729 ( .ip1(n9461), .ip2(n14824), .op(n9415) );
  or2_1 U9730 ( .ip1(n9415), .ip2(n9287), .op(n9288) );
  nand2_1 U9731 ( .ip1(n9289), .ip2(n9288), .op(n9365) );
  nand2_1 U9732 ( .ip1(m1Inputs[136]), .ip2(\STAGE_1/weightReg [5]), .op(n9290) );
  nand2_1 U9733 ( .ip1(m1Inputs[136]), .ip2(n13637), .op(n9367) );
  nor3_1 U9734 ( .ip1(n9495), .ip2(n4624), .ip3(n9367), .op(n9294) );
  or2_1 U9735 ( .ip1(n9290), .ip2(n9294), .op(n9293) );
  or2_1 U9736 ( .ip1(n9291), .ip2(n9294), .op(n9292) );
  nand2_1 U9737 ( .ip1(n9293), .ip2(n9292), .op(n9414) );
  or2_1 U9738 ( .ip1(n9414), .ip2(n9294), .op(n9296) );
  nor2_1 U9739 ( .ip1(n9540), .ip2(n14188), .op(n9413) );
  or2_1 U9740 ( .ip1(n9413), .ip2(n9294), .op(n9295) );
  nand2_1 U9741 ( .ip1(n9296), .ip2(n9295), .op(n9364) );
  xor2_1 U9742 ( .ip1(n9298), .ip2(n9297), .op(n9363) );
  nand2_1 U9743 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[132]), .op(n9515) );
  nor3_1 U9744 ( .ip1(n12083), .ip2(n9299), .ip3(n9515), .op(n9379) );
  or2_1 U9745 ( .ip1(m1Inputs[133]), .ip2(n9300), .op(n9302) );
  or2_1 U9746 ( .ip1(n14838), .ip2(n9300), .op(n9301) );
  nand2_1 U9747 ( .ip1(n9302), .ip2(n9301), .op(n9378) );
  nand2_1 U9748 ( .ip1(m1Inputs[131]), .ip2(\STAGE_1/weightReg [10]), .op(
        n9380) );
  nor2_1 U9749 ( .ip1(n9378), .ip2(n9380), .op(n9303) );
  nor2_1 U9750 ( .ip1(n9379), .ip2(n9303), .op(n9362) );
  nand2_1 U9751 ( .ip1(n4672), .ip2(m1Inputs[139]), .op(n9305) );
  nand2_1 U9752 ( .ip1(n10507), .ip2(m1Inputs[139]), .op(n9336) );
  nor3_1 U9753 ( .ip1(n10555), .ip2(n9304), .ip3(n9336), .op(n9309) );
  or2_1 U9754 ( .ip1(n9305), .ip2(n9309), .op(n9308) );
  or2_1 U9755 ( .ip1(n9306), .ip2(n9309), .op(n9307) );
  nand2_1 U9756 ( .ip1(n9308), .ip2(n9307), .op(n9351) );
  or2_1 U9757 ( .ip1(n9351), .ip2(n9309), .op(n9312) );
  nand2_1 U9758 ( .ip1(column[133]), .ip2(n14768), .op(n9350) );
  inv_1 U9759 ( .ip(n9350), .op(n9310) );
  or2_1 U9760 ( .ip1(n9310), .ip2(n9309), .op(n9311) );
  nand2_1 U9761 ( .ip1(n9312), .ip2(n9311), .op(n9361) );
  nand2_1 U9762 ( .ip1(m1Inputs[131]), .ip2(\STAGE_1/weightReg [11]), .op(
        n9360) );
  inv_1 U9763 ( .ip(n9313), .op(n9661) );
  fulladder U9764 ( .a(n9316), .b(n9315), .ci(n9314), .co(n9313), .s(n9317) );
  inv_1 U9765 ( .ip(n9317), .op(n9665) );
  fulladder U9766 ( .a(n9320), .b(n9319), .ci(n9318), .co(n9245), .s(n9385) );
  fulladder U9767 ( .a(n9323), .b(n9322), .ci(n9321), .co(n9314), .s(n9384) );
  fulladder U9768 ( .a(n9326), .b(n9325), .ci(n9324), .co(n9318), .s(n9393) );
  fulladder U9769 ( .a(n9329), .b(n9328), .ci(n9327), .co(n9208), .s(n9330) );
  inv_1 U9770 ( .ip(n9330), .op(n9392) );
  fulladder U9771 ( .a(n9333), .b(n9332), .ci(n9331), .co(n9329), .s(n9334) );
  inv_1 U9772 ( .ip(n9334), .op(n9422) );
  nand2_1 U9773 ( .ip1(n4672), .ip2(m1Inputs[138]), .op(n9335) );
  nand2_1 U9774 ( .ip1(n10507), .ip2(m1Inputs[138]), .op(n9441) );
  nor3_1 U9775 ( .ip1(n10555), .ip2(n9449), .ip3(n9441), .op(n9339) );
  or2_1 U9776 ( .ip1(n9335), .ip2(n9339), .op(n9338) );
  or2_1 U9777 ( .ip1(n9336), .ip2(n9339), .op(n9337) );
  nand2_1 U9778 ( .ip1(n9338), .ip2(n9337), .op(n9466) );
  or2_1 U9779 ( .ip1(n9466), .ip2(n9339), .op(n9342) );
  nand2_1 U9780 ( .ip1(column[132]), .ip2(n14768), .op(n9465) );
  inv_1 U9781 ( .ip(n9465), .op(n9340) );
  or2_1 U9782 ( .ip1(n9340), .ip2(n9339), .op(n9341) );
  nand2_1 U9783 ( .ip1(n9342), .ip2(n9341), .op(n9439) );
  nand2_1 U9784 ( .ip1(n14835), .ip2(m1Inputs[133]), .op(n9343) );
  nand2_1 U9785 ( .ip1(n13749), .ip2(m1Inputs[133]), .op(n9458) );
  nor3_1 U9786 ( .ip1(n14587), .ip2(n14368), .ip3(n9458), .op(n9347) );
  or2_1 U9787 ( .ip1(n9343), .ip2(n9347), .op(n9346) );
  or2_1 U9788 ( .ip1(n9344), .ip2(n9347), .op(n9345) );
  nand2_1 U9789 ( .ip1(n9346), .ip2(n9345), .op(n9478) );
  or2_1 U9790 ( .ip1(n9478), .ip2(n9347), .op(n9349) );
  nor2_1 U9791 ( .ip1(n9461), .ip2(n13594), .op(n9477) );
  or2_1 U9792 ( .ip1(n9477), .ip2(n9347), .op(n9348) );
  nand2_1 U9793 ( .ip1(n9349), .ip2(n9348), .op(n9438) );
  xor2_1 U9794 ( .ip1(n9351), .ip2(n9350), .op(n9437) );
  nor2_1 U9795 ( .ip1(n9353), .ip2(n9352), .op(n9355) );
  xor2_1 U9796 ( .ip1(n9355), .ip2(n9354), .op(n9408) );
  nor2_1 U9797 ( .ip1(n9357), .ip2(n9356), .op(n9359) );
  xor2_1 U9798 ( .ip1(n9359), .ip2(n9358), .op(n9407) );
  fulladder U9799 ( .a(n9362), .b(n9361), .ci(n9360), .co(n9395), .s(n9429) );
  fulladder U9800 ( .a(n9365), .b(n9364), .ci(n9363), .co(n9396), .s(n9428) );
  nand2_1 U9801 ( .ip1(m1Inputs[135]), .ip2(\STAGE_1/weightReg [5]), .op(n9366) );
  nand2_1 U9802 ( .ip1(m1Inputs[135]), .ip2(n13637), .op(n9469) );
  nor3_1 U9803 ( .ip1(n14635), .ip2(n4624), .ip3(n9469), .op(n9370) );
  or2_1 U9804 ( .ip1(n9366), .ip2(n9370), .op(n9369) );
  or2_1 U9805 ( .ip1(n9367), .ip2(n9370), .op(n9368) );
  nand2_1 U9806 ( .ip1(n9369), .ip2(n9368), .op(n9476) );
  or2_1 U9807 ( .ip1(n9476), .ip2(n9370), .op(n9372) );
  nor2_1 U9808 ( .ip1(n9540), .ip2(n14824), .op(n9475) );
  or2_1 U9809 ( .ip1(n9475), .ip2(n9370), .op(n9371) );
  nand2_1 U9810 ( .ip1(n9372), .ip2(n9371), .op(n9432) );
  nor3_1 U9811 ( .ip1(n10476), .ip2(n9495), .ip3(n9373), .op(n9517) );
  nor2_1 U9812 ( .ip1(n13801), .ip2(n9495), .op(n9374) );
  or2_1 U9813 ( .ip1(m1Inputs[140]), .ip2(n9374), .op(n9376) );
  or2_1 U9814 ( .ip1(n13803), .ip2(n9374), .op(n9375) );
  nand2_1 U9815 ( .ip1(n9376), .ip2(n9375), .op(n9516) );
  nand2_1 U9816 ( .ip1(m1Inputs[128]), .ip2(\STAGE_1/weightReg [12]), .op(
        n9518) );
  nor2_1 U9817 ( .ip1(n9516), .ip2(n9518), .op(n9377) );
  nor2_1 U9818 ( .ip1(n9517), .ip2(n9377), .op(n9431) );
  nor2_1 U9819 ( .ip1(n9379), .ip2(n9378), .op(n9381) );
  xor2_1 U9820 ( .ip1(n9381), .ip2(n9380), .op(n9430) );
  inv_1 U9821 ( .ip(n9382), .op(n9664) );
  fulladder U9822 ( .a(n9385), .b(n9384), .ci(n9383), .co(n9382), .s(n9386) );
  inv_1 U9823 ( .ip(n9386), .op(n9668) );
  fulladder U9824 ( .a(n9389), .b(n9388), .ci(n9387), .co(n9321), .s(n9390) );
  inv_1 U9825 ( .ip(n9390), .op(n9419) );
  fulladder U9826 ( .a(n9393), .b(n9392), .ci(n9391), .co(n9383), .s(n9394) );
  inv_1 U9827 ( .ip(n9394), .op(n9418) );
  fulladder U9828 ( .a(n9397), .b(n9396), .ci(n9395), .co(n9387), .s(n9398) );
  inv_1 U9829 ( .ip(n9398), .op(n9425) );
  fulladder U9830 ( .a(n9401), .b(n9400), .ci(n9399), .co(n9388), .s(n9402) );
  inv_1 U9831 ( .ip(n9402), .op(n9424) );
  fulladder U9832 ( .a(n9405), .b(n9404), .ci(n9403), .co(n9401), .s(n9406) );
  inv_1 U9833 ( .ip(n9406), .op(n9486) );
  fulladder U9834 ( .a(n9409), .b(n9408), .ci(n9407), .co(n9421), .s(n9410) );
  inv_1 U9835 ( .ip(n9410), .op(n9485) );
  xor2_1 U9836 ( .ip1(n9412), .ip2(n9411), .op(n9435) );
  xor2_1 U9837 ( .ip1(n9414), .ip2(n9413), .op(n9434) );
  xor2_1 U9838 ( .ip1(n9416), .ip2(n9415), .op(n9433) );
  fulladder U9839 ( .a(n9419), .b(n9418), .ci(n9417), .co(n9667), .s(n9671) );
  fulladder U9840 ( .a(n9422), .b(n9421), .ci(n9420), .co(n9391), .s(n9482) );
  fulladder U9841 ( .a(n9425), .b(n9424), .ci(n9423), .co(n9417), .s(n9426) );
  inv_1 U9842 ( .ip(n9426), .op(n9481) );
  fulladder U9843 ( .a(n9429), .b(n9428), .ci(n9427), .co(n9420), .s(n9490) );
  fulladder U9844 ( .a(n9432), .b(n9431), .ci(n9430), .co(n9427), .s(n9553) );
  fulladder U9845 ( .a(n9435), .b(n9434), .ci(n9433), .co(n9484), .s(n9436) );
  inv_1 U9846 ( .ip(n9436), .op(n9552) );
  fulladder U9847 ( .a(n9439), .b(n9438), .ci(n9437), .co(n9409), .s(n9551) );
  nand2_1 U9848 ( .ip1(n4619), .ip2(m1Inputs[137]), .op(n9440) );
  nand2_1 U9849 ( .ip1(\STAGE_1/weightReg [1]), .ip2(m1Inputs[137]), .op(n9497) );
  nor3_1 U9850 ( .ip1(n10555), .ip2(n14650), .ip3(n9497), .op(n9444) );
  or2_1 U9851 ( .ip1(n9440), .ip2(n9444), .op(n9443) );
  or2_1 U9852 ( .ip1(n9441), .ip2(n9444), .op(n9442) );
  nand2_1 U9853 ( .ip1(n9443), .ip2(n9442), .op(n9545) );
  or2_1 U9854 ( .ip1(n9545), .ip2(n9444), .op(n9447) );
  nand2_1 U9855 ( .ip1(column[131]), .ip2(n13498), .op(n9544) );
  inv_1 U9856 ( .ip(n9544), .op(n9445) );
  or2_1 U9857 ( .ip1(n9445), .ip2(n9444), .op(n9446) );
  nand2_1 U9858 ( .ip1(n9447), .ip2(n9446), .op(n9514) );
  nand2_1 U9859 ( .ip1(m1Inputs[131]), .ip2(n14994), .op(n9513) );
  nand2_1 U9860 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[136]), .op(n9450) );
  nor3_1 U9861 ( .ip1(n13801), .ip2(n9449), .ip3(n9448), .op(n9454) );
  or2_1 U9862 ( .ip1(n9450), .ip2(n9454), .op(n9453) );
  or2_1 U9863 ( .ip1(n9451), .ip2(n9454), .op(n9452) );
  nand2_1 U9864 ( .ip1(n9453), .ip2(n9452), .op(n9528) );
  or2_1 U9865 ( .ip1(n9528), .ip2(n9454), .op(n9456) );
  nor2_1 U9866 ( .ip1(n9509), .ip2(n14824), .op(n9527) );
  or2_1 U9867 ( .ip1(n9527), .ip2(n9454), .op(n9455) );
  nand2_1 U9868 ( .ip1(n9456), .ip2(n9455), .op(n9522) );
  nand2_1 U9869 ( .ip1(m1Inputs[132]), .ip2(\STAGE_1/weightReg [7]), .op(n9457) );
  nor2_1 U9870 ( .ip1(n9530), .ip2(n14836), .op(n9531) );
  and3_1 U9871 ( .ip1(n4627), .ip2(m1Inputs[133]), .ip3(n9531), .op(n9462) );
  or2_1 U9872 ( .ip1(n9457), .ip2(n9462), .op(n9460) );
  or2_1 U9873 ( .ip1(n9458), .ip2(n9462), .op(n9459) );
  nand2_1 U9874 ( .ip1(n9460), .ip2(n9459), .op(n9524) );
  or2_1 U9875 ( .ip1(n9524), .ip2(n9462), .op(n9464) );
  nor2_1 U9876 ( .ip1(n9461), .ip2(n12083), .op(n9523) );
  or2_1 U9877 ( .ip1(n9523), .ip2(n9462), .op(n9463) );
  nand2_1 U9878 ( .ip1(n9464), .ip2(n9463), .op(n9521) );
  xor2_1 U9879 ( .ip1(n9466), .ip2(n9465), .op(n9520) );
  nand2_1 U9880 ( .ip1(m1Inputs[134]), .ip2(\STAGE_1/weightReg [5]), .op(n9468) );
  nand2_1 U9881 ( .ip1(m1Inputs[134]), .ip2(n13637), .op(n9537) );
  nor3_1 U9882 ( .ip1(n9467), .ip2(n4624), .ip3(n9537), .op(n9472) );
  or2_1 U9883 ( .ip1(n9468), .ip2(n9472), .op(n9471) );
  or2_1 U9884 ( .ip1(n9469), .ip2(n9472), .op(n9470) );
  nand2_1 U9885 ( .ip1(n9471), .ip2(n9470), .op(n9526) );
  or2_1 U9886 ( .ip1(n9526), .ip2(n9472), .op(n9474) );
  nor2_1 U9887 ( .ip1(n9540), .ip2(n13594), .op(n9525) );
  or2_1 U9888 ( .ip1(n9525), .ip2(n9472), .op(n9473) );
  nand2_1 U9889 ( .ip1(n9474), .ip2(n9473), .op(n9559) );
  xnor2_1 U9890 ( .ip1(n9476), .ip2(n9475), .op(n9558) );
  xnor2_1 U9891 ( .ip1(n9478), .ip2(n9477), .op(n9557) );
  inv_1 U9892 ( .ip(n9479), .op(n9670) );
  fulladder U9893 ( .a(n9482), .b(n9481), .ci(n9480), .co(n9479), .s(n9483) );
  inv_1 U9894 ( .ip(n9483), .op(n9674) );
  fulladder U9895 ( .a(n9486), .b(n9485), .ci(n9484), .co(n9423), .s(n9487) );
  inv_1 U9896 ( .ip(n9487), .op(n9549) );
  fulladder U9897 ( .a(n9490), .b(n9489), .ci(n9488), .co(n9480), .s(n9548) );
  fulladder U9898 ( .a(n9493), .b(n9492), .ci(n9491), .co(n9488), .s(n9556) );
  nand2_1 U9899 ( .ip1(n4619), .ip2(m1Inputs[136]), .op(n9496) );
  nor3_1 U9900 ( .ip1(n10555), .ip2(n9495), .ip3(n9494), .op(n9500) );
  or2_1 U9901 ( .ip1(n9496), .ip2(n9500), .op(n9499) );
  or2_1 U9902 ( .ip1(n9497), .ip2(n9500), .op(n9498) );
  nand2_1 U9903 ( .ip1(n9499), .ip2(n9498), .op(n9588) );
  or2_1 U9904 ( .ip1(n9588), .ip2(n9500), .op(n9503) );
  nand2_1 U9905 ( .ip1(column[130]), .ip2(n13498), .op(n9587) );
  inv_1 U9906 ( .ip(n9587), .op(n9501) );
  or2_1 U9907 ( .ip1(n9501), .ip2(n9500), .op(n9502) );
  nand2_1 U9908 ( .ip1(n9503), .ip2(n9502), .op(n9565) );
  nand2_1 U9909 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[135]), .op(n9505) );
  nor3_1 U9910 ( .ip1(n13801), .ip2(n14650), .ip3(n9504), .op(n9510) );
  or2_1 U9911 ( .ip1(n9505), .ip2(n9510), .op(n9508) );
  or2_1 U9912 ( .ip1(n9506), .ip2(n9510), .op(n9507) );
  nand2_1 U9913 ( .ip1(n9508), .ip2(n9507), .op(n9608) );
  or2_1 U9914 ( .ip1(n9608), .ip2(n9510), .op(n9512) );
  nor2_1 U9915 ( .ip1(n9509), .ip2(n13594), .op(n9607) );
  or2_1 U9916 ( .ip1(n9607), .ip2(n9510), .op(n9511) );
  nand2_1 U9917 ( .ip1(n9512), .ip2(n9511), .op(n9564) );
  nand2_1 U9918 ( .ip1(m1Inputs[131]), .ip2(n14975), .op(n9563) );
  fulladder U9919 ( .a(n9515), .b(n9514), .ci(n9513), .co(n9493), .s(n9561) );
  nor2_1 U9920 ( .ip1(n9517), .ip2(n9516), .op(n9519) );
  xor2_1 U9921 ( .ip1(n9519), .ip2(n9518), .op(n9560) );
  fulladder U9922 ( .a(n9522), .b(n9521), .ci(n9520), .co(n9492), .s(n9596) );
  xor2_1 U9923 ( .ip1(n9524), .ip2(n9523), .op(n9605) );
  xor2_1 U9924 ( .ip1(n9526), .ip2(n9525), .op(n9604) );
  xor2_1 U9925 ( .ip1(n9528), .ip2(n9527), .op(n9603) );
  inv_1 U9926 ( .ip(n9529), .op(n9595) );
  nor3_1 U9927 ( .ip1(n9530), .ip2(n14368), .ip3(n9613), .op(n9567) );
  or2_1 U9928 ( .ip1(\STAGE_1/weightReg [7]), .ip2(n9531), .op(n9533) );
  or2_1 U9929 ( .ip1(m1Inputs[131]), .ip2(n9531), .op(n9532) );
  nand2_1 U9930 ( .ip1(n9533), .ip2(n9532), .op(n9566) );
  nand2_1 U9931 ( .ip1(m1Inputs[130]), .ip2(n14975), .op(n9568) );
  nor2_1 U9932 ( .ip1(n9566), .ip2(n9568), .op(n9534) );
  nor2_1 U9933 ( .ip1(n9567), .ip2(n9534), .op(n9602) );
  nand2_1 U9934 ( .ip1(n14369), .ip2(m1Inputs[133]), .op(n9536) );
  nor3_1 U9935 ( .ip1(n14587), .ip2(n12746), .ip3(n9535), .op(n9541) );
  or2_1 U9936 ( .ip1(n9536), .ip2(n9541), .op(n9539) );
  or2_1 U9937 ( .ip1(n9537), .ip2(n9541), .op(n9538) );
  nand2_1 U9938 ( .ip1(n9539), .ip2(n9538), .op(n9575) );
  or2_1 U9939 ( .ip1(n9575), .ip2(n9541), .op(n9543) );
  nor2_1 U9940 ( .ip1(n9540), .ip2(n13766), .op(n9574) );
  or2_1 U9941 ( .ip1(n9574), .ip2(n9541), .op(n9542) );
  nand2_1 U9942 ( .ip1(n9543), .ip2(n9542), .op(n9601) );
  xor2_1 U9943 ( .ip1(n9545), .ip2(n9544), .op(n9600) );
  inv_1 U9944 ( .ip(n9546), .op(n9673) );
  fulladder U9945 ( .a(n9549), .b(n9548), .ci(n9547), .co(n9546), .s(n9550) );
  inv_1 U9946 ( .ip(n9550), .op(n9677) );
  fulladder U9947 ( .a(n9553), .b(n9552), .ci(n9551), .co(n9489), .s(n9592) );
  fulladder U9948 ( .a(n9556), .b(n9555), .ci(n9554), .co(n9547), .s(n9591) );
  fulladder U9949 ( .a(n9559), .b(n9558), .ci(n9557), .co(n9491), .s(n9599) );
  fulladder U9950 ( .a(n9562), .b(n9561), .ci(n9560), .co(n9555), .s(n9598) );
  fulladder U9951 ( .a(n9565), .b(n9564), .ci(n9563), .co(n9562), .s(n9622) );
  nor2_1 U9952 ( .ip1(n9567), .ip2(n9566), .op(n9569) );
  xor2_1 U9953 ( .ip1(n9569), .ip2(n9568), .op(n9631) );
  nor2_1 U9954 ( .ip1(n9571), .ip2(n9570), .op(n9572) );
  nor2_1 U9955 ( .ip1(n9573), .ip2(n9572), .op(n9630) );
  xnor2_1 U9956 ( .ip1(n9575), .ip2(n9574), .op(n9629) );
  or2_1 U9957 ( .ip1(n9576), .ip2(n9577), .op(n9580) );
  or2_1 U9958 ( .ip1(n9578), .ip2(n9577), .op(n9579) );
  nand2_1 U9959 ( .ip1(n9580), .ip2(n9579), .op(n9628) );
  or2_1 U9960 ( .ip1(n9581), .ip2(n9583), .op(n9586) );
  inv_1 U9961 ( .ip(n9582), .op(n9584) );
  or2_1 U9962 ( .ip1(n9584), .ip2(n9583), .op(n9585) );
  nand2_1 U9963 ( .ip1(n9586), .ip2(n9585), .op(n9627) );
  xor2_1 U9964 ( .ip1(n9588), .ip2(n9587), .op(n9626) );
  inv_1 U9965 ( .ip(n9589), .op(n9676) );
  fulladder U9966 ( .a(n9592), .b(n9591), .ci(n9590), .co(n9589), .s(n9593) );
  inv_1 U9967 ( .ip(n9593), .op(n9680) );
  fulladder U9968 ( .a(n9596), .b(n9595), .ci(n9594), .co(n9554), .s(n9618) );
  fulladder U9969 ( .a(n9599), .b(n9598), .ci(n9597), .co(n9590), .s(n9617) );
  fulladder U9970 ( .a(n9602), .b(n9601), .ci(n9600), .co(n9594), .s(n9625) );
  fulladder U9971 ( .a(n9605), .b(n9604), .ci(n9603), .co(n9529), .s(n9606) );
  inv_1 U9972 ( .ip(n9606), .op(n9624) );
  xnor2_1 U9973 ( .ip1(n9608), .ip2(n9607), .op(n9642) );
  fulladder U9974 ( .a(n9611), .b(n9610), .ci(n9609), .co(n9641), .s(n8975) );
  fulladder U9975 ( .a(n9614), .b(n9613), .ci(n9612), .co(n9640), .s(n8960) );
  inv_1 U9976 ( .ip(n9615), .op(n9679) );
  fulladder U9977 ( .a(n9618), .b(n9617), .ci(n9616), .co(n9615), .s(n9619) );
  inv_1 U9978 ( .ip(n9619), .op(n9683) );
  fulladder U9979 ( .a(n9622), .b(n9621), .ci(n9620), .co(n9597), .s(n9638) );
  fulladder U9980 ( .a(n9625), .b(n9624), .ci(n9623), .co(n9616), .s(n9637) );
  fulladder U9981 ( .a(n9628), .b(n9627), .ci(n9626), .co(n9620), .s(n9646) );
  fulladder U9982 ( .a(n9631), .b(n9630), .ci(n9629), .co(n9621), .s(n9645) );
  fulladder U9983 ( .a(n9634), .b(n9633), .ci(n9632), .co(n9644), .s(n8954) );
  inv_1 U9984 ( .ip(n9635), .op(n9682) );
  fulladder U9985 ( .a(n9638), .b(n9637), .ci(n9636), .co(n9635), .s(n9639) );
  inv_1 U9986 ( .ip(n9639), .op(n9686) );
  fulladder U9987 ( .a(n9642), .b(n9641), .ci(n9640), .co(n9623), .s(n9643) );
  inv_1 U9988 ( .ip(n9643), .op(n9653) );
  fulladder U9989 ( .a(n9646), .b(n9645), .ci(n9644), .co(n9636), .s(n9647) );
  inv_1 U9990 ( .ip(n9647), .op(n9652) );
  fulladder U9991 ( .a(n9650), .b(n9649), .ci(n9648), .co(n9651), .s(n9658) );
  fulladder U9992 ( .a(n9653), .b(n9652), .ci(n9651), .co(n9685), .s(n9689) );
  fulladder U9993 ( .a(n9656), .b(n9655), .ci(n9654), .co(n9688), .s(
        \STAGE_1/M9/sum [1]) );
  fulladder U9994 ( .a(n9659), .b(n9658), .ci(n9657), .co(n9687), .s(n9656) );
  fulladder U9995 ( .a(n9662), .b(n9661), .ci(n9660), .co(n14618), .s(
        \STAGE_1/M9/sum [11]) );
  fulladder U9996 ( .a(n9665), .b(n9664), .ci(n9663), .co(n9660), .s(
        \STAGE_1/M9/sum [10]) );
  fulladder U9997 ( .a(n9668), .b(n9667), .ci(n9666), .co(n9663), .s(
        \STAGE_1/M9/sum [9]) );
  fulladder U9998 ( .a(n9671), .b(n9670), .ci(n9669), .co(n9666), .s(
        \STAGE_1/M9/sum [8]) );
  fulladder U9999 ( .a(n9674), .b(n9673), .ci(n9672), .co(n9669), .s(
        \STAGE_1/M9/sum [7]) );
  fulladder U10000 ( .a(n9677), .b(n9676), .ci(n9675), .co(n9672), .s(
        \STAGE_1/M9/sum [6]) );
  fulladder U10001 ( .a(n9680), .b(n9679), .ci(n9678), .co(n9675), .s(
        \STAGE_1/M9/sum [5]) );
  fulladder U10002 ( .a(n9683), .b(n9682), .ci(n9681), .co(n9678), .s(
        \STAGE_1/M9/sum [4]) );
  fulladder U10003 ( .a(n9686), .b(n9685), .ci(n9684), .co(n9681), .s(
        \STAGE_1/M9/sum [3]) );
  fulladder U10004 ( .a(n9689), .b(n9688), .ci(n9687), .co(n9684), .s(
        \STAGE_1/M9/sum [2]) );
  or2_1 U10005 ( .ip1(n9690), .ip2(n9691), .op(n9694) );
  or2_1 U10006 ( .ip1(n9692), .ip2(n9691), .op(n9693) );
  nand2_1 U10007 ( .ip1(n9694), .ip2(n9693), .op(n10304) );
  or2_1 U10008 ( .ip1(n9695), .ip2(n9696), .op(n9699) );
  or2_1 U10009 ( .ip1(n9697), .ip2(n9696), .op(n9698) );
  nand2_1 U10010 ( .ip1(n9699), .ip2(n9698), .op(n10303) );
  nand2_1 U10011 ( .ip1(n4672), .ip2(m1Inputs[10]), .op(n9701) );
  nor3_1 U10012 ( .ip1(n10555), .ip2(n10083), .ip3(n9700), .op(n10203) );
  or2_1 U10013 ( .ip1(n9701), .ip2(n10203), .op(n9703) );
  nand2_1 U10014 ( .ip1(n10507), .ip2(m1Inputs[11]), .op(n10171) );
  or2_1 U10015 ( .ip1(n10171), .ip2(n10203), .op(n9702) );
  nand2_1 U10016 ( .ip1(n9703), .ip2(n9702), .op(n10201) );
  nand2_1 U10017 ( .ip1(column[4]), .ip2(n13859), .op(n10202) );
  xor2_1 U10018 ( .ip1(n10201), .ip2(n10202), .op(n10302) );
  fulladder U10019 ( .a(n9706), .b(n9705), .ci(n9704), .co(n9707), .s(n6147)
         );
  inv_1 U10020 ( .ip(n9707), .op(n10325) );
  fulladder U10021 ( .a(n9710), .b(n9709), .ci(n9708), .co(n10324), .s(n9743)
         );
  or2_1 U10022 ( .ip1(n9711), .ip2(n9712), .op(n9715) );
  or2_1 U10023 ( .ip1(n9713), .ip2(n9712), .op(n9714) );
  nand2_1 U10024 ( .ip1(n9715), .ip2(n9714), .op(n10307) );
  nand2_1 U10025 ( .ip1(m1Inputs[7]), .ip2(\STAGE_1/weightReg [5]), .op(n9717)
         );
  nor3_1 U10026 ( .ip1(n10072), .ip2(n4624), .ip3(n9716), .op(n10229) );
  or2_1 U10027 ( .ip1(n9717), .ip2(n10229), .op(n9719) );
  nand2_1 U10028 ( .ip1(m1Inputs[8]), .ip2(\STAGE_1/weightReg [4]), .op(n10154) );
  or2_1 U10029 ( .ip1(n10154), .ip2(n10229), .op(n9718) );
  nand2_1 U10030 ( .ip1(n9719), .ip2(n9718), .op(n10228) );
  nor2_1 U10031 ( .ip1(n10160), .ip2(n13579), .op(n10230) );
  xnor2_1 U10032 ( .ip1(n10228), .ip2(n10230), .op(n10306) );
  nand2_1 U10033 ( .ip1(m1Inputs[5]), .ip2(\STAGE_1/weightReg [7]), .op(n9721)
         );
  nor3_1 U10034 ( .ip1(n9908), .ip2(n14368), .ip3(n9720), .op(n10208) );
  or2_1 U10035 ( .ip1(n9721), .ip2(n10208), .op(n9723) );
  nand2_1 U10036 ( .ip1(m1Inputs[6]), .ip2(n13749), .op(n10144) );
  or2_1 U10037 ( .ip1(n10144), .ip2(n10208), .op(n9722) );
  nand2_1 U10038 ( .ip1(n9723), .ip2(n9722), .op(n10207) );
  nor2_1 U10039 ( .ip1(n10150), .ip2(n13594), .op(n10209) );
  xnor2_1 U10040 ( .ip1(n10207), .ip2(n10209), .op(n10305) );
  fulladder U10041 ( .a(n9726), .b(n9725), .ci(n9724), .co(n10323), .s(n9740)
         );
  nand2_1 U10042 ( .ip1(n14838), .ip2(m1Inputs[4]), .op(n10301) );
  or2_1 U10043 ( .ip1(n9727), .ip2(n9729), .op(n9732) );
  inv_1 U10044 ( .ip(n9728), .op(n9730) );
  or2_1 U10045 ( .ip1(n9730), .ip2(n9729), .op(n9731) );
  nand2_1 U10046 ( .ip1(n9732), .ip2(n9731), .op(n10300) );
  nand2_1 U10047 ( .ip1(m1Inputs[3]), .ip2(n14994), .op(n10299) );
  nand2_1 U10048 ( .ip1(n9733), .ip2(m1Inputs[12]), .op(n10053) );
  nor3_1 U10049 ( .ip1(n10476), .ip2(n10155), .ip3(n10053), .op(n10236) );
  nor2_1 U10050 ( .ip1(n13082), .ip2(n10155), .op(n9734) );
  or2_1 U10051 ( .ip1(m1Inputs[12]), .ip2(n9734), .op(n9736) );
  or2_1 U10052 ( .ip1(n13803), .ip2(n9734), .op(n9735) );
  nand2_1 U10053 ( .ip1(n9736), .ip2(n9735), .op(n10234) );
  nor2_1 U10054 ( .ip1(n10236), .ip2(n10234), .op(n9737) );
  nand2_1 U10055 ( .ip1(m1Inputs[0]), .ip2(n15025), .op(n10233) );
  xor2_1 U10056 ( .ip1(n9737), .ip2(n10233), .op(n10321) );
  fulladder U10057 ( .a(n9740), .b(n9739), .ci(n9738), .co(n10336), .s(n9747)
         );
  fulladder U10058 ( .a(n9743), .b(n9742), .ci(n9741), .co(n10346), .s(n9746)
         );
  inv_1 U10059 ( .ip(n9744), .op(n10344) );
  fulladder U10060 ( .a(n9747), .b(n9746), .ci(n9745), .co(n9748), .s(n6165)
         );
  inv_1 U10061 ( .ip(n9748), .op(n10343) );
  fulladder U10062 ( .a(n9751), .b(n9750), .ci(n9749), .co(n10342), .s(
        \STAGE_1/M1/sum [3]) );
  inv_1 U10063 ( .ip(m1Inputs[12]), .op(n10172) );
  nor2_1 U10064 ( .ip1(n10172), .ip2(n13766), .op(n9796) );
  inv_1 U10065 ( .ip(m1Inputs[14]), .op(n9969) );
  nor2_1 U10066 ( .ip1(n9969), .ip2(n14384), .op(n9795) );
  nand2_1 U10067 ( .ip1(n14976), .ip2(m1Inputs[6]), .op(n9794) );
  inv_1 U10068 ( .ip(n9752), .op(n9800) );
  nand2_1 U10069 ( .ip1(n15025), .ip2(m1Inputs[9]), .op(n9782) );
  nand2_1 U10070 ( .ip1(m1Inputs[13]), .ip2(n14975), .op(n9781) );
  nand2_1 U10071 ( .ip1(m1Inputs[12]), .ip2(\STAGE_1/weightReg [8]), .op(n9769) );
  nand2_1 U10072 ( .ip1(m1Inputs[14]), .ip2(n13749), .op(n9767) );
  nor2_1 U10073 ( .ip1(n10155), .ip2(n14373), .op(n10403) );
  nand3_1 U10074 ( .ip1(n14847), .ip2(m1Inputs[7]), .ip3(n10403), .op(n9756)
         );
  nand2_1 U10075 ( .ip1(m1Inputs[7]), .ip2(n15028), .op(n9754) );
  nand2_1 U10076 ( .ip1(m1Inputs[9]), .ip2(n14847), .op(n9753) );
  xor2_1 U10077 ( .ip1(n9754), .ip2(n9753), .op(n9815) );
  nand3_1 U10078 ( .ip1(n14816), .ip2(m1Inputs[6]), .ip3(n9815), .op(n9755) );
  nand2_1 U10079 ( .ip1(n9756), .ip2(n9755), .op(n9810) );
  nand2_1 U10080 ( .ip1(n14876), .ip2(m1Inputs[11]), .op(n9757) );
  nand2_1 U10081 ( .ip1(n14847), .ip2(m1Inputs[11]), .op(n9784) );
  nand2_1 U10082 ( .ip1(n14629), .ip2(m1Inputs[10]), .op(n9824) );
  nor2_1 U10083 ( .ip1(n9784), .ip2(n9824), .op(n9790) );
  or2_1 U10084 ( .ip1(n9757), .ip2(n9790), .op(n9760) );
  nand2_1 U10085 ( .ip1(n14847), .ip2(m1Inputs[10]), .op(n9758) );
  or2_1 U10086 ( .ip1(n9758), .ip2(n9790), .op(n9759) );
  nand2_1 U10087 ( .ip1(n9760), .ip2(n9759), .op(n9791) );
  inv_1 U10088 ( .ip(n9791), .op(n9762) );
  nand2_1 U10089 ( .ip1(column[13]), .ip2(n13859), .op(n9761) );
  mux2_1 U10090 ( .ip1(n9762), .ip2(n9791), .s(n9761), .op(n9809) );
  inv_1 U10091 ( .ip(m1Inputs[13]), .op(n10037) );
  nor2_1 U10092 ( .ip1(n10037), .ip2(n14368), .op(n9765) );
  nor2_1 U10093 ( .ip1(n14902), .ip2(n10072), .op(n9816) );
  nand2_1 U10094 ( .ip1(n14976), .ip2(m1Inputs[5]), .op(n9764) );
  inv_1 U10095 ( .ip(n9763), .op(n9838) );
  fulladder U10096 ( .a(n9765), .b(n9816), .ci(n9764), .co(n9808), .s(n9766)
         );
  inv_1 U10097 ( .ip(n9766), .op(n9864) );
  fulladder U10098 ( .a(n9769), .b(n9768), .ci(n9767), .co(n9798), .s(n9863)
         );
  nor3_1 U10099 ( .ip1(n10072), .ip2(n6503), .ip3(n9824), .op(n9773) );
  nand2_1 U10100 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[10]), .op(n9771) );
  nand2_1 U10101 ( .ip1(m1Inputs[8]), .ip2(\STAGE_1/weightReg [10]), .op(n9770) );
  xor2_1 U10102 ( .ip1(n9771), .ip2(n9770), .op(n9882) );
  and3_1 U10103 ( .ip1(column[10]), .ip2(n13498), .ip3(n9882), .op(n9772) );
  nor2_1 U10104 ( .ip1(n9773), .ip2(n9772), .op(n9872) );
  nand2_1 U10105 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[6]), .op(n9871) );
  nand2_1 U10106 ( .ip1(n14847), .ip2(m1Inputs[7]), .op(n9774) );
  nand2_1 U10107 ( .ip1(n14847), .ip2(m1Inputs[12]), .op(n10395) );
  nand2_1 U10108 ( .ip1(m1Inputs[7]), .ip2(n13749), .op(n10147) );
  nor2_1 U10109 ( .ip1(n10395), .ip2(n10147), .op(n9778) );
  or2_1 U10110 ( .ip1(n9774), .ip2(n9778), .op(n9777) );
  nand2_1 U10111 ( .ip1(m1Inputs[12]), .ip2(\STAGE_1/weightReg [6]), .op(n9775) );
  or2_1 U10112 ( .ip1(n9775), .ip2(n9778), .op(n9776) );
  nand2_1 U10113 ( .ip1(n9777), .ip2(n9776), .op(n9934) );
  or2_1 U10114 ( .ip1(n9934), .ip2(n9778), .op(n9780) );
  nor2_1 U10115 ( .ip1(n14842), .ip2(n10088), .op(n9933) );
  or2_1 U10116 ( .ip1(n9933), .ip2(n9778), .op(n9779) );
  nand2_1 U10117 ( .ip1(n9780), .ip2(n9779), .op(n9870) );
  fulladder U10118 ( .a(n9783), .b(n9782), .ci(n9781), .co(n10400), .s(n9799)
         );
  nand4_1 U10119 ( .ip1(\STAGE_1/weightReg [11]), .ip2(m1Inputs[12]), .ip3(
        \STAGE_1/weightReg [10]), .ip4(m1Inputs[11]), .op(n10425) );
  inv_1 U10120 ( .ip(n10425), .op(n9785) );
  or2_1 U10121 ( .ip1(n9784), .ip2(n9785), .op(n9788) );
  nand2_1 U10122 ( .ip1(m1Inputs[12]), .ip2(n14629), .op(n9786) );
  or2_1 U10123 ( .ip1(n9786), .ip2(n9785), .op(n9787) );
  nand2_1 U10124 ( .ip1(n9788), .ip2(n9787), .op(n10424) );
  nand2_1 U10125 ( .ip1(column[14]), .ip2(n13859), .op(n9789) );
  xor2_1 U10126 ( .ip1(n10424), .ip2(n9789), .op(n10399) );
  nand2_1 U10127 ( .ip1(n14816), .ip2(m1Inputs[8]), .op(n10387) );
  nand2_1 U10128 ( .ip1(m1Inputs[13]), .ip2(n14994), .op(n10386) );
  inv_1 U10129 ( .ip(n9790), .op(n9793) );
  nand3_1 U10130 ( .ip1(column[13]), .ip2(n15042), .ip3(n9791), .op(n9792) );
  nand2_1 U10131 ( .ip1(n9793), .ip2(n9792), .op(n10402) );
  fulladder U10132 ( .a(n9796), .b(n9795), .ci(n9794), .co(n10401), .s(n9752)
         );
  inv_1 U10133 ( .ip(n9797), .op(n10440) );
  fulladder U10134 ( .a(n9800), .b(n9799), .ci(n9798), .co(n10439), .s(n9839)
         );
  inv_1 U10135 ( .ip(n9801), .op(n10433) );
  nor2_1 U10136 ( .ip1(n14842), .ip2(n10145), .op(n9813) );
  nor2_1 U10137 ( .ip1(n10072), .ip2(n14373), .op(n9812) );
  nand4_1 U10138 ( .ip1(\STAGE_1/weightReg [10]), .ip2(m1Inputs[11]), .ip3(
        m1Inputs[10]), .ip4(n14994), .op(n9807) );
  inv_1 U10139 ( .ip(n9807), .op(n9802) );
  or2_1 U10140 ( .ip1(n9824), .ip2(n9802), .op(n9805) );
  nand2_1 U10141 ( .ip1(m1Inputs[11]), .ip2(n14994), .op(n9803) );
  or2_1 U10142 ( .ip1(n9803), .ip2(n9802), .op(n9804) );
  nand2_1 U10143 ( .ip1(n9805), .ip2(n9804), .op(n9822) );
  nand3_1 U10144 ( .ip1(column[12]), .ip2(n15042), .ip3(n9822), .op(n9806) );
  nand2_1 U10145 ( .ip1(n9807), .ip2(n9806), .op(n9811) );
  nor2_1 U10146 ( .ip1(n14902), .ip2(n10122), .op(n10391) );
  nor2_1 U10147 ( .ip1(n6503), .ip2(n9969), .op(n10390) );
  nand2_1 U10148 ( .ip1(n14976), .ip2(m1Inputs[7]), .op(n10389) );
  fulladder U10149 ( .a(n9810), .b(n9809), .ci(n9808), .co(n10436), .s(n9763)
         );
  fulladder U10150 ( .a(n9813), .b(n9812), .ci(n9811), .co(n10438), .s(n9835)
         );
  nand2_1 U10151 ( .ip1(n14816), .ip2(m1Inputs[6]), .op(n9814) );
  xor2_1 U10152 ( .ip1(n9815), .ip2(n9814), .op(n9868) );
  and3_1 U10153 ( .ip1(\STAGE_1/weightReg [11]), .ip2(m1Inputs[7]), .ip3(n9816), .op(n9819) );
  nand2_1 U10154 ( .ip1(m1Inputs[8]), .ip2(n13718), .op(n9818) );
  nor2_1 U10155 ( .ip1(n14902), .ip2(n10145), .op(n9817) );
  xor2_1 U10156 ( .ip1(n9818), .ip2(n9817), .op(n9844) );
  nor3_1 U10157 ( .ip1(n14842), .ip2(n10166), .ip3(n9844), .op(n9845) );
  nor2_1 U10158 ( .ip1(n9819), .ip2(n9845), .op(n9867) );
  nand2_1 U10159 ( .ip1(m1Inputs[12]), .ip2(n4627), .op(n9850) );
  nand2_1 U10160 ( .ip1(m1Inputs[14]), .ip2(\STAGE_1/weightReg [5]), .op(n9849) );
  inv_1 U10161 ( .ip(n9820), .op(n9834) );
  inv_1 U10162 ( .ip(n9822), .op(n9823) );
  nand2_1 U10163 ( .ip1(column[12]), .ip2(n13859), .op(n9821) );
  mux2_1 U10164 ( .ip1(n9823), .ip2(n9822), .s(n9821), .op(n9842) );
  nand2_1 U10165 ( .ip1(m1Inputs[9]), .ip2(n14994), .op(n9917) );
  nor2_1 U10166 ( .ip1(n9824), .ip2(n9917), .op(n9826) );
  inv_1 U10167 ( .ip(n9826), .op(n9831) );
  nand2_1 U10168 ( .ip1(m1Inputs[10]), .ip2(n14994), .op(n9825) );
  or2_1 U10169 ( .ip1(n9825), .ip2(n9826), .op(n9829) );
  nand2_1 U10170 ( .ip1(n14876), .ip2(m1Inputs[9]), .op(n9827) );
  or2_1 U10171 ( .ip1(n9827), .ip2(n9826), .op(n9828) );
  nand2_1 U10172 ( .ip1(n9829), .ip2(n9828), .op(n9858) );
  nand3_1 U10173 ( .ip1(column[11]), .ip2(n15042), .ip3(n9858), .op(n9830) );
  nand2_1 U10174 ( .ip1(n9831), .ip2(n9830), .op(n9841) );
  nor2_1 U10175 ( .ip1(n10037), .ip2(n14289), .op(n9855) );
  nor2_1 U10176 ( .ip1(n10083), .ip2(n6503), .op(n9854) );
  nand2_1 U10177 ( .ip1(n14976), .ip2(m1Inputs[4]), .op(n9853) );
  inv_1 U10178 ( .ip(n9832), .op(n10407) );
  fulladder U10179 ( .a(n9835), .b(n9834), .ci(n9833), .co(n10431), .s(n9836)
         );
  inv_1 U10180 ( .ip(n9836), .op(n9861) );
  fulladder U10181 ( .a(n9839), .b(n9838), .ci(n9837), .co(n10408), .s(n9860)
         );
  fulladder U10182 ( .a(n9842), .b(n9841), .ci(n9840), .co(n9833), .s(n9843)
         );
  inv_1 U10183 ( .ip(n9843), .op(n9887) );
  or2_1 U10184 ( .ip1(n9844), .ip2(n9845), .op(n9848) );
  nand2_1 U10185 ( .ip1(n14816), .ip2(m1Inputs[5]), .op(n9846) );
  or2_1 U10186 ( .ip1(n9846), .ip2(n9845), .op(n9847) );
  nand2_1 U10187 ( .ip1(n9848), .ip2(n9847), .op(n9931) );
  fulladder U10188 ( .a(n9851), .b(n9850), .ci(n9849), .co(n9866), .s(n9852)
         );
  inv_1 U10189 ( .ip(n9852), .op(n9930) );
  fulladder U10190 ( .a(n9855), .b(n9854), .ci(n9853), .co(n9840), .s(n9929)
         );
  inv_1 U10191 ( .ip(n9856), .op(n9886) );
  nand2_1 U10192 ( .ip1(column[11]), .ip2(n13859), .op(n9857) );
  xor2_1 U10193 ( .ip1(n9858), .ip2(n9857), .op(n9928) );
  nand2_1 U10194 ( .ip1(m1Inputs[13]), .ip2(n12699), .op(n9919) );
  nor2_1 U10195 ( .ip1(n10003), .ip2(n14853), .op(n9918) );
  nand2_1 U10196 ( .ip1(m1Inputs[11]), .ip2(n4627), .op(n9915) );
  nand2_1 U10197 ( .ip1(m1Inputs[14]), .ip2(n11974), .op(n9913) );
  fulladder U10198 ( .a(n9861), .b(n9860), .ci(n9859), .co(n10406), .s(n9942)
         );
  fulladder U10199 ( .a(n9864), .b(n9863), .ci(n9862), .co(n9837), .s(n9865)
         );
  inv_1 U10200 ( .ip(n9865), .op(n9945) );
  fulladder U10201 ( .a(n9868), .b(n9867), .ci(n9866), .co(n9820), .s(n9869)
         );
  inv_1 U10202 ( .ip(n9869), .op(n9944) );
  fulladder U10203 ( .a(n9872), .b(n9871), .ci(n9870), .co(n9862), .s(n9873)
         );
  inv_1 U10204 ( .ip(n9873), .op(n9890) );
  nand2_1 U10205 ( .ip1(m1Inputs[11]), .ip2(\STAGE_1/weightReg [6]), .op(n9874) );
  nor3_1 U10206 ( .ip1(n10122), .ip2(n14289), .ip3(n9915), .op(n9878) );
  or2_1 U10207 ( .ip1(n9874), .ip2(n9878), .op(n9877) );
  nand2_1 U10208 ( .ip1(m1Inputs[10]), .ip2(n14835), .op(n9875) );
  or2_1 U10209 ( .ip1(n9875), .ip2(n9878), .op(n9876) );
  nand2_1 U10210 ( .ip1(n9877), .ip2(n9876), .op(n9907) );
  or2_1 U10211 ( .ip1(n9907), .ip2(n9878), .op(n9880) );
  nor2_1 U10212 ( .ip1(n10172), .ip2(n13835), .op(n9906) );
  or2_1 U10213 ( .ip1(n9906), .ip2(n9878), .op(n9879) );
  nand2_1 U10214 ( .ip1(n9880), .ip2(n9879), .op(n9956) );
  nand2_1 U10215 ( .ip1(m1Inputs[13]), .ip2(n13637), .op(n9962) );
  nor2_1 U10216 ( .ip1(n10150), .ip2(n14853), .op(n9961) );
  nand2_1 U10217 ( .ip1(m1Inputs[9]), .ip2(n14975), .op(n9960) );
  nand2_1 U10218 ( .ip1(column[10]), .ip2(n13859), .op(n9881) );
  xor2_1 U10219 ( .ip1(n9882), .ip2(n9881), .op(n9954) );
  inv_1 U10220 ( .ip(n9883), .op(n9889) );
  nor2_1 U10221 ( .ip1(n14340), .ip2(n10166), .op(n9893) );
  nor2_1 U10222 ( .ip1(n14902), .ip2(n9908), .op(n9892) );
  nor2_1 U10223 ( .ip1(n10072), .ip2(n13766), .op(n9903) );
  and2_1 U10224 ( .ip1(column[9]), .ip2(n13498), .op(n9902) );
  nand2_1 U10225 ( .ip1(column[8]), .ip2(n13498), .op(n9997) );
  inv_1 U10226 ( .ip(n9997), .op(n9901) );
  inv_1 U10227 ( .ip(n9884), .op(n9941) );
  fulladder U10228 ( .a(n9887), .b(n9886), .ci(n9885), .co(n9859), .s(n9948)
         );
  fulladder U10229 ( .a(n9890), .b(n9889), .ci(n9888), .co(n9943), .s(n10015)
         );
  fulladder U10230 ( .a(n9893), .b(n9892), .ci(n9891), .co(n9888), .s(n9984)
         );
  nand2_1 U10231 ( .ip1(m1Inputs[9]), .ip2(\STAGE_1/weightReg [6]), .op(n9988)
         );
  nor3_1 U10232 ( .ip1(n10122), .ip2(n14368), .ip3(n9988), .op(n9898) );
  nor2_1 U10233 ( .ip1(n10122), .ip2(n14289), .op(n9894) );
  or2_1 U10234 ( .ip1(\STAGE_1/weightReg [7]), .ip2(n9894), .op(n9896) );
  or2_1 U10235 ( .ip1(m1Inputs[9]), .ip2(n9894), .op(n9895) );
  nand2_1 U10236 ( .ip1(n9896), .ip2(n9895), .op(n9897) );
  nor2_1 U10237 ( .ip1(n9898), .ip2(n9897), .op(n10007) );
  or2_1 U10238 ( .ip1(n10007), .ip2(n9898), .op(n9900) );
  nor2_1 U10239 ( .ip1(n10083), .ip2(n12746), .op(n10006) );
  or2_1 U10240 ( .ip1(n10006), .ip2(n9898), .op(n9899) );
  nand2_1 U10241 ( .ip1(n9900), .ip2(n9899), .op(n10026) );
  nand2_1 U10242 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[13]), .op(
        n10120) );
  nand2_1 U10243 ( .ip1(m1Inputs[2]), .ip2(n14816), .op(n10031) );
  fulladder U10244 ( .a(n9903), .b(n9902), .ci(n9901), .co(n9891), .s(n9904)
         );
  inv_1 U10245 ( .ip(n9904), .op(n10024) );
  inv_1 U10246 ( .ip(n9905), .op(n9983) );
  xor2_1 U10247 ( .ip1(n9907), .ip2(n9906), .op(n10029) );
  nor2_1 U10248 ( .ip1(n13594), .ip2(n9908), .op(n9921) );
  and3_1 U10249 ( .ip1(\STAGE_1/weightReg [11]), .ip2(m1Inputs[7]), .ip3(n9921), .op(n9936) );
  nor2_1 U10250 ( .ip1(n14824), .ip2(n9908), .op(n9909) );
  or2_1 U10251 ( .ip1(m1Inputs[7]), .ip2(n9909), .op(n9911) );
  or2_1 U10252 ( .ip1(n14876), .ip2(n9909), .op(n9910) );
  nand2_1 U10253 ( .ip1(n9911), .ip2(n9910), .op(n9912) );
  nor2_1 U10254 ( .ip1(n9936), .ip2(n9912), .op(n9935) );
  nor2_1 U10255 ( .ip1(n14340), .ip2(n10088), .op(n9937) );
  xor2_1 U10256 ( .ip1(n9935), .ip2(n9937), .op(n10028) );
  nor2_1 U10257 ( .ip1(n10172), .ip2(n14783), .op(n10035) );
  nor2_1 U10258 ( .ip1(n10072), .ip2(n6503), .op(n10034) );
  nand2_1 U10259 ( .ip1(m1Inputs[1]), .ip2(n14976), .op(n10033) );
  fulladder U10260 ( .a(n9915), .b(n9914), .ci(n9913), .co(n9926), .s(n9916)
         );
  inv_1 U10261 ( .ip(n9916), .op(n9981) );
  fulladder U10262 ( .a(n9919), .b(n9918), .ci(n9917), .co(n9927), .s(n9920)
         );
  inv_1 U10263 ( .ip(n9920), .op(n9980) );
  nor2_1 U10264 ( .ip1(n14902), .ip2(n10166), .op(n9987) );
  or2_1 U10265 ( .ip1(m1Inputs[5]), .ip2(n9921), .op(n9923) );
  or2_1 U10266 ( .ip1(n14847), .ip2(n9921), .op(n9922) );
  nand2_1 U10267 ( .ip1(n9923), .ip2(n9922), .op(n10001) );
  nor3_1 U10268 ( .ip1(n10001), .ip2(n10003), .ip3(n14340), .op(n9924) );
  nor2_1 U10269 ( .ip1(n13594), .ip2(n10166), .op(n10089) );
  and3_1 U10270 ( .ip1(\STAGE_1/weightReg [11]), .ip2(m1Inputs[6]), .ip3(
        n10089), .op(n10002) );
  or2_1 U10271 ( .ip1(n9924), .ip2(n10002), .op(n9986) );
  nor2_1 U10272 ( .ip1(n6745), .ip2(n9969), .op(n9998) );
  nor2_1 U10273 ( .ip1(n13766), .ip2(n10145), .op(n9996) );
  inv_1 U10274 ( .ip(n9925), .op(n9947) );
  fulladder U10275 ( .a(n9928), .b(n9927), .ci(n9926), .co(n9885), .s(n9952)
         );
  fulladder U10276 ( .a(n9931), .b(n9930), .ci(n9929), .co(n9856), .s(n9932)
         );
  inv_1 U10277 ( .ip(n9932), .op(n9951) );
  xnor2_1 U10278 ( .ip1(n9934), .ip2(n9933), .op(n9959) );
  or2_1 U10279 ( .ip1(n9935), .ip2(n9936), .op(n9939) );
  or2_1 U10280 ( .ip1(n9937), .ip2(n9936), .op(n9938) );
  nand2_1 U10281 ( .ip1(n9939), .ip2(n9938), .op(n9958) );
  nand2_1 U10282 ( .ip1(n13614), .ip2(m1Inputs[14]), .op(n10081) );
  nand2_1 U10283 ( .ip1(m1Inputs[3]), .ip2(n14816), .op(n9963) );
  fulladder U10284 ( .a(n9942), .b(n9941), .ci(n9940), .co(n10410), .s(n10352)
         );
  fulladder U10285 ( .a(n9945), .b(n9944), .ci(n9943), .co(n9884), .s(n10011)
         );
  fulladder U10286 ( .a(n9948), .b(n9947), .ci(n9946), .co(n9940), .s(n9949)
         );
  inv_1 U10287 ( .ip(n9949), .op(n10010) );
  fulladder U10288 ( .a(n9952), .b(n9951), .ci(n9950), .co(n9946), .s(n9953)
         );
  inv_1 U10289 ( .ip(n9953), .op(n10019) );
  fulladder U10290 ( .a(n9956), .b(n9955), .ci(n9954), .co(n9883), .s(n10023)
         );
  fulladder U10291 ( .a(n9959), .b(n9958), .ci(n9957), .co(n9950), .s(n10022)
         );
  fulladder U10292 ( .a(n9962), .b(n9961), .ci(n9960), .co(n9955), .s(n10048)
         );
  fulladder U10293 ( .a(n10081), .b(n9964), .ci(n9963), .co(n9957), .s(n10047)
         );
  nor2_1 U10294 ( .ip1(n10145), .ip2(n14384), .op(n10073) );
  and2_1 U10295 ( .ip1(n10034), .ip2(n10073), .op(n10078) );
  nor2_1 U10296 ( .ip1(n10072), .ip2(n14384), .op(n9965) );
  or2_1 U10297 ( .ip1(m1Inputs[7]), .ip2(n9965), .op(n9967) );
  or2_1 U10298 ( .ip1(n14838), .ip2(n9965), .op(n9966) );
  nand2_1 U10299 ( .ip1(n9967), .ip2(n9966), .op(n10077) );
  nand2_1 U10300 ( .ip1(m1Inputs[2]), .ip2(n15028), .op(n10079) );
  nor2_1 U10301 ( .ip1(n10077), .ip2(n10079), .op(n9968) );
  nor2_1 U10302 ( .ip1(n10078), .ip2(n9968), .op(n10067) );
  nand2_1 U10303 ( .ip1(n4672), .ip2(m1Inputs[13]), .op(n9970) );
  nand2_1 U10304 ( .ip1(n13707), .ip2(m1Inputs[13]), .op(n10039) );
  nor3_1 U10305 ( .ip1(n10555), .ip2(n9969), .ip3(n10039), .op(n9974) );
  or2_1 U10306 ( .ip1(n9970), .ip2(n9974), .op(n9973) );
  nand2_1 U10307 ( .ip1(n10507), .ip2(m1Inputs[14]), .op(n9971) );
  or2_1 U10308 ( .ip1(n9971), .ip2(n9974), .op(n9972) );
  nand2_1 U10309 ( .ip1(n9973), .ip2(n9972), .op(n10095) );
  or2_1 U10310 ( .ip1(n10095), .ip2(n9974), .op(n9977) );
  nand2_1 U10311 ( .ip1(column[7]), .ip2(n13859), .op(n10094) );
  inv_1 U10312 ( .ip(n10094), .op(n9975) );
  or2_1 U10313 ( .ip1(n9975), .ip2(n9974), .op(n9976) );
  nand2_1 U10314 ( .ip1(n9977), .ip2(n9976), .op(n10066) );
  nand2_1 U10315 ( .ip1(n15025), .ip2(m1Inputs[4]), .op(n10065) );
  inv_1 U10316 ( .ip(n9978), .op(n10018) );
  fulladder U10317 ( .a(n9981), .b(n9980), .ci(n9979), .co(n10013), .s(n10101)
         );
  fulladder U10318 ( .a(n9984), .b(n9983), .ci(n9982), .co(n10014), .s(n10100)
         );
  fulladder U10319 ( .a(n9987), .b(n9986), .ci(n9985), .co(n9979), .s(n10108)
         );
  nand2_1 U10320 ( .ip1(m1Inputs[9]), .ip2(\STAGE_1/weightReg [4]), .op(n10157) );
  nor3_1 U10321 ( .ip1(n10083), .ip2(n14289), .ip3(n10157), .op(n9992) );
  or2_1 U10322 ( .ip1(n9988), .ip2(n9992), .op(n9991) );
  nand2_1 U10323 ( .ip1(m1Inputs[11]), .ip2(n11974), .op(n9989) );
  or2_1 U10324 ( .ip1(n9989), .ip2(n9992), .op(n9990) );
  nand2_1 U10325 ( .ip1(n9991), .ip2(n9990), .op(n10056) );
  or2_1 U10326 ( .ip1(n10056), .ip2(n9992), .op(n9994) );
  nor2_1 U10327 ( .ip1(n10160), .ip2(n14842), .op(n10055) );
  or2_1 U10328 ( .ip1(n10055), .ip2(n9992), .op(n9993) );
  nand2_1 U10329 ( .ip1(n9994), .ip2(n9993), .op(n10062) );
  nor2_1 U10330 ( .ip1(n13646), .ip2(n9995), .op(n10052) );
  nand2_1 U10331 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[6]), .op(n10051) );
  fulladder U10332 ( .a(n9998), .b(n9997), .ci(n9996), .co(n9985), .s(n9999)
         );
  inv_1 U10333 ( .ip(n9999), .op(n10060) );
  inv_1 U10334 ( .ip(n10000), .op(n10107) );
  nor2_1 U10335 ( .ip1(n10002), .ip2(n10001), .op(n10005) );
  nor2_1 U10336 ( .ip1(n10003), .ip2(n14373), .op(n10004) );
  xor2_1 U10337 ( .ip1(n10005), .ip2(n10004), .op(n10059) );
  xor2_1 U10338 ( .ip1(n10007), .ip2(n10006), .op(n10058) );
  nor2_1 U10339 ( .ip1(n10122), .ip2(n12746), .op(n10050) );
  nand2_1 U10340 ( .ip1(m1Inputs[0]), .ip2(n14976), .op(n10049) );
  inv_1 U10341 ( .ip(n10008), .op(n10351) );
  fulladder U10342 ( .a(n10011), .b(n10010), .ci(n10009), .co(n10008), .s(
        n10012) );
  inv_1 U10343 ( .ip(n10012), .op(n10356) );
  fulladder U10344 ( .a(n10015), .b(n10014), .ci(n10013), .co(n9925), .s(
        n10016) );
  inv_1 U10345 ( .ip(n10016), .op(n10098) );
  fulladder U10346 ( .a(n10019), .b(n10018), .ci(n10017), .co(n10009), .s(
        n10020) );
  inv_1 U10347 ( .ip(n10020), .op(n10097) );
  fulladder U10348 ( .a(n10023), .b(n10022), .ci(n10021), .co(n9978), .s(
        n10105) );
  fulladder U10349 ( .a(n10026), .b(n10025), .ci(n10024), .co(n9905), .s(
        n10112) );
  fulladder U10350 ( .a(n10029), .b(n10028), .ci(n10027), .co(n9982), .s(
        n10030) );
  inv_1 U10351 ( .ip(n10030), .op(n10111) );
  fulladder U10352 ( .a(n10032), .b(n10120), .ci(n10031), .co(n10025), .s(
        n10115) );
  fulladder U10353 ( .a(n10035), .b(n10034), .ci(n10033), .co(n10027), .s(
        n10036) );
  inv_1 U10354 ( .ip(n10036), .op(n10114) );
  nand2_1 U10355 ( .ip1(n4619), .ip2(m1Inputs[12]), .op(n10038) );
  nand2_1 U10356 ( .ip1(n10507), .ip2(m1Inputs[12]), .op(n10174) );
  nor3_1 U10357 ( .ip1(n10555), .ip2(n10037), .ip3(n10174), .op(n10042) );
  or2_1 U10358 ( .ip1(n10038), .ip2(n10042), .op(n10041) );
  or2_1 U10359 ( .ip1(n10039), .ip2(n10042), .op(n10040) );
  nand2_1 U10360 ( .ip1(n10041), .ip2(n10040), .op(n10165) );
  or2_1 U10361 ( .ip1(n10165), .ip2(n10042), .op(n10045) );
  nand2_1 U10362 ( .ip1(column[6]), .ip2(n13859), .op(n10164) );
  inv_1 U10363 ( .ip(n10164), .op(n10043) );
  or2_1 U10364 ( .ip1(n10043), .ip2(n10042), .op(n10044) );
  nand2_1 U10365 ( .ip1(n10045), .ip2(n10044), .op(n10143) );
  nand2_1 U10366 ( .ip1(m1Inputs[3]), .ip2(n15025), .op(n10142) );
  nand2_1 U10367 ( .ip1(n14847), .ip2(m1Inputs[4]), .op(n10141) );
  fulladder U10368 ( .a(n10048), .b(n10047), .ci(n10046), .co(n10021), .s(
        n10189) );
  fulladder U10369 ( .a(n10050), .b(n10089), .ci(n10049), .co(n10057), .s(
        n10199) );
  fulladder U10370 ( .a(n10053), .b(n10052), .ci(n10051), .co(n10061), .s(
        n10054) );
  inv_1 U10371 ( .ip(n10054), .op(n10198) );
  xor2_1 U10372 ( .ip1(n10056), .ip2(n10055), .op(n10197) );
  fulladder U10373 ( .a(n10059), .b(n10058), .ci(n10057), .co(n10106), .s(
        n10191) );
  fulladder U10374 ( .a(n10062), .b(n10061), .ci(n10060), .co(n10000), .s(
        n10063) );
  inv_1 U10375 ( .ip(n10063), .op(n10190) );
  inv_1 U10376 ( .ip(n10064), .op(n10188) );
  fulladder U10377 ( .a(n10067), .b(n10066), .ci(n10065), .co(n10046), .s(
        n10196) );
  nor3_1 U10378 ( .ip1(n10122), .ip2(n4624), .ip3(n10157), .op(n10215) );
  nor2_1 U10379 ( .ip1(n10155), .ip2(n12746), .op(n10068) );
  or2_1 U10380 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n10068), .op(n10070) );
  or2_1 U10381 ( .ip1(m1Inputs[10]), .ip2(n10068), .op(n10069) );
  nand2_1 U10382 ( .ip1(n10070), .ip2(n10069), .op(n10214) );
  nand2_1 U10383 ( .ip1(n14975), .ip2(m1Inputs[6]), .op(n10216) );
  nor2_1 U10384 ( .ip1(n10214), .ip2(n10216), .op(n10071) );
  nor2_1 U10385 ( .ip1(n10215), .ip2(n10071), .op(n10137) );
  nor3_1 U10386 ( .ip1(n10072), .ip2(n14368), .ip3(n10147), .op(n10117) );
  or2_1 U10387 ( .ip1(n13749), .ip2(n10073), .op(n10075) );
  or2_1 U10388 ( .ip1(m1Inputs[8]), .ip2(n10073), .op(n10074) );
  nand2_1 U10389 ( .ip1(n10075), .ip2(n10074), .op(n10116) );
  nand2_1 U10390 ( .ip1(m1Inputs[1]), .ip2(n15028), .op(n10118) );
  nor2_1 U10391 ( .ip1(n10116), .ip2(n10118), .op(n10076) );
  nor2_1 U10392 ( .ip1(n10117), .ip2(n10076), .op(n10136) );
  nor2_1 U10393 ( .ip1(n10078), .ip2(n10077), .op(n10080) );
  xor2_1 U10394 ( .ip1(n10080), .ip2(n10079), .op(n10135) );
  nor2_1 U10395 ( .ip1(n10082), .ip2(n10081), .op(n10219) );
  nor2_1 U10396 ( .ip1(n13082), .ip2(n10083), .op(n10084) );
  or2_1 U10397 ( .ip1(m1Inputs[14]), .ip2(n10084), .op(n10086) );
  or2_1 U10398 ( .ip1(n13803), .ip2(n10084), .op(n10085) );
  nand2_1 U10399 ( .ip1(n10086), .ip2(n10085), .op(n10218) );
  nand2_1 U10400 ( .ip1(m1Inputs[0]), .ip2(n14816), .op(n10220) );
  nor2_1 U10401 ( .ip1(n10218), .ip2(n10220), .op(n10087) );
  nor2_1 U10402 ( .ip1(n10219), .ip2(n10087), .op(n10140) );
  inv_1 U10403 ( .ip(\STAGE_1/weightReg [9]), .op(n12083) );
  nor2_1 U10404 ( .ip1(n12083), .ip2(n10088), .op(n10167) );
  and2_1 U10405 ( .ip1(n10167), .ip2(n10089), .op(n10132) );
  nor2_1 U10406 ( .ip1(n13766), .ip2(n10166), .op(n10090) );
  or2_1 U10407 ( .ip1(m1Inputs[4]), .ip2(n10090), .op(n10092) );
  or2_1 U10408 ( .ip1(n14876), .ip2(n10090), .op(n10091) );
  nand2_1 U10409 ( .ip1(n10092), .ip2(n10091), .op(n10131) );
  nand2_1 U10410 ( .ip1(m1Inputs[2]), .ip2(n15025), .op(n10133) );
  nor2_1 U10411 ( .ip1(n10131), .ip2(n10133), .op(n10093) );
  nor2_1 U10412 ( .ip1(n10132), .ip2(n10093), .op(n10139) );
  xor2_1 U10413 ( .ip1(n10095), .ip2(n10094), .op(n10138) );
  fulladder U10414 ( .a(n10098), .b(n10097), .ci(n10096), .co(n10355), .s(
        n10360) );
  fulladder U10415 ( .a(n10101), .b(n10100), .ci(n10099), .co(n10017), .s(
        n10102) );
  inv_1 U10416 ( .ip(n10102), .op(n10183) );
  fulladder U10417 ( .a(n10105), .b(n10104), .ci(n10103), .co(n10096), .s(
        n10182) );
  fulladder U10418 ( .a(n10108), .b(n10107), .ci(n10106), .co(n10099), .s(
        n10109) );
  inv_1 U10419 ( .ip(n10109), .op(n10186) );
  fulladder U10420 ( .a(n10112), .b(n10111), .ci(n10110), .co(n10104), .s(
        n10185) );
  fulladder U10421 ( .a(n10115), .b(n10114), .ci(n10113), .co(n10110), .s(
        n10246) );
  nor2_1 U10422 ( .ip1(n10117), .ip2(n10116), .op(n10119) );
  xor2_1 U10423 ( .ip1(n10119), .ip2(n10118), .op(n10262) );
  nor2_1 U10424 ( .ip1(n10121), .ip2(n10120), .op(n10128) );
  nor2_1 U10425 ( .ip1(n13801), .ip2(n10122), .op(n10123) );
  or2_1 U10426 ( .ip1(m1Inputs[13]), .ip2(n10123), .op(n10125) );
  or2_1 U10427 ( .ip1(n13803), .ip2(n10123), .op(n10124) );
  nand2_1 U10428 ( .ip1(n10125), .ip2(n10124), .op(n10126) );
  nor2_1 U10429 ( .ip1(n10128), .ip2(n10126), .op(n10269) );
  or2_1 U10430 ( .ip1(n10269), .ip2(n10128), .op(n10130) );
  nor2_1 U10431 ( .ip1(n10127), .ip2(n14373), .op(n10268) );
  or2_1 U10432 ( .ip1(n10268), .ip2(n10128), .op(n10129) );
  nand2_1 U10433 ( .ip1(n10130), .ip2(n10129), .op(n10261) );
  nor2_1 U10434 ( .ip1(n10132), .ip2(n10131), .op(n10134) );
  xor2_1 U10435 ( .ip1(n10134), .ip2(n10133), .op(n10260) );
  fulladder U10436 ( .a(n10137), .b(n10136), .ci(n10135), .co(n10195), .s(
        n10257) );
  fulladder U10437 ( .a(n10140), .b(n10139), .ci(n10138), .co(n10194), .s(
        n10256) );
  fulladder U10438 ( .a(n10143), .b(n10142), .ci(n10141), .co(n10113), .s(
        n10254) );
  nand2_1 U10439 ( .ip1(m1Inputs[6]), .ip2(\STAGE_1/weightReg [7]), .op(n10146) );
  nor3_1 U10440 ( .ip1(n10145), .ip2(n14368), .ip3(n10144), .op(n10151) );
  or2_1 U10441 ( .ip1(n10146), .ip2(n10151), .op(n10149) );
  or2_1 U10442 ( .ip1(n10147), .ip2(n10151), .op(n10148) );
  nand2_1 U10443 ( .ip1(n10149), .ip2(n10148), .op(n10273) );
  or2_1 U10444 ( .ip1(n10273), .ip2(n10151), .op(n10153) );
  nor2_1 U10445 ( .ip1(n10150), .ip2(n14824), .op(n10272) );
  or2_1 U10446 ( .ip1(n10272), .ip2(n10151), .op(n10152) );
  nand2_1 U10447 ( .ip1(n10153), .ip2(n10152), .op(n10227) );
  nand2_1 U10448 ( .ip1(m1Inputs[8]), .ip2(\STAGE_1/weightReg [5]), .op(n10156) );
  nor3_1 U10449 ( .ip1(n10155), .ip2(n4624), .ip3(n10154), .op(n10161) );
  or2_1 U10450 ( .ip1(n10156), .ip2(n10161), .op(n10159) );
  or2_1 U10451 ( .ip1(n10157), .ip2(n10161), .op(n10158) );
  nand2_1 U10452 ( .ip1(n10159), .ip2(n10158), .op(n10271) );
  or2_1 U10453 ( .ip1(n10271), .ip2(n10161), .op(n10163) );
  nor2_1 U10454 ( .ip1(n10160), .ip2(n14188), .op(n10270) );
  or2_1 U10455 ( .ip1(n10270), .ip2(n10161), .op(n10162) );
  nand2_1 U10456 ( .ip1(n10163), .ip2(n10162), .op(n10226) );
  xor2_1 U10457 ( .ip1(n10165), .ip2(n10164), .op(n10225) );
  nor3_1 U10458 ( .ip1(n13766), .ip2(n10166), .ip3(n10301), .op(n10238) );
  or2_1 U10459 ( .ip1(m1Inputs[5]), .ip2(n10167), .op(n10169) );
  or2_1 U10460 ( .ip1(n14838), .ip2(n10167), .op(n10168) );
  nand2_1 U10461 ( .ip1(n10169), .ip2(n10168), .op(n10237) );
  nand2_1 U10462 ( .ip1(m1Inputs[3]), .ip2(\STAGE_1/weightReg [10]), .op(
        n10239) );
  nor2_1 U10463 ( .ip1(n10237), .ip2(n10239), .op(n10170) );
  nor2_1 U10464 ( .ip1(n10238), .ip2(n10170), .op(n10224) );
  nand2_1 U10465 ( .ip1(n4672), .ip2(m1Inputs[11]), .op(n10173) );
  nor3_1 U10466 ( .ip1(n10555), .ip2(n10172), .ip3(n10171), .op(n10177) );
  or2_1 U10467 ( .ip1(n10173), .ip2(n10177), .op(n10176) );
  or2_1 U10468 ( .ip1(n10174), .ip2(n10177), .op(n10175) );
  nand2_1 U10469 ( .ip1(n10176), .ip2(n10175), .op(n10213) );
  or2_1 U10470 ( .ip1(n10213), .ip2(n10177), .op(n10180) );
  nand2_1 U10471 ( .ip1(column[5]), .ip2(n13859), .op(n10212) );
  inv_1 U10472 ( .ip(n10212), .op(n10178) );
  or2_1 U10473 ( .ip1(n10178), .ip2(n10177), .op(n10179) );
  nand2_1 U10474 ( .ip1(n10180), .ip2(n10179), .op(n10223) );
  nand2_1 U10475 ( .ip1(m1Inputs[3]), .ip2(n13718), .op(n10222) );
  fulladder U10476 ( .a(n10183), .b(n10182), .ci(n10181), .co(n10359), .s(
        n10364) );
  fulladder U10477 ( .a(n10186), .b(n10185), .ci(n10184), .co(n10181), .s(
        n10243) );
  fulladder U10478 ( .a(n10189), .b(n10188), .ci(n10187), .co(n10103), .s(
        n10242) );
  fulladder U10479 ( .a(n10192), .b(n10191), .ci(n10190), .co(n10064), .s(
        n10193) );
  inv_1 U10480 ( .ip(n10193), .op(n10250) );
  fulladder U10481 ( .a(n10196), .b(n10195), .ci(n10194), .co(n10187), .s(
        n10249) );
  fulladder U10482 ( .a(n10199), .b(n10198), .ci(n10197), .co(n10192), .s(
        n10200) );
  inv_1 U10483 ( .ip(n10200), .op(n10285) );
  or2_1 U10484 ( .ip1(n10201), .ip2(n10203), .op(n10206) );
  inv_1 U10485 ( .ip(n10202), .op(n10204) );
  or2_1 U10486 ( .ip1(n10204), .ip2(n10203), .op(n10205) );
  nand2_1 U10487 ( .ip1(n10206), .ip2(n10205), .op(n10295) );
  or2_1 U10488 ( .ip1(n10207), .ip2(n10208), .op(n10211) );
  or2_1 U10489 ( .ip1(n10209), .ip2(n10208), .op(n10210) );
  nand2_1 U10490 ( .ip1(n10211), .ip2(n10210), .op(n10294) );
  xor2_1 U10491 ( .ip1(n10213), .ip2(n10212), .op(n10293) );
  nor2_1 U10492 ( .ip1(n10215), .ip2(n10214), .op(n10217) );
  xor2_1 U10493 ( .ip1(n10217), .ip2(n10216), .op(n10265) );
  nor2_1 U10494 ( .ip1(n10219), .ip2(n10218), .op(n10221) );
  xor2_1 U10495 ( .ip1(n10221), .ip2(n10220), .op(n10264) );
  fulladder U10496 ( .a(n10224), .b(n10223), .ci(n10222), .co(n10252), .s(
        n10298) );
  fulladder U10497 ( .a(n10227), .b(n10226), .ci(n10225), .co(n10253), .s(
        n10297) );
  or2_1 U10498 ( .ip1(n10228), .ip2(n10229), .op(n10232) );
  or2_1 U10499 ( .ip1(n10230), .ip2(n10229), .op(n10231) );
  nand2_1 U10500 ( .ip1(n10232), .ip2(n10231), .op(n10288) );
  nor2_1 U10501 ( .ip1(n10234), .ip2(n10233), .op(n10235) );
  nor2_1 U10502 ( .ip1(n10236), .ip2(n10235), .op(n10287) );
  nor2_1 U10503 ( .ip1(n10238), .ip2(n10237), .op(n10240) );
  xor2_1 U10504 ( .ip1(n10240), .ip2(n10239), .op(n10286) );
  fulladder U10505 ( .a(n10243), .b(n10242), .ci(n10241), .co(n10363), .s(
        n10368) );
  fulladder U10506 ( .a(n10246), .b(n10245), .ci(n10244), .co(n10184), .s(
        n10247) );
  inv_1 U10507 ( .ip(n10247), .op(n10277) );
  fulladder U10508 ( .a(n10250), .b(n10249), .ci(n10248), .co(n10241), .s(
        n10251) );
  inv_1 U10509 ( .ip(n10251), .op(n10276) );
  fulladder U10510 ( .a(n10254), .b(n10253), .ci(n10252), .co(n10244), .s(
        n10255) );
  inv_1 U10511 ( .ip(n10255), .op(n10281) );
  fulladder U10512 ( .a(n10258), .b(n10257), .ci(n10256), .co(n10245), .s(
        n10259) );
  inv_1 U10513 ( .ip(n10259), .op(n10280) );
  fulladder U10514 ( .a(n10262), .b(n10261), .ci(n10260), .co(n10258), .s(
        n10263) );
  inv_1 U10515 ( .ip(n10263), .op(n10313) );
  fulladder U10516 ( .a(n10266), .b(n10265), .ci(n10264), .co(n10284), .s(
        n10267) );
  inv_1 U10517 ( .ip(n10267), .op(n10312) );
  xor2_1 U10518 ( .ip1(n10269), .ip2(n10268), .op(n10291) );
  xor2_1 U10519 ( .ip1(n10271), .ip2(n10270), .op(n10290) );
  xor2_1 U10520 ( .ip1(n10273), .ip2(n10272), .op(n10289) );
  inv_1 U10521 ( .ip(n10274), .op(n10367) );
  fulladder U10522 ( .a(n10277), .b(n10276), .ci(n10275), .co(n10274), .s(
        n10278) );
  inv_1 U10523 ( .ip(n10278), .op(n10372) );
  fulladder U10524 ( .a(n10281), .b(n10280), .ci(n10279), .co(n10275), .s(
        n10282) );
  inv_1 U10525 ( .ip(n10282), .op(n10310) );
  fulladder U10526 ( .a(n10285), .b(n10284), .ci(n10283), .co(n10248), .s(
        n10309) );
  fulladder U10527 ( .a(n10288), .b(n10287), .ci(n10286), .co(n10296), .s(
        n10332) );
  fulladder U10528 ( .a(n10291), .b(n10290), .ci(n10289), .co(n10311), .s(
        n10292) );
  inv_1 U10529 ( .ip(n10292), .op(n10331) );
  fulladder U10530 ( .a(n10295), .b(n10294), .ci(n10293), .co(n10266), .s(
        n10330) );
  fulladder U10531 ( .a(n10298), .b(n10297), .ci(n10296), .co(n10283), .s(
        n10316) );
  fulladder U10532 ( .a(n10301), .b(n10300), .ci(n10299), .co(n10320), .s(
        n10322) );
  fulladder U10533 ( .a(n10304), .b(n10303), .ci(n10302), .co(n10319), .s(
        n10326) );
  fulladder U10534 ( .a(n10307), .b(n10306), .ci(n10305), .co(n10318), .s(
        n10338) );
  fulladder U10535 ( .a(n10310), .b(n10309), .ci(n10308), .co(n10371), .s(
        n10376) );
  fulladder U10536 ( .a(n10313), .b(n10312), .ci(n10311), .co(n10279), .s(
        n10314) );
  inv_1 U10537 ( .ip(n10314), .op(n10329) );
  fulladder U10538 ( .a(n10317), .b(n10316), .ci(n10315), .co(n10308), .s(
        n10328) );
  fulladder U10539 ( .a(n10320), .b(n10319), .ci(n10318), .co(n10315), .s(
        n10335) );
  fulladder U10540 ( .a(n10323), .b(n10322), .ci(n10321), .co(n10334), .s(
        n10337) );
  fulladder U10541 ( .a(n10326), .b(n10325), .ci(n10324), .co(n10333), .s(
        n10348) );
  fulladder U10542 ( .a(n10329), .b(n10328), .ci(n10327), .co(n10375), .s(
        n10380) );
  fulladder U10543 ( .a(n10332), .b(n10331), .ci(n10330), .co(n10317), .s(
        n10341) );
  fulladder U10544 ( .a(n10335), .b(n10334), .ci(n10333), .co(n10327), .s(
        n10340) );
  fulladder U10545 ( .a(n10338), .b(n10337), .ci(n10336), .co(n10339), .s(
        n10347) );
  fulladder U10546 ( .a(n10341), .b(n10340), .ci(n10339), .co(n10379), .s(
        n10384) );
  fulladder U10547 ( .a(n10344), .b(n10343), .ci(n10342), .co(n10345), .s(
        \STAGE_1/M1/sum [4]) );
  inv_1 U10548 ( .ip(n10345), .op(n10383) );
  fulladder U10549 ( .a(n10348), .b(n10347), .ci(n10346), .co(n10382), .s(
        n9744) );
  inv_1 U10550 ( .ip(n10349), .op(\STAGE_1/M1/sum [14]) );
  fulladder U10551 ( .a(n10352), .b(n10351), .ci(n10350), .co(n10409), .s(
        n10353) );
  inv_1 U10552 ( .ip(n10353), .op(\STAGE_1/M1/sum [13]) );
  fulladder U10553 ( .a(n10356), .b(n10355), .ci(n10354), .co(n10350), .s(
        n10357) );
  inv_1 U10554 ( .ip(n10357), .op(\STAGE_1/M1/sum [12]) );
  fulladder U10555 ( .a(n10360), .b(n10359), .ci(n10358), .co(n10354), .s(
        n10361) );
  inv_1 U10556 ( .ip(n10361), .op(\STAGE_1/M1/sum [11]) );
  fulladder U10557 ( .a(n10364), .b(n10363), .ci(n10362), .co(n10358), .s(
        n10365) );
  inv_1 U10558 ( .ip(n10365), .op(\STAGE_1/M1/sum [10]) );
  fulladder U10559 ( .a(n10368), .b(n10367), .ci(n10366), .co(n10362), .s(
        n10369) );
  inv_1 U10560 ( .ip(n10369), .op(\STAGE_1/M1/sum [9]) );
  fulladder U10561 ( .a(n10372), .b(n10371), .ci(n10370), .co(n10366), .s(
        n10373) );
  inv_1 U10562 ( .ip(n10373), .op(\STAGE_1/M1/sum [8]) );
  fulladder U10563 ( .a(n10376), .b(n10375), .ci(n10374), .co(n10370), .s(
        n10377) );
  inv_1 U10564 ( .ip(n10377), .op(\STAGE_1/M1/sum [7]) );
  fulladder U10565 ( .a(n10380), .b(n10379), .ci(n10378), .co(n10374), .s(
        n10381) );
  inv_1 U10566 ( .ip(n10381), .op(\STAGE_1/M1/sum [6]) );
  fulladder U10567 ( .a(n10384), .b(n10383), .ci(n10382), .co(n10378), .s(
        n10385) );
  inv_1 U10568 ( .ip(n10385), .op(\STAGE_1/M1/sum [5]) );
  fulladder U10569 ( .a(n10388), .b(n10387), .ci(n10386), .co(n10393), .s(
        n10398) );
  fulladder U10570 ( .a(n10391), .b(n10390), .ci(n10389), .co(n10392), .s(
        n10437) );
  xor2_1 U10571 ( .ip1(n10393), .ip2(n10392), .op(n10394) );
  xor2_1 U10572 ( .ip1(n10395), .ip2(n10394), .op(n10423) );
  nand2_1 U10573 ( .ip1(m1Inputs[10]), .ip2(n15028), .op(n10397) );
  nand2_1 U10574 ( .ip1(m1Inputs[13]), .ip2(n14629), .op(n10396) );
  xor2_1 U10575 ( .ip1(n10397), .ip2(n10396), .op(n10421) );
  fulladder U10576 ( .a(n10400), .b(n10399), .ci(n10398), .co(n10405), .s(
        n10441) );
  fulladder U10577 ( .a(n10403), .b(n10402), .ci(n10401), .co(n10404), .s(
        n9797) );
  xor2_1 U10578 ( .ip1(n10405), .ip2(n10404), .op(n10415) );
  fulladder U10579 ( .a(n10408), .b(n10407), .ci(n10406), .co(n10413), .s(
        n10411) );
  fulladder U10580 ( .a(n10411), .b(n10410), .ci(n10409), .co(n10412), .s(
        n10349) );
  xor2_1 U10581 ( .ip1(n10413), .ip2(n10412), .op(n10414) );
  xor2_1 U10582 ( .ip1(n10415), .ip2(n10414), .op(n10416) );
  xor2_1 U10583 ( .ip1(n10417), .ip2(n10416), .op(n10419) );
  nand2_1 U10584 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[14]), .op(
        n10418) );
  xor2_1 U10585 ( .ip1(n10419), .ip2(n10418), .op(n10420) );
  xor2_1 U10586 ( .ip1(n10421), .ip2(n10420), .op(n10422) );
  xor2_1 U10587 ( .ip1(n10423), .ip2(n10422), .op(n10451) );
  nand2_1 U10588 ( .ip1(n15042), .ip2(column[15]), .op(n10428) );
  nand3_1 U10589 ( .ip1(column[14]), .ip2(n10424), .ip3(n14768), .op(n10426)
         );
  nand2_1 U10590 ( .ip1(n10426), .ip2(n10425), .op(n10427) );
  xor2_1 U10591 ( .ip1(n10428), .ip2(n10427), .op(n10449) );
  nand2_1 U10592 ( .ip1(m1Inputs[8]), .ip2(n14976), .op(n10430) );
  nand2_1 U10593 ( .ip1(m1Inputs[9]), .ip2(n14816), .op(n10429) );
  xor2_1 U10594 ( .ip1(n10430), .ip2(n10429), .op(n10435) );
  fulladder U10595 ( .a(n10433), .b(n10432), .ci(n10431), .co(n10434), .s(
        n9832) );
  xor2_1 U10596 ( .ip1(n10435), .ip2(n10434), .op(n10445) );
  fulladder U10597 ( .a(n10438), .b(n10437), .ci(n10436), .co(n10443), .s(
        n10432) );
  fulladder U10598 ( .a(n10441), .b(n10440), .ci(n10439), .co(n10442), .s(
        n9801) );
  xor2_1 U10599 ( .ip1(n10443), .ip2(n10442), .op(n10444) );
  xor2_1 U10600 ( .ip1(n10445), .ip2(n10444), .op(n10447) );
  nand2_1 U10601 ( .ip1(n15025), .ip2(m1Inputs[11]), .op(n10446) );
  xor2_1 U10602 ( .ip1(n10447), .ip2(n10446), .op(n10448) );
  xor2_1 U10603 ( .ip1(n10449), .ip2(n10448), .op(n10450) );
  xor2_1 U10604 ( .ip1(n10451), .ip2(n10450), .op(\STAGE_1/M1/sum [15]) );
  nor2_1 U10605 ( .ip1(n14902), .ip2(n10866), .op(n10897) );
  nor2_1 U10606 ( .ip1(n13594), .ip2(n10867), .op(n10491) );
  or2_1 U10607 ( .ip1(m1Inputs[21]), .ip2(n10491), .op(n10453) );
  or2_1 U10608 ( .ip1(n14847), .ip2(n10491), .op(n10452) );
  nand2_1 U10609 ( .ip1(n10453), .ip2(n10452), .op(n10459) );
  nor3_1 U10610 ( .ip1(n10459), .ip2(n10461), .ip3(n14340), .op(n10454) );
  nor2_1 U10611 ( .ip1(n13594), .ip2(n10866), .op(n10598) );
  and3_1 U10612 ( .ip1(n13718), .ip2(m1Inputs[22]), .ip3(n10598), .op(n10460)
         );
  or2_1 U10613 ( .ip1(n10454), .ip2(n10460), .op(n10896) );
  inv_1 U10614 ( .ip(m1Inputs[30]), .op(n10828) );
  nor2_1 U10615 ( .ip1(n13854), .ip2(n10828), .op(n10466) );
  nand2_1 U10616 ( .ip1(column[24]), .ip2(n13859), .op(n10482) );
  nor2_1 U10617 ( .ip1(n12083), .ip2(n10734), .op(n10465) );
  inv_1 U10618 ( .ip(n10455), .op(n10949) );
  nor2_1 U10619 ( .ip1(n10753), .ip2(n14836), .op(n10468) );
  and3_1 U10620 ( .ip1(m1Inputs[26]), .ip2(n4627), .ip3(n10468), .op(n10478)
         );
  nor2_1 U10621 ( .ip1(n10827), .ip2(n14836), .op(n10484) );
  or2_1 U10622 ( .ip1(\STAGE_1/weightReg [7]), .ip2(n10484), .op(n10457) );
  or2_1 U10623 ( .ip1(m1Inputs[25]), .ip2(n10484), .op(n10456) );
  nand2_1 U10624 ( .ip1(n10457), .ip2(n10456), .op(n10458) );
  nor2_1 U10625 ( .ip1(n10478), .ip2(n10458), .op(n10477) );
  nor2_1 U10626 ( .ip1(n10751), .ip2(n4624), .op(n10479) );
  xor2_1 U10627 ( .ip1(n10477), .ip2(n10479), .op(n10607) );
  nor2_1 U10628 ( .ip1(n10827), .ip2(n12746), .op(n10597) );
  nand2_1 U10629 ( .ip1(m1Inputs[16]), .ip2(n14976), .op(n10596) );
  nor2_1 U10630 ( .ip1(n10460), .ip2(n10459), .op(n10463) );
  nor2_1 U10631 ( .ip1(n10461), .ip2(n14340), .op(n10462) );
  xor2_1 U10632 ( .ip1(n10463), .ip2(n10462), .op(n10605) );
  inv_1 U10633 ( .ip(n10464), .op(n10948) );
  fulladder U10634 ( .a(n10466), .b(n10482), .ci(n10465), .co(n10895), .s(
        n10467) );
  inv_1 U10635 ( .ip(n10467), .op(n10610) );
  nor3_1 U10636 ( .ip1(n10751), .ip2(n14836), .ip3(n10530), .op(n10473) );
  or2_1 U10637 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n10468), .op(n10470) );
  or2_1 U10638 ( .ip1(m1Inputs[27]), .ip2(n10468), .op(n10469) );
  nand2_1 U10639 ( .ip1(n10470), .ip2(n10469), .op(n10471) );
  nor2_1 U10640 ( .ip1(n10473), .ip2(n10471), .op(n10604) );
  or2_1 U10641 ( .ip1(n10604), .ip2(n10473), .op(n10475) );
  nor2_1 U10642 ( .ip1(n10472), .ip2(n14842), .op(n10603) );
  or2_1 U10643 ( .ip1(n10603), .ip2(n10473), .op(n10474) );
  nand2_1 U10644 ( .ip1(n10475), .ip2(n10474), .op(n10609) );
  inv_1 U10645 ( .ip(m1Inputs[31]), .op(n10738) );
  nor2_1 U10646 ( .ip1(n10476), .ip2(n10738), .op(n10601) );
  nand2_1 U10647 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[22]), .op(
        n10599) );
  or2_1 U10648 ( .ip1(n10477), .ip2(n10478), .op(n10481) );
  or2_1 U10649 ( .ip1(n10479), .ip2(n10478), .op(n10480) );
  nand2_1 U10650 ( .ip1(n10481), .ip2(n10480), .op(n10884) );
  nor2_1 U10651 ( .ip1(n13570), .ip2(n10738), .op(n10500) );
  nand2_1 U10652 ( .ip1(m1Inputs[18]), .ip2(n14816), .op(n10499) );
  nor2_1 U10653 ( .ip1(n12083), .ip2(n10812), .op(n10870) );
  and2_1 U10654 ( .ip1(column[25]), .ip2(n13498), .op(n10869) );
  inv_1 U10655 ( .ip(n10482), .op(n10868) );
  inv_1 U10656 ( .ip(n10483), .op(n10882) );
  nand2_1 U10657 ( .ip1(m1Inputs[27]), .ip2(n13749), .op(n10485) );
  nor2_1 U10658 ( .ip1(n10751), .ip2(n14368), .op(n10891) );
  and2_1 U10659 ( .ip1(n10484), .ip2(n10891), .op(n10856) );
  or2_1 U10660 ( .ip1(n10485), .ip2(n10856), .op(n10488) );
  nand2_1 U10661 ( .ip1(m1Inputs[26]), .ip2(\STAGE_1/weightReg [7]), .op(
        n10486) );
  or2_1 U10662 ( .ip1(n10486), .ip2(n10856), .op(n10487) );
  nand2_1 U10663 ( .ip1(n10488), .ip2(n10487), .op(n10855) );
  nor2_1 U10664 ( .ip1(n11033), .ip2(n8942), .op(n10857) );
  xor2_1 U10665 ( .ip1(n10855), .ip2(n10857), .op(n10888) );
  nand2_1 U10666 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[20]), .op(
        n10494) );
  nand2_1 U10667 ( .ip1(m1Inputs[23]), .ip2(\STAGE_1/weightReg [10]), .op(
        n10490) );
  nand2_1 U10668 ( .ip1(n13718), .ip2(m1Inputs[22]), .op(n10489) );
  nand2_1 U10669 ( .ip1(n10490), .ip2(n10489), .op(n10492) );
  nor2_1 U10670 ( .ip1(n14824), .ip2(n10734), .op(n10778) );
  nand2_1 U10671 ( .ip1(n10778), .ip2(n10491), .op(n10911) );
  nand2_1 U10672 ( .ip1(n10492), .ip2(n10911), .op(n10495) );
  nor3_1 U10673 ( .ip1(n14340), .ip2(n10493), .ip3(n10495), .op(n10912) );
  or2_1 U10674 ( .ip1(n10494), .ip2(n10912), .op(n10497) );
  or2_1 U10675 ( .ip1(n10495), .ip2(n10912), .op(n10496) );
  nand2_1 U10676 ( .ip1(n10497), .ip2(n10496), .op(n10887) );
  nor2_1 U10677 ( .ip1(n11033), .ip2(n14783), .op(n10503) );
  nor2_1 U10678 ( .ip1(n6503), .ip2(n10812), .op(n10540) );
  nand2_1 U10679 ( .ip1(m1Inputs[17]), .ip2(n14976), .op(n10502) );
  inv_1 U10680 ( .ip(n10498), .op(n10961) );
  fulladder U10681 ( .a(n10501), .b(n10500), .ci(n10499), .co(n10883), .s(
        n10516) );
  fulladder U10682 ( .a(n10503), .b(n10540), .ci(n10502), .co(n10886), .s(
        n10504) );
  inv_1 U10683 ( .ip(n10504), .op(n10515) );
  nand2_1 U10684 ( .ip1(n4672), .ip2(m1Inputs[28]), .op(n10506) );
  inv_1 U10685 ( .ip(m1Inputs[29]), .op(n10813) );
  nor3_1 U10686 ( .ip1(n10555), .ip2(n10813), .ip3(n10505), .op(n10510) );
  or2_1 U10687 ( .ip1(n10506), .ip2(n10510), .op(n10509) );
  nand2_1 U10688 ( .ip1(n10507), .ip2(m1Inputs[29]), .op(n10554) );
  or2_1 U10689 ( .ip1(n10554), .ip2(n10510), .op(n10508) );
  nand2_1 U10690 ( .ip1(n10509), .ip2(n10508), .op(n10574) );
  or2_1 U10691 ( .ip1(n10574), .ip2(n10510), .op(n10513) );
  nand2_1 U10692 ( .ip1(column[22]), .ip2(n13859), .op(n10573) );
  inv_1 U10693 ( .ip(n10573), .op(n10511) );
  or2_1 U10694 ( .ip1(n10511), .ip2(n10510), .op(n10512) );
  nand2_1 U10695 ( .ip1(n10513), .ip2(n10512), .op(n10562) );
  nand2_1 U10696 ( .ip1(m1Inputs[19]), .ip2(n15025), .op(n10561) );
  nand2_1 U10697 ( .ip1(n13718), .ip2(m1Inputs[20]), .op(n10560) );
  fulladder U10698 ( .a(n10516), .b(n10515), .ci(n10514), .co(n10960), .s(
        n10656) );
  nor3_1 U10699 ( .ip1(n10812), .ip2(n14368), .ip3(n10777), .op(n10538) );
  nor2_1 U10700 ( .ip1(n10734), .ip2(n14384), .op(n10539) );
  or2_1 U10701 ( .ip1(n13749), .ip2(n10539), .op(n10518) );
  or2_1 U10702 ( .ip1(m1Inputs[24]), .ip2(n10539), .op(n10517) );
  nand2_1 U10703 ( .ip1(n10518), .ip2(n10517), .op(n10536) );
  nor2_1 U10704 ( .ip1(n10538), .ip2(n10536), .op(n10519) );
  nand2_1 U10705 ( .ip1(m1Inputs[17]), .ip2(n15028), .op(n10535) );
  xor2_1 U10706 ( .ip1(n10519), .ip2(n10535), .op(n10672) );
  or2_1 U10707 ( .ip1(n10520), .ip2(n10521), .op(n10524) );
  or2_1 U10708 ( .ip1(n10522), .ip2(n10521), .op(n10523) );
  nand2_1 U10709 ( .ip1(n10524), .ip2(n10523), .op(n10671) );
  and2_1 U10710 ( .ip1(n10525), .ip2(n10598), .op(n10553) );
  nor2_1 U10711 ( .ip1(n12083), .ip2(n10866), .op(n10526) );
  or2_1 U10712 ( .ip1(m1Inputs[20]), .ip2(n10526), .op(n10528) );
  or2_1 U10713 ( .ip1(n14876), .ip2(n10526), .op(n10527) );
  nand2_1 U10714 ( .ip1(n10528), .ip2(n10527), .op(n10551) );
  nor2_1 U10715 ( .ip1(n10553), .ip2(n10551), .op(n10529) );
  nand2_1 U10716 ( .ip1(m1Inputs[18]), .ip2(n15025), .op(n10550) );
  xor2_1 U10717 ( .ip1(n10529), .ip2(n10550), .op(n10670) );
  nor3_1 U10718 ( .ip1(n10827), .ip2(n4624), .ip3(n10530), .op(n10637) );
  nor2_1 U10719 ( .ip1(n10753), .ip2(n12746), .op(n10531) );
  or2_1 U10720 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n10531), .op(n10533) );
  or2_1 U10721 ( .ip1(m1Inputs[26]), .ip2(n10531), .op(n10532) );
  nand2_1 U10722 ( .ip1(n10533), .ip2(n10532), .op(n10636) );
  nand2_1 U10723 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[22]), .op(
        n10638) );
  nor2_1 U10724 ( .ip1(n10636), .ip2(n10638), .op(n10534) );
  nor2_1 U10725 ( .ip1(n10637), .ip2(n10534), .op(n10618) );
  nor2_1 U10726 ( .ip1(n10536), .ip2(n10535), .op(n10537) );
  nor2_1 U10727 ( .ip1(n10538), .ip2(n10537), .op(n10617) );
  and2_1 U10728 ( .ip1(n10540), .ip2(n10539), .op(n10589) );
  nor2_1 U10729 ( .ip1(n10812), .ip2(n12156), .op(n10541) );
  or2_1 U10730 ( .ip1(m1Inputs[23]), .ip2(n10541), .op(n10543) );
  or2_1 U10731 ( .ip1(n14838), .ip2(n10541), .op(n10542) );
  nand2_1 U10732 ( .ip1(n10543), .ip2(n10542), .op(n10587) );
  nor2_1 U10733 ( .ip1(n10589), .ip2(n10587), .op(n10544) );
  nand2_1 U10734 ( .ip1(m1Inputs[18]), .ip2(n15028), .op(n10586) );
  xor2_1 U10735 ( .ip1(n10544), .ip2(n10586), .op(n10616) );
  nand2_1 U10736 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[30]), .op(
        n10915) );
  nor2_1 U10737 ( .ip1(n10545), .ip2(n10915), .op(n10641) );
  nor2_1 U10738 ( .ip1(n13801), .ip2(n10751), .op(n10546) );
  or2_1 U10739 ( .ip1(m1Inputs[30]), .ip2(n10546), .op(n10548) );
  or2_1 U10740 ( .ip1(n13803), .ip2(n10546), .op(n10547) );
  nand2_1 U10741 ( .ip1(n10548), .ip2(n10547), .op(n10640) );
  nand2_1 U10742 ( .ip1(m1Inputs[16]), .ip2(n14816), .op(n10642) );
  nor2_1 U10743 ( .ip1(n10640), .ip2(n10642), .op(n10549) );
  nor2_1 U10744 ( .ip1(n10641), .ip2(n10549), .op(n10621) );
  nor2_1 U10745 ( .ip1(n10551), .ip2(n10550), .op(n10552) );
  nor2_1 U10746 ( .ip1(n10553), .ip2(n10552), .op(n10620) );
  nand2_1 U10747 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[29]), .op(
        n10556) );
  nor3_1 U10748 ( .ip1(n10555), .ip2(n10828), .ip3(n10554), .op(n10592) );
  or2_1 U10749 ( .ip1(n10556), .ip2(n10592), .op(n10559) );
  nand2_1 U10750 ( .ip1(n12809), .ip2(m1Inputs[30]), .op(n10557) );
  or2_1 U10751 ( .ip1(n10557), .ip2(n10592), .op(n10558) );
  nand2_1 U10752 ( .ip1(n10559), .ip2(n10558), .op(n10590) );
  nand2_1 U10753 ( .ip1(column[23]), .ip2(n13859), .op(n10591) );
  xor2_1 U10754 ( .ip1(n10590), .ip2(n10591), .op(n10619) );
  fulladder U10755 ( .a(n10562), .b(n10561), .ci(n10560), .co(n10514), .s(
        n10664) );
  or2_1 U10756 ( .ip1(n10563), .ip2(n10564), .op(n10567) );
  or2_1 U10757 ( .ip1(n10565), .ip2(n10564), .op(n10566) );
  nand2_1 U10758 ( .ip1(n10567), .ip2(n10566), .op(n10649) );
  or2_1 U10759 ( .ip1(n10568), .ip2(n10569), .op(n10572) );
  or2_1 U10760 ( .ip1(n10570), .ip2(n10569), .op(n10571) );
  nand2_1 U10761 ( .ip1(n10572), .ip2(n10571), .op(n10648) );
  xor2_1 U10762 ( .ip1(n10574), .ip2(n10573), .op(n10647) );
  nor2_1 U10763 ( .ip1(n10576), .ip2(n10575), .op(n10577) );
  nor2_1 U10764 ( .ip1(n10578), .ip2(n10577), .op(n10646) );
  or2_1 U10765 ( .ip1(n10579), .ip2(n10581), .op(n10584) );
  inv_1 U10766 ( .ip(n10580), .op(n10582) );
  or2_1 U10767 ( .ip1(n10582), .ip2(n10581), .op(n10583) );
  nand2_1 U10768 ( .ip1(n10584), .ip2(n10583), .op(n10645) );
  nand2_1 U10769 ( .ip1(m1Inputs[19]), .ip2(n13718), .op(n10644) );
  nand2_1 U10770 ( .ip1(m1Inputs[29]), .ip2(n11974), .op(n10862) );
  nor2_1 U10771 ( .ip1(n10585), .ip2(n14853), .op(n10861) );
  nand2_1 U10772 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[25]), .op(
        n10860) );
  nor2_1 U10773 ( .ip1(n6745), .ip2(n10738), .op(n10916) );
  nand2_1 U10774 ( .ip1(m1Inputs[19]), .ip2(n14816), .op(n10914) );
  nor2_1 U10775 ( .ip1(n10587), .ip2(n10586), .op(n10588) );
  nor2_1 U10776 ( .ip1(n10589), .ip2(n10588), .op(n10615) );
  or2_1 U10777 ( .ip1(n10590), .ip2(n10592), .op(n10595) );
  inv_1 U10778 ( .ip(n10591), .op(n10593) );
  or2_1 U10779 ( .ip1(n10593), .ip2(n10592), .op(n10594) );
  nand2_1 U10780 ( .ip1(n10595), .ip2(n10594), .op(n10614) );
  nand2_1 U10781 ( .ip1(n15025), .ip2(m1Inputs[20]), .op(n10613) );
  fulladder U10782 ( .a(n10598), .b(n10597), .ci(n10596), .co(n10606), .s(
        n10631) );
  fulladder U10783 ( .a(n10601), .b(n10600), .ci(n10599), .co(n10608), .s(
        n10602) );
  inv_1 U10784 ( .ip(n10602), .op(n10630) );
  xor2_1 U10785 ( .ip1(n10604), .ip2(n10603), .op(n10629) );
  fulladder U10786 ( .a(n10607), .b(n10606), .ci(n10605), .co(n10464), .s(
        n10623) );
  fulladder U10787 ( .a(n10610), .b(n10609), .ci(n10608), .co(n10947), .s(
        n10611) );
  inv_1 U10788 ( .ip(n10611), .op(n10622) );
  inv_1 U10789 ( .ip(n10612), .op(n10967) );
  fulladder U10790 ( .a(n10615), .b(n10614), .ci(n10613), .co(n10936), .s(
        n10628) );
  fulladder U10791 ( .a(n10618), .b(n10617), .ci(n10616), .co(n10627), .s(
        n10667) );
  fulladder U10792 ( .a(n10621), .b(n10620), .ci(n10619), .co(n10626), .s(
        n10666) );
  fulladder U10793 ( .a(n10624), .b(n10623), .ci(n10622), .co(n10612), .s(
        n10625) );
  inv_1 U10794 ( .ip(n10625), .op(n10660) );
  fulladder U10795 ( .a(n10628), .b(n10627), .ci(n10626), .co(n10966), .s(
        n10659) );
  fulladder U10796 ( .a(n10631), .b(n10630), .ci(n10629), .co(n10624), .s(
        n10632) );
  inv_1 U10797 ( .ip(n10632), .op(n10684) );
  fulladder U10798 ( .a(n10635), .b(n10634), .ci(n10633), .co(n10676), .s(
        n10692) );
  nor2_1 U10799 ( .ip1(n10637), .ip2(n10636), .op(n10639) );
  xor2_1 U10800 ( .ip1(n10639), .ip2(n10638), .op(n10675) );
  nor2_1 U10801 ( .ip1(n10641), .ip2(n10640), .op(n10643) );
  xor2_1 U10802 ( .ip1(n10643), .ip2(n10642), .op(n10674) );
  fulladder U10803 ( .a(n10646), .b(n10645), .ci(n10644), .co(n10662), .s(
        n10691) );
  fulladder U10804 ( .a(n10649), .b(n10648), .ci(n10647), .co(n10663), .s(
        n10690) );
  fulladder U10805 ( .a(n10652), .b(n10651), .ci(n10650), .co(n10689), .s(
        n10694) );
  inv_1 U10806 ( .ip(n10653), .op(n10986) );
  fulladder U10807 ( .a(n10656), .b(n10655), .ci(n10654), .co(n10978), .s(
        n10657) );
  inv_1 U10808 ( .ip(n10657), .op(n10724) );
  fulladder U10809 ( .a(n10660), .b(n10659), .ci(n10658), .co(n10988), .s(
        n10661) );
  inv_1 U10810 ( .ip(n10661), .op(n10723) );
  fulladder U10811 ( .a(n10664), .b(n10663), .ci(n10662), .co(n10654), .s(
        n10665) );
  inv_1 U10812 ( .ip(n10665), .op(n10687) );
  fulladder U10813 ( .a(n10668), .b(n10667), .ci(n10666), .co(n10655), .s(
        n10669) );
  inv_1 U10814 ( .ip(n10669), .op(n10686) );
  fulladder U10815 ( .a(n10672), .b(n10671), .ci(n10670), .co(n10668), .s(
        n10673) );
  inv_1 U10816 ( .ip(n10673), .op(n10703) );
  fulladder U10817 ( .a(n10676), .b(n10675), .ci(n10674), .co(n10683), .s(
        n10677) );
  inv_1 U10818 ( .ip(n10677), .op(n10702) );
  fulladder U10819 ( .a(n10680), .b(n10679), .ci(n10678), .co(n10701), .s(
        n6519) );
  inv_1 U10820 ( .ip(n10681), .op(n11010) );
  fulladder U10821 ( .a(n10684), .b(n10683), .ci(n10682), .co(n10658), .s(
        n10700) );
  fulladder U10822 ( .a(n10687), .b(n10686), .ci(n10685), .co(n10722), .s(
        n10688) );
  inv_1 U10823 ( .ip(n10688), .op(n10699) );
  fulladder U10824 ( .a(n10691), .b(n10690), .ci(n10689), .co(n10682), .s(
        n10707) );
  fulladder U10825 ( .a(n10694), .b(n10693), .ci(n10692), .co(n10706), .s(
        n10720) );
  fulladder U10826 ( .a(n10697), .b(n10696), .ci(n10695), .co(n10705), .s(
        n10710) );
  fulladder U10827 ( .a(n10700), .b(n10699), .ci(n10698), .co(n11009), .s(
        n11014) );
  fulladder U10828 ( .a(n10703), .b(n10702), .ci(n10701), .co(n10685), .s(
        n10704) );
  inv_1 U10829 ( .ip(n10704), .op(n10713) );
  fulladder U10830 ( .a(n10707), .b(n10706), .ci(n10705), .co(n10698), .s(
        n10712) );
  fulladder U10831 ( .a(n10710), .b(n10709), .ci(n10708), .co(n10711), .s(
        n10719) );
  fulladder U10832 ( .a(n10713), .b(n10712), .ci(n10711), .co(n11013), .s(
        n11018) );
  fulladder U10833 ( .a(n10716), .b(n10715), .ci(n10714), .co(n10717), .s(
        \STAGE_1/M2/sum [5]) );
  inv_1 U10834 ( .ip(n10717), .op(n11017) );
  fulladder U10835 ( .a(n10720), .b(n10719), .ci(n10718), .co(n11016), .s(
        n6652) );
  inv_1 U10836 ( .ip(n10721), .op(n10985) );
  fulladder U10837 ( .a(n10724), .b(n10723), .ci(n10722), .co(n10984), .s(
        n10681) );
  nor2_1 U10838 ( .ip1(n14842), .ip2(n10734), .op(n10826) );
  nor2_1 U10839 ( .ip1(n14373), .ip2(n10812), .op(n10825) );
  nand4_1 U10840 ( .ip1(\STAGE_1/weightReg [10]), .ip2(n14994), .ip3(
        m1Inputs[27]), .ip4(m1Inputs[26]), .op(n10730) );
  nand2_1 U10841 ( .ip1(n14629), .ip2(m1Inputs[26]), .op(n10772) );
  inv_1 U10842 ( .ip(n10730), .op(n10725) );
  or2_1 U10843 ( .ip1(n10772), .ip2(n10725), .op(n10728) );
  nand2_1 U10844 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[27]), .op(
        n10726) );
  or2_1 U10845 ( .ip1(n10726), .ip2(n10725), .op(n10727) );
  nand2_1 U10846 ( .ip1(n10728), .ip2(n10727), .op(n10749) );
  nand3_1 U10847 ( .ip1(column[28]), .ip2(n15042), .ip3(n10749), .op(n10729)
         );
  nand2_1 U10848 ( .ip1(n10730), .ip2(n10729), .op(n10824) );
  nand2_1 U10849 ( .ip1(m1Inputs[23]), .ip2(n15028), .op(n10732) );
  nand2_1 U10850 ( .ip1(m1Inputs[25]), .ip2(n14847), .op(n10731) );
  xor2_1 U10851 ( .ip1(n10732), .ip2(n10731), .op(n10754) );
  nand2_1 U10852 ( .ip1(n14816), .ip2(m1Inputs[22]), .op(n10733) );
  xor2_1 U10853 ( .ip1(n10754), .ip2(n10733), .op(n10849) );
  nor2_1 U10854 ( .ip1(n14902), .ip2(n10812), .op(n10765) );
  and2_1 U10855 ( .ip1(n10778), .ip2(n10765), .op(n10737) );
  nand2_1 U10856 ( .ip1(m1Inputs[24]), .ip2(n14847), .op(n10736) );
  nor2_1 U10857 ( .ip1(n14902), .ip2(n10734), .op(n10735) );
  xor2_1 U10858 ( .ip1(n10736), .ip2(n10735), .op(n10786) );
  nor3_1 U10859 ( .ip1(n14842), .ip2(n10866), .ip3(n10786), .op(n10787) );
  nor2_1 U10860 ( .ip1(n10737), .ip2(n10787), .op(n10848) );
  nand2_1 U10861 ( .ip1(m1Inputs[28]), .ip2(\STAGE_1/weightReg [7]), .op(
        n10793) );
  nor2_1 U10862 ( .ip1(n10738), .ip2(n14783), .op(n10792) );
  nand2_1 U10863 ( .ip1(m1Inputs[30]), .ip2(n12699), .op(n10791) );
  inv_1 U10864 ( .ip(n10739), .op(n10833) );
  nor2_1 U10865 ( .ip1(n12083), .ip2(n10753), .op(n10893) );
  inv_1 U10866 ( .ip(n10893), .op(n10740) );
  nor2_1 U10867 ( .ip1(n10772), .ip2(n10740), .op(n10742) );
  inv_1 U10868 ( .ip(n10742), .op(n10747) );
  nand2_1 U10869 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[26]), .op(
        n10741) );
  or2_1 U10870 ( .ip1(n10741), .ip2(n10742), .op(n10745) );
  nand2_1 U10871 ( .ip1(n14629), .ip2(m1Inputs[25]), .op(n10743) );
  or2_1 U10872 ( .ip1(n10743), .ip2(n10742), .op(n10744) );
  nand2_1 U10873 ( .ip1(n10745), .ip2(n10744), .op(n10799) );
  nand3_1 U10874 ( .ip1(column[27]), .ip2(n15042), .ip3(n10799), .op(n10746)
         );
  nand2_1 U10875 ( .ip1(n10747), .ip2(n10746), .op(n10785) );
  inv_1 U10876 ( .ip(n10749), .op(n10750) );
  nand2_1 U10877 ( .ip1(column[28]), .ip2(n13859), .op(n10748) );
  mux2_1 U10878 ( .ip1(n10750), .ip2(n10749), .s(n10748), .op(n10784) );
  nor2_1 U10879 ( .ip1(n10813), .ip2(n14289), .op(n10797) );
  nor2_1 U10880 ( .ip1(n6503), .ip2(n10751), .op(n10796) );
  nand2_1 U10881 ( .ip1(n14976), .ip2(m1Inputs[20]), .op(n10795) );
  nor2_1 U10882 ( .ip1(n12083), .ip2(n11033), .op(n10820) );
  nor2_1 U10883 ( .ip1(n10828), .ip2(n14384), .op(n10819) );
  nand2_1 U10884 ( .ip1(n14976), .ip2(m1Inputs[22]), .op(n10818) );
  nor2_1 U10885 ( .ip1(n14902), .ip2(n10753), .op(n10804) );
  nor2_1 U10886 ( .ip1(n6503), .ip2(n10813), .op(n10803) );
  nand2_1 U10887 ( .ip1(m1Inputs[31]), .ip2(n13749), .op(n10802) );
  nor2_1 U10888 ( .ip1(n10828), .ip2(n14836), .op(n10770) );
  nor2_1 U10889 ( .ip1(n6503), .ip2(n11033), .op(n10769) );
  nand2_1 U10890 ( .ip1(m1Inputs[31]), .ip2(n12699), .op(n10768) );
  inv_1 U10891 ( .ip(n10752), .op(n10838) );
  nor2_1 U10892 ( .ip1(n14340), .ip2(n10753), .op(n11027) );
  nand2_1 U10893 ( .ip1(n10778), .ip2(n11027), .op(n10756) );
  nand3_1 U10894 ( .ip1(n14816), .ip2(m1Inputs[22]), .ip3(n10754), .op(n10755)
         );
  nand2_1 U10895 ( .ip1(n10756), .ip2(n10755), .op(n10831) );
  nand2_1 U10896 ( .ip1(n14629), .ip2(m1Inputs[27]), .op(n10757) );
  nand2_1 U10897 ( .ip1(n13718), .ip2(m1Inputs[27]), .op(n10805) );
  nor2_1 U10898 ( .ip1(n10805), .ip2(n10772), .op(n10814) );
  or2_1 U10899 ( .ip1(n10757), .ip2(n10814), .op(n10760) );
  nand2_1 U10900 ( .ip1(n14847), .ip2(m1Inputs[26]), .op(n10758) );
  or2_1 U10901 ( .ip1(n10758), .ip2(n10814), .op(n10759) );
  nand2_1 U10902 ( .ip1(n10760), .ip2(n10759), .op(n10815) );
  inv_1 U10903 ( .ip(n10815), .op(n10762) );
  nand2_1 U10904 ( .ip1(column[29]), .ip2(n13859), .op(n10761) );
  mux2_1 U10905 ( .ip1(n10762), .ip2(n10815), .s(n10761), .op(n10830) );
  nor2_1 U10906 ( .ip1(n10813), .ip2(n12156), .op(n10766) );
  nand2_1 U10907 ( .ip1(\STAGE_1/weightReg [15]), .ip2(m1Inputs[21]), .op(
        n10764) );
  inv_1 U10908 ( .ip(n10763), .op(n10837) );
  fulladder U10909 ( .a(n10766), .b(n10765), .ci(n10764), .co(n10829), .s(
        n10767) );
  inv_1 U10910 ( .ip(n10767), .op(n10845) );
  fulladder U10911 ( .a(n10770), .b(n10769), .ci(n10768), .co(n10821), .s(
        n10771) );
  inv_1 U10912 ( .ip(n10771), .op(n10844) );
  nor3_1 U10913 ( .ip1(n6503), .ip2(n10812), .ip3(n10772), .op(n10776) );
  nand2_1 U10914 ( .ip1(m1Inputs[26]), .ip2(n14975), .op(n10774) );
  nand2_1 U10915 ( .ip1(m1Inputs[24]), .ip2(\STAGE_1/weightReg [10]), .op(
        n10773) );
  xor2_1 U10916 ( .ip1(n10774), .ip2(n10773), .op(n10864) );
  and3_1 U10917 ( .ip1(column[26]), .ip2(n15042), .ip3(n10864), .op(n10775) );
  nor2_1 U10918 ( .ip1(n10776), .ip2(n10775), .op(n10853) );
  nand2_1 U10919 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[22]), .op(
        n10852) );
  nor3_1 U10920 ( .ip1(n14824), .ip2(n11033), .ip3(n10777), .op(n10908) );
  or2_1 U10921 ( .ip1(n13749), .ip2(n10778), .op(n10780) );
  or2_1 U10922 ( .ip1(m1Inputs[28]), .ip2(n10778), .op(n10779) );
  nand2_1 U10923 ( .ip1(n10780), .ip2(n10779), .op(n10907) );
  nand2_1 U10924 ( .ip1(n14816), .ip2(m1Inputs[20]), .op(n10909) );
  nor2_1 U10925 ( .ip1(n10907), .ip2(n10909), .op(n10781) );
  nor2_1 U10926 ( .ip1(n10908), .ip2(n10781), .op(n10851) );
  inv_1 U10927 ( .ip(n10782), .op(n10840) );
  fulladder U10928 ( .a(n10785), .b(n10784), .ci(n10783), .co(n10832), .s(
        n10874) );
  or2_1 U10929 ( .ip1(n10786), .ip2(n10787), .op(n10790) );
  nand2_1 U10930 ( .ip1(n14816), .ip2(m1Inputs[21]), .op(n10788) );
  or2_1 U10931 ( .ip1(n10788), .ip2(n10787), .op(n10789) );
  nand2_1 U10932 ( .ip1(n10790), .ip2(n10789), .op(n10905) );
  fulladder U10933 ( .a(n10793), .b(n10792), .ci(n10791), .co(n10847), .s(
        n10794) );
  inv_1 U10934 ( .ip(n10794), .op(n10904) );
  fulladder U10935 ( .a(n10797), .b(n10796), .ci(n10795), .co(n10783), .s(
        n10903) );
  inv_1 U10936 ( .ip(n10799), .op(n10800) );
  nand2_1 U10937 ( .ip1(column[27]), .ip2(n13859), .op(n10798) );
  mux2_1 U10938 ( .ip1(n10800), .ip2(n10799), .s(n10798), .op(n10901) );
  nor2_1 U10939 ( .ip1(n10828), .ip2(n14783), .op(n10890) );
  nand2_1 U10940 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[31]), .op(
        n10889) );
  nor2_1 U10941 ( .ip1(n10813), .ip2(n12746), .op(n10894) );
  nand2_1 U10942 ( .ip1(m1Inputs[19]), .ip2(n14976), .op(n10892) );
  inv_1 U10943 ( .ip(n10801), .op(n11044) );
  fulladder U10944 ( .a(n10804), .b(n10803), .ci(n10802), .co(n11070), .s(
        n10822) );
  nand4_1 U10945 ( .ip1(\STAGE_1/weightReg [11]), .ip2(\STAGE_1/weightReg [10]), .ip3(m1Inputs[28]), .ip4(m1Inputs[27]), .op(n11021) );
  inv_1 U10946 ( .ip(n11021), .op(n10806) );
  or2_1 U10947 ( .ip1(n10805), .ip2(n10806), .op(n10809) );
  nand2_1 U10948 ( .ip1(n14629), .ip2(m1Inputs[28]), .op(n10807) );
  or2_1 U10949 ( .ip1(n10807), .ip2(n10806), .op(n10808) );
  nand2_1 U10950 ( .ip1(n10809), .ip2(n10808), .op(n11020) );
  inv_1 U10951 ( .ip(n11020), .op(n10811) );
  nand2_1 U10952 ( .ip1(column[30]), .ip2(n13039), .op(n10810) );
  mux2_1 U10953 ( .ip1(n10811), .ip2(n11020), .s(n10810), .op(n11069) );
  nor2_1 U10954 ( .ip1(n14842), .ip2(n10812), .op(n11047) );
  nor2_1 U10955 ( .ip1(n12083), .ip2(n10813), .op(n11046) );
  nand2_1 U10956 ( .ip1(m1Inputs[31]), .ip2(n4627), .op(n11045) );
  inv_1 U10957 ( .ip(n10814), .op(n10817) );
  nand3_1 U10958 ( .ip1(column[29]), .ip2(n15042), .ip3(n10815), .op(n10816)
         );
  nand2_1 U10959 ( .ip1(n10817), .ip2(n10816), .op(n11026) );
  fulladder U10960 ( .a(n10820), .b(n10819), .ci(n10818), .co(n11025), .s(
        n10823) );
  fulladder U10961 ( .a(n10823), .b(n10822), .ci(n10821), .co(n11034), .s(
        n10752) );
  fulladder U10962 ( .a(n10826), .b(n10825), .ci(n10824), .co(n11030), .s(
        n10834) );
  nor2_1 U10963 ( .ip1(n14902), .ip2(n10827), .op(n11039) );
  nor2_1 U10964 ( .ip1(n6503), .ip2(n10828), .op(n11038) );
  nand2_1 U10965 ( .ip1(n14976), .ip2(m1Inputs[23]), .op(n11037) );
  fulladder U10966 ( .a(n10831), .b(n10830), .ci(n10829), .co(n11028), .s(
        n10763) );
  fulladder U10967 ( .a(n10834), .b(n10833), .ci(n10832), .co(n11073), .s(
        n10841) );
  inv_1 U10968 ( .ip(n10835), .op(n11043) );
  fulladder U10969 ( .a(n10838), .b(n10837), .ci(n10836), .co(n11042), .s(
        n10782) );
  fulladder U10970 ( .a(n10841), .b(n10840), .ci(n10839), .co(n10801), .s(
        n10842) );
  inv_1 U10971 ( .ip(n10842), .op(n10919) );
  fulladder U10972 ( .a(n10845), .b(n10844), .ci(n10843), .co(n10836), .s(
        n10846) );
  inv_1 U10973 ( .ip(n10846), .op(n10922) );
  fulladder U10974 ( .a(n10849), .b(n10848), .ci(n10847), .co(n10739), .s(
        n10850) );
  inv_1 U10975 ( .ip(n10850), .op(n10921) );
  fulladder U10976 ( .a(n10853), .b(n10852), .ci(n10851), .co(n10843), .s(
        n10854) );
  inv_1 U10977 ( .ip(n10854), .op(n10878) );
  or2_1 U10978 ( .ip1(n10855), .ip2(n10856), .op(n10859) );
  or2_1 U10979 ( .ip1(n10857), .ip2(n10856), .op(n10858) );
  nand2_1 U10980 ( .ip1(n10859), .ip2(n10858), .op(n10932) );
  fulladder U10981 ( .a(n10862), .b(n10861), .ci(n10860), .co(n10931), .s(
        n10938) );
  nand2_1 U10982 ( .ip1(column[26]), .ip2(n13859), .op(n10863) );
  xor2_1 U10983 ( .ip1(n10864), .ip2(n10863), .op(n10930) );
  inv_1 U10984 ( .ip(n10865), .op(n10877) );
  nor2_1 U10985 ( .ip1(n14340), .ip2(n10866), .op(n10881) );
  nor2_1 U10986 ( .ip1(n14902), .ip2(n10867), .op(n10880) );
  fulladder U10987 ( .a(n10870), .b(n10869), .ci(n10868), .co(n10879), .s(
        n10483) );
  inv_1 U10988 ( .ip(n10871), .op(n10918) );
  fulladder U10989 ( .a(n10874), .b(n10873), .ci(n10872), .co(n10839), .s(
        n10875) );
  inv_1 U10990 ( .ip(n10875), .op(n10926) );
  fulladder U10991 ( .a(n10878), .b(n10877), .ci(n10876), .co(n10920), .s(
        n10958) );
  fulladder U10992 ( .a(n10881), .b(n10880), .ci(n10879), .co(n10876), .s(
        n10945) );
  fulladder U10993 ( .a(n10884), .b(n10883), .ci(n10882), .co(n10885), .s(
        n10962) );
  inv_1 U10994 ( .ip(n10885), .op(n10944) );
  fulladder U10995 ( .a(n10888), .b(n10887), .ci(n10886), .co(n10943), .s(
        n10498) );
  fulladder U10996 ( .a(n10891), .b(n10890), .ci(n10889), .co(n10900), .s(
        n10941) );
  fulladder U10997 ( .a(n10894), .b(n10893), .ci(n10892), .co(n10899), .s(
        n10940) );
  fulladder U10998 ( .a(n10897), .b(n10896), .ci(n10895), .co(n10939), .s(
        n10455) );
  inv_1 U10999 ( .ip(n10898), .op(n10925) );
  fulladder U11000 ( .a(n10901), .b(n10900), .ci(n10899), .co(n10872), .s(
        n10902) );
  inv_1 U11001 ( .ip(n10902), .op(n10929) );
  fulladder U11002 ( .a(n10905), .b(n10904), .ci(n10903), .co(n10873), .s(
        n10906) );
  inv_1 U11003 ( .ip(n10906), .op(n10928) );
  nor2_1 U11004 ( .ip1(n10908), .ip2(n10907), .op(n10910) );
  xor2_1 U11005 ( .ip1(n10910), .ip2(n10909), .op(n10935) );
  inv_1 U11006 ( .ip(n10911), .op(n10913) );
  nor2_1 U11007 ( .ip1(n10913), .ip2(n10912), .op(n10934) );
  fulladder U11008 ( .a(n10916), .b(n10915), .ci(n10914), .co(n10933), .s(
        n10937) );
  fulladder U11009 ( .a(n10919), .b(n10918), .ci(n10917), .co(n11077), .s(
        n10994) );
  fulladder U11010 ( .a(n10922), .b(n10921), .ci(n10920), .co(n10871), .s(
        n10923) );
  inv_1 U11011 ( .ip(n10923), .op(n10952) );
  fulladder U11012 ( .a(n10926), .b(n10925), .ci(n10924), .co(n10917), .s(
        n10951) );
  fulladder U11013 ( .a(n10929), .b(n10928), .ci(n10927), .co(n10924), .s(
        n10955) );
  fulladder U11014 ( .a(n10932), .b(n10931), .ci(n10930), .co(n10865), .s(
        n10965) );
  fulladder U11015 ( .a(n10935), .b(n10934), .ci(n10933), .co(n10927), .s(
        n10964) );
  fulladder U11016 ( .a(n10938), .b(n10937), .ci(n10936), .co(n10963), .s(
        n10968) );
  fulladder U11017 ( .a(n10941), .b(n10940), .ci(n10939), .co(n10956), .s(
        n10942) );
  inv_1 U11018 ( .ip(n10942), .op(n10974) );
  fulladder U11019 ( .a(n10945), .b(n10944), .ci(n10943), .co(n10957), .s(
        n10946) );
  inv_1 U11020 ( .ip(n10946), .op(n10973) );
  fulladder U11021 ( .a(n10949), .b(n10948), .ci(n10947), .co(n10972), .s(
        n10980) );
  fulladder U11022 ( .a(n10952), .b(n10951), .ci(n10950), .co(n10993), .s(
        n10998) );
  fulladder U11023 ( .a(n10955), .b(n10954), .ci(n10953), .co(n10950), .s(
        n10971) );
  fulladder U11024 ( .a(n10958), .b(n10957), .ci(n10956), .co(n10898), .s(
        n10959) );
  inv_1 U11025 ( .ip(n10959), .op(n10970) );
  fulladder U11026 ( .a(n10962), .b(n10961), .ci(n10960), .co(n10977), .s(
        n10979) );
  fulladder U11027 ( .a(n10965), .b(n10964), .ci(n10963), .co(n10954), .s(
        n10976) );
  fulladder U11028 ( .a(n10968), .b(n10967), .ci(n10966), .co(n10975), .s(
        n10989) );
  fulladder U11029 ( .a(n10971), .b(n10970), .ci(n10969), .co(n10997), .s(
        n11002) );
  fulladder U11030 ( .a(n10974), .b(n10973), .ci(n10972), .co(n10953), .s(
        n10983) );
  fulladder U11031 ( .a(n10977), .b(n10976), .ci(n10975), .co(n10969), .s(
        n10982) );
  fulladder U11032 ( .a(n10980), .b(n10979), .ci(n10978), .co(n10981), .s(
        n10990) );
  fulladder U11033 ( .a(n10983), .b(n10982), .ci(n10981), .co(n11001), .s(
        n11006) );
  fulladder U11034 ( .a(n10986), .b(n10985), .ci(n10984), .co(n10987), .s(
        \STAGE_1/M2/sum [9]) );
  inv_1 U11035 ( .ip(n10987), .op(n11005) );
  fulladder U11036 ( .a(n10990), .b(n10989), .ci(n10988), .co(n11004), .s(
        n10653) );
  inv_1 U11037 ( .ip(n10991), .op(\STAGE_1/M2/sum [14]) );
  fulladder U11038 ( .a(n10994), .b(n10993), .ci(n10992), .co(n11076), .s(
        n10995) );
  inv_1 U11039 ( .ip(n10995), .op(\STAGE_1/M2/sum [13]) );
  fulladder U11040 ( .a(n10998), .b(n10997), .ci(n10996), .co(n10992), .s(
        n10999) );
  inv_1 U11041 ( .ip(n10999), .op(\STAGE_1/M2/sum [12]) );
  fulladder U11042 ( .a(n11002), .b(n11001), .ci(n11000), .co(n10996), .s(
        n11003) );
  inv_1 U11043 ( .ip(n11003), .op(\STAGE_1/M2/sum [11]) );
  fulladder U11044 ( .a(n11006), .b(n11005), .ci(n11004), .co(n11000), .s(
        n11007) );
  inv_1 U11045 ( .ip(n11007), .op(\STAGE_1/M2/sum [10]) );
  fulladder U11046 ( .a(n11010), .b(n11009), .ci(n11008), .co(n10721), .s(
        n11011) );
  inv_1 U11047 ( .ip(n11011), .op(\STAGE_1/M2/sum [8]) );
  fulladder U11048 ( .a(n11014), .b(n11013), .ci(n11012), .co(n11008), .s(
        n11015) );
  inv_1 U11049 ( .ip(n11015), .op(\STAGE_1/M2/sum [7]) );
  fulladder U11050 ( .a(n11018), .b(n11017), .ci(n11016), .co(n11012), .s(
        n11019) );
  inv_1 U11051 ( .ip(n11019), .op(\STAGE_1/M2/sum [6]) );
  nand2_1 U11052 ( .ip1(column[31]), .ip2(n13039), .op(n11024) );
  nand3_1 U11053 ( .ip1(column[30]), .ip2(n15042), .ip3(n11020), .op(n11022)
         );
  nand2_1 U11054 ( .ip1(n11022), .ip2(n11021), .op(n11023) );
  xor2_1 U11055 ( .ip1(n11024), .ip2(n11023), .op(n11057) );
  fulladder U11056 ( .a(n11027), .b(n11026), .ci(n11025), .co(n11032), .s(
        n11035) );
  fulladder U11057 ( .a(n11030), .b(n11029), .ci(n11028), .co(n11031), .s(
        n11074) );
  xor2_1 U11058 ( .ip1(n11032), .ip2(n11031), .op(n11055) );
  nor2_1 U11059 ( .ip1(n14824), .ip2(n11033), .op(n11053) );
  fulladder U11060 ( .a(n11036), .b(n11035), .ci(n11034), .co(n11041), .s(
        n11075) );
  fulladder U11061 ( .a(n11039), .b(n11038), .ci(n11037), .co(n11040), .s(
        n11029) );
  xor2_1 U11062 ( .ip1(n11041), .ip2(n11040), .op(n11051) );
  fulladder U11063 ( .a(n11044), .b(n11043), .ci(n11042), .co(n11049), .s(
        n11078) );
  fulladder U11064 ( .a(n11047), .b(n11046), .ci(n11045), .co(n11048), .s(
        n11068) );
  xor2_1 U11065 ( .ip1(n11049), .ip2(n11048), .op(n11050) );
  xor2_1 U11066 ( .ip1(n11051), .ip2(n11050), .op(n11052) );
  xor2_1 U11067 ( .ip1(n11053), .ip2(n11052), .op(n11054) );
  xor2_1 U11068 ( .ip1(n11055), .ip2(n11054), .op(n11056) );
  xor2_1 U11069 ( .ip1(n11057), .ip2(n11056), .op(n11065) );
  nand2_1 U11070 ( .ip1(m1Inputs[26]), .ip2(n15028), .op(n11059) );
  nand2_1 U11071 ( .ip1(m1Inputs[29]), .ip2(n14629), .op(n11058) );
  xor2_1 U11072 ( .ip1(n11059), .ip2(n11058), .op(n11063) );
  nand2_1 U11073 ( .ip1(m1Inputs[30]), .ip2(n14994), .op(n11061) );
  nand2_1 U11074 ( .ip1(m1Inputs[31]), .ip2(n14975), .op(n11060) );
  xor2_1 U11075 ( .ip1(n11061), .ip2(n11060), .op(n11062) );
  xor2_1 U11076 ( .ip1(n11063), .ip2(n11062), .op(n11064) );
  xor2_1 U11077 ( .ip1(n11065), .ip2(n11064), .op(n11086) );
  nand2_1 U11078 ( .ip1(m1Inputs[24]), .ip2(n14976), .op(n11067) );
  nand2_1 U11079 ( .ip1(m1Inputs[25]), .ip2(n14816), .op(n11066) );
  xor2_1 U11080 ( .ip1(n11067), .ip2(n11066), .op(n11072) );
  fulladder U11081 ( .a(n11070), .b(n11069), .ci(n11068), .co(n11071), .s(
        n11036) );
  xor2_1 U11082 ( .ip1(n11072), .ip2(n11071), .op(n11082) );
  fulladder U11083 ( .a(n11075), .b(n11074), .ci(n11073), .co(n11080), .s(
        n10835) );
  fulladder U11084 ( .a(n11078), .b(n11077), .ci(n11076), .co(n11079), .s(
        n10991) );
  xor2_1 U11085 ( .ip1(n11080), .ip2(n11079), .op(n11081) );
  xor2_1 U11086 ( .ip1(n11082), .ip2(n11081), .op(n11084) );
  nand2_1 U11087 ( .ip1(m1Inputs[27]), .ip2(n15025), .op(n11083) );
  xor2_1 U11088 ( .ip1(n11084), .ip2(n11083), .op(n11085) );
  xor2_1 U11089 ( .ip1(n11086), .ip2(n11085), .op(\STAGE_1/M2/sum [15]) );
  or2_1 U11090 ( .ip1(n11087), .ip2(n11088), .op(n11091) );
  or2_1 U11091 ( .ip1(n11089), .ip2(n11088), .op(n11090) );
  nand2_1 U11092 ( .ip1(n11091), .ip2(n11090), .op(n11693) );
  or2_1 U11093 ( .ip1(n11092), .ip2(n11093), .op(n11096) );
  or2_1 U11094 ( .ip1(n11094), .ip2(n11093), .op(n11095) );
  nand2_1 U11095 ( .ip1(n11096), .ip2(n11095), .op(n11692) );
  nand2_1 U11096 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[42]), .op(
        n11098) );
  nor3_1 U11097 ( .ip1(n13709), .ip2(n11472), .ip3(n11097), .op(n11592) );
  or2_1 U11098 ( .ip1(n11098), .ip2(n11592), .op(n11100) );
  nand2_1 U11099 ( .ip1(n12809), .ip2(m1Inputs[43]), .op(n11560) );
  or2_1 U11100 ( .ip1(n11560), .ip2(n11592), .op(n11099) );
  nand2_1 U11101 ( .ip1(n11100), .ip2(n11099), .op(n11590) );
  nand2_1 U11102 ( .ip1(column[36]), .ip2(n13039), .op(n11591) );
  xor2_1 U11103 ( .ip1(n11590), .ip2(n11591), .op(n11691) );
  fulladder U11104 ( .a(n11103), .b(n11102), .ci(n11101), .co(n11104), .s(
        n6299) );
  inv_1 U11105 ( .ip(n11104), .op(n11714) );
  fulladder U11106 ( .a(n11107), .b(n11106), .ci(n11105), .co(n11713), .s(
        n11139) );
  or2_1 U11107 ( .ip1(n11108), .ip2(n11109), .op(n11112) );
  or2_1 U11108 ( .ip1(n11110), .ip2(n11109), .op(n11111) );
  nand2_1 U11109 ( .ip1(n11112), .ip2(n11111), .op(n11696) );
  nand2_1 U11110 ( .ip1(m1Inputs[39]), .ip2(n12699), .op(n11114) );
  nor3_1 U11111 ( .ip1(n11461), .ip2(n13835), .ip3(n11113), .op(n11618) );
  or2_1 U11112 ( .ip1(n11114), .ip2(n11618), .op(n11116) );
  nand2_1 U11113 ( .ip1(m1Inputs[40]), .ip2(n11974), .op(n11543) );
  or2_1 U11114 ( .ip1(n11543), .ip2(n11618), .op(n11115) );
  nand2_1 U11115 ( .ip1(n11116), .ip2(n11115), .op(n11617) );
  nor2_1 U11116 ( .ip1(n11549), .ip2(n13579), .op(n11619) );
  xnor2_1 U11117 ( .ip1(n11617), .ip2(n11619), .op(n11695) );
  nand2_1 U11118 ( .ip1(n14835), .ip2(m1Inputs[37]), .op(n11118) );
  nor3_1 U11119 ( .ip1(n11283), .ip2(n14384), .ip3(n11117), .op(n11597) );
  or2_1 U11120 ( .ip1(n11118), .ip2(n11597), .op(n11120) );
  nand2_1 U11121 ( .ip1(m1Inputs[38]), .ip2(n12981), .op(n11533) );
  or2_1 U11122 ( .ip1(n11533), .ip2(n11597), .op(n11119) );
  nand2_1 U11123 ( .ip1(n11120), .ip2(n11119), .op(n11596) );
  nor2_1 U11124 ( .ip1(n11539), .ip2(n13594), .op(n11598) );
  xnor2_1 U11125 ( .ip1(n11596), .ip2(n11598), .op(n11694) );
  fulladder U11126 ( .a(n11123), .b(n11122), .ci(n11121), .co(n11712), .s(
        n11136) );
  nand2_1 U11127 ( .ip1(n14975), .ip2(m1Inputs[36]), .op(n11690) );
  or2_1 U11128 ( .ip1(n11124), .ip2(n11126), .op(n11129) );
  inv_1 U11129 ( .ip(n11125), .op(n11127) );
  or2_1 U11130 ( .ip1(n11127), .ip2(n11126), .op(n11128) );
  nand2_1 U11131 ( .ip1(n11129), .ip2(n11128), .op(n11689) );
  nand2_1 U11132 ( .ip1(m1Inputs[35]), .ip2(n14994), .op(n11688) );
  nand2_1 U11133 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[44]), .op(
        n11440) );
  nor3_1 U11134 ( .ip1(n10476), .ip2(n11544), .ip3(n11440), .op(n11625) );
  nor2_1 U11135 ( .ip1(n13801), .ip2(n11544), .op(n11130) );
  or2_1 U11136 ( .ip1(m1Inputs[44]), .ip2(n11130), .op(n11132) );
  or2_1 U11137 ( .ip1(n13803), .ip2(n11130), .op(n11131) );
  nand2_1 U11138 ( .ip1(n11132), .ip2(n11131), .op(n11623) );
  nor2_1 U11139 ( .ip1(n11625), .ip2(n11623), .op(n11133) );
  nand2_1 U11140 ( .ip1(m1Inputs[32]), .ip2(n15025), .op(n11622) );
  xor2_1 U11141 ( .ip1(n11133), .ip2(n11622), .op(n11710) );
  fulladder U11142 ( .a(n11136), .b(n11135), .ci(n11134), .co(n11725), .s(
        n11143) );
  fulladder U11143 ( .a(n11139), .b(n11138), .ci(n11137), .co(n11735), .s(
        n11142) );
  inv_1 U11144 ( .ip(n11140), .op(n11733) );
  fulladder U11145 ( .a(n11143), .b(n11142), .ci(n11141), .co(n11144), .s(
        n6317) );
  inv_1 U11146 ( .ip(n11144), .op(n11732) );
  fulladder U11147 ( .a(n11147), .b(n11146), .ci(n11145), .co(n11731), .s(
        \STAGE_1/M3/sum [3]) );
  nand2_1 U11148 ( .ip1(m1Inputs[46]), .ip2(\STAGE_1/weightReg [7]), .op(
        n11231) );
  nor2_1 U11149 ( .ip1(n14853), .ip2(n11283), .op(n11230) );
  nand2_1 U11150 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[44]), .op(
        n11229) );
  nand2_1 U11151 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[45]), .op(
        n11224) );
  nand2_1 U11152 ( .ip1(n15025), .ip2(m1Inputs[41]), .op(n11223) );
  nand2_1 U11153 ( .ip1(m1Inputs[46]), .ip2(\STAGE_1/weightReg [6]), .op(
        n11161) );
  nand2_1 U11154 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[44]), .op(
        n11159) );
  nand2_1 U11155 ( .ip1(m1Inputs[39]), .ip2(\STAGE_1/weightReg [13]), .op(
        n11149) );
  nand2_1 U11156 ( .ip1(m1Inputs[41]), .ip2(n13718), .op(n11148) );
  xor2_1 U11157 ( .ip1(n11149), .ip2(n11148), .op(n11186) );
  nor2_1 U11158 ( .ip1(n14824), .ip2(n11534), .op(n11162) );
  inv_1 U11159 ( .ip(n11162), .op(n11181) );
  nand2_1 U11160 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[41]), .op(
        n11789) );
  nor2_1 U11161 ( .ip1(n11181), .ip2(n11789), .op(n11150) );
  or2_1 U11162 ( .ip1(n11186), .ip2(n11150), .op(n11152) );
  nor2_1 U11163 ( .ip1(n14842), .ip2(n11283), .op(n11185) );
  or2_1 U11164 ( .ip1(n11185), .ip2(n11150), .op(n11151) );
  nand2_1 U11165 ( .ip1(n11152), .ip2(n11151), .op(n11241) );
  nand2_1 U11166 ( .ip1(n14629), .ip2(m1Inputs[43]), .op(n11173) );
  nand2_1 U11167 ( .ip1(n13718), .ip2(m1Inputs[43]), .op(n11217) );
  nand2_1 U11168 ( .ip1(n14629), .ip2(m1Inputs[42]), .op(n11174) );
  nor2_1 U11169 ( .ip1(n11217), .ip2(n11174), .op(n11228) );
  or2_1 U11170 ( .ip1(n11173), .ip2(n11228), .op(n11155) );
  nand2_1 U11171 ( .ip1(n13718), .ip2(m1Inputs[42]), .op(n11153) );
  or2_1 U11172 ( .ip1(n11153), .ip2(n11228), .op(n11154) );
  nand2_1 U11173 ( .ip1(n11155), .ip2(n11154), .op(n11226) );
  nand2_1 U11174 ( .ip1(column[45]), .ip2(n13039), .op(n11156) );
  xor2_1 U11175 ( .ip1(n11226), .ip2(n11156), .op(n11240) );
  nor2_1 U11176 ( .ip1(n14853), .ip2(n11555), .op(n11158) );
  nand2_1 U11177 ( .ip1(n15025), .ip2(m1Inputs[40]), .op(n11180) );
  nand2_1 U11178 ( .ip1(m1Inputs[45]), .ip2(n4627), .op(n11157) );
  fulladder U11179 ( .a(n11158), .b(n11180), .ci(n11157), .co(n11239), .s(
        n11254) );
  fulladder U11180 ( .a(n11161), .b(n11160), .ci(n11159), .co(n11232), .s(
        n11253) );
  nand2_1 U11181 ( .ip1(n13718), .ip2(m1Inputs[44]), .op(n11810) );
  nand2_1 U11182 ( .ip1(m1Inputs[39]), .ip2(n12981), .op(n11536) );
  nor2_1 U11183 ( .ip1(n11810), .ip2(n11536), .op(n11280) );
  or2_1 U11184 ( .ip1(n13749), .ip2(n11162), .op(n11164) );
  or2_1 U11185 ( .ip1(m1Inputs[44]), .ip2(n11162), .op(n11163) );
  nand2_1 U11186 ( .ip1(n11164), .ip2(n11163), .op(n11279) );
  nand2_1 U11187 ( .ip1(n14816), .ip2(m1Inputs[36]), .op(n11281) );
  nor2_1 U11188 ( .ip1(n11279), .ip2(n11281), .op(n11165) );
  nor2_1 U11189 ( .ip1(n11280), .ip2(n11165), .op(n11258) );
  nand2_1 U11190 ( .ip1(m1Inputs[42]), .ip2(n14975), .op(n11167) );
  nand2_1 U11191 ( .ip1(m1Inputs[40]), .ip2(\STAGE_1/weightReg [10]), .op(
        n11166) );
  xor2_1 U11192 ( .ip1(n11167), .ip2(n11166), .op(n11266) );
  nor2_1 U11193 ( .ip1(n6503), .ip2(n11461), .op(n11423) );
  and3_1 U11194 ( .ip1(\STAGE_1/weightReg [10]), .ip2(m1Inputs[42]), .ip3(
        n11423), .op(n11168) );
  or2_1 U11195 ( .ip1(n11266), .ip2(n11168), .op(n11171) );
  nand2_1 U11196 ( .ip1(column[42]), .ip2(n13039), .op(n11265) );
  inv_1 U11197 ( .ip(n11265), .op(n11169) );
  or2_1 U11198 ( .ip1(n11169), .ip2(n11168), .op(n11170) );
  nand2_1 U11199 ( .ip1(n11171), .ip2(n11170), .op(n11257) );
  nand2_1 U11200 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[38]), .op(
        n11256) );
  inv_1 U11201 ( .ip(n11172), .op(n11270) );
  nand2_1 U11202 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[40]), .op(
        n11237) );
  nand2_1 U11203 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[42]), .op(
        n11192) );
  nor2_1 U11204 ( .ip1(n11173), .ip2(n11192), .op(n11188) );
  inv_1 U11205 ( .ip(n11174), .op(n11191) );
  or2_1 U11206 ( .ip1(m1Inputs[43]), .ip2(n11191), .op(n11176) );
  or2_1 U11207 ( .ip1(\STAGE_1/weightReg [9]), .ip2(n11191), .op(n11175) );
  nand2_1 U11208 ( .ip1(n11176), .ip2(n11175), .op(n11187) );
  nand2_1 U11209 ( .ip1(column[44]), .ip2(n13039), .op(n11189) );
  nor2_1 U11210 ( .ip1(n11187), .ip2(n11189), .op(n11177) );
  nor2_1 U11211 ( .ip1(n11188), .ip2(n11177), .op(n11236) );
  nand2_1 U11212 ( .ip1(n14816), .ip2(m1Inputs[39]), .op(n11235) );
  nand2_1 U11213 ( .ip1(m1Inputs[39]), .ip2(n15025), .op(n11179) );
  nand2_1 U11214 ( .ip1(m1Inputs[40]), .ip2(n13718), .op(n11178) );
  xor2_1 U11215 ( .ip1(n11179), .ip2(n11178), .op(n11204) );
  nor2_1 U11216 ( .ip1(n11181), .ip2(n11180), .op(n11182) );
  or2_1 U11217 ( .ip1(n11204), .ip2(n11182), .op(n11184) );
  nor2_1 U11218 ( .ip1(n14842), .ip2(n11555), .op(n11203) );
  or2_1 U11219 ( .ip1(n11203), .ip2(n11182), .op(n11183) );
  nand2_1 U11220 ( .ip1(n11184), .ip2(n11183), .op(n11250) );
  nand2_1 U11221 ( .ip1(m1Inputs[44]), .ip2(\STAGE_1/weightReg [7]), .op(
        n11206) );
  nand2_1 U11222 ( .ip1(m1Inputs[46]), .ip2(n12699), .op(n11205) );
  xnor2_1 U11223 ( .ip1(n11186), .ip2(n11185), .op(n11248) );
  nor2_1 U11224 ( .ip1(n11188), .ip2(n11187), .op(n11190) );
  xor2_1 U11225 ( .ip1(n11190), .ip2(n11189), .op(n11201) );
  nor2_1 U11226 ( .ip1(n12083), .ip2(n11544), .op(n11325) );
  nand2_1 U11227 ( .ip1(n11191), .ip2(n11325), .op(n11194) );
  inv_1 U11228 ( .ip(n11194), .op(n11197) );
  nand2_1 U11229 ( .ip1(m1Inputs[41]), .ip2(\STAGE_1/weightReg [10]), .op(
        n11193) );
  nand2_1 U11230 ( .ip1(n11193), .ip2(n11192), .op(n11195) );
  nand2_1 U11231 ( .ip1(n11195), .ip2(n11194), .op(n11214) );
  nand2_1 U11232 ( .ip1(column[43]), .ip2(n13039), .op(n11213) );
  nor2_1 U11233 ( .ip1(n11214), .ip2(n11213), .op(n11196) );
  nor2_1 U11234 ( .ip1(n11197), .ip2(n11196), .op(n11200) );
  nor2_1 U11235 ( .ip1(n14853), .ip2(n11477), .op(n11211) );
  nand2_1 U11236 ( .ip1(m1Inputs[45]), .ip2(\STAGE_1/weightReg [6]), .op(
        n11210) );
  nand2_1 U11237 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[43]), .op(
        n11209) );
  inv_1 U11238 ( .ip(n11198), .op(n11269) );
  fulladder U11239 ( .a(n11201), .b(n11200), .ci(n11199), .co(n11242), .s(
        n11202) );
  inv_1 U11240 ( .ip(n11202), .op(n11294) );
  xor2_1 U11241 ( .ip1(n11204), .ip2(n11203), .op(n11277) );
  fulladder U11242 ( .a(n11207), .b(n11206), .ci(n11205), .co(n11249), .s(
        n11208) );
  inv_1 U11243 ( .ip(n11208), .op(n11276) );
  fulladder U11244 ( .a(n11211), .b(n11210), .ci(n11209), .co(n11199), .s(
        n11212) );
  inv_1 U11245 ( .ip(n11212), .op(n11275) );
  xor2_1 U11246 ( .ip1(n11214), .ip2(n11213), .op(n11273) );
  nand2_1 U11247 ( .ip1(m1Inputs[46]), .ip2(n11974), .op(n11321) );
  nand2_1 U11248 ( .ip1(m1Inputs[43]), .ip2(\STAGE_1/weightReg [7]), .op(
        n11320) );
  inv_1 U11249 ( .ip(n11215), .op(n11272) );
  inv_1 U11250 ( .ip(m1Inputs[45]), .op(n11426) );
  nor2_1 U11251 ( .ip1(n11426), .ip2(n4624), .op(n11326) );
  nand2_1 U11252 ( .ip1(m1Inputs[35]), .ip2(n14976), .op(n11324) );
  inv_1 U11253 ( .ip(n11216), .op(n11784) );
  nand4_1 U11254 ( .ip1(\STAGE_1/weightReg [11]), .ip2(\STAGE_1/weightReg [10]), .ip3(m1Inputs[44]), .ip4(m1Inputs[43]), .op(n11776) );
  inv_1 U11255 ( .ip(n11776), .op(n11218) );
  or2_1 U11256 ( .ip1(n11217), .ip2(n11218), .op(n11221) );
  nand2_1 U11257 ( .ip1(n14629), .ip2(m1Inputs[44]), .op(n11219) );
  or2_1 U11258 ( .ip1(n11219), .ip2(n11218), .op(n11220) );
  nand2_1 U11259 ( .ip1(n11221), .ip2(n11220), .op(n11775) );
  nand2_1 U11260 ( .ip1(column[46]), .ip2(n13039), .op(n11222) );
  xor2_1 U11261 ( .ip1(n11775), .ip2(n11222), .op(n11824) );
  nand2_1 U11262 ( .ip1(n14816), .ip2(m1Inputs[40]), .op(n11791) );
  nand2_1 U11263 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[45]), .op(
        n11790) );
  fulladder U11264 ( .a(n11225), .b(n11224), .ci(n11223), .co(n11822), .s(
        n11233) );
  and3_1 U11265 ( .ip1(column[45]), .ip2(n13498), .ip3(n11226), .op(n11227) );
  nor2_1 U11266 ( .ip1(n11228), .ip2(n11227), .op(n11788) );
  fulladder U11267 ( .a(n11231), .b(n11230), .ci(n11229), .co(n11787), .s(
        n11234) );
  fulladder U11268 ( .a(n11234), .b(n11233), .ci(n11232), .co(n11811), .s(
        n11247) );
  fulladder U11269 ( .a(n11237), .b(n11236), .ci(n11235), .co(n11821), .s(
        n11244) );
  nor2_1 U11270 ( .ip1(n14902), .ip2(n11511), .op(n11803) );
  inv_1 U11271 ( .ip(m1Inputs[46]), .op(n11391) );
  nor2_1 U11272 ( .ip1(n6503), .ip2(n11391), .op(n11802) );
  nand2_1 U11273 ( .ip1(n14976), .ip2(m1Inputs[39]), .op(n11801) );
  inv_1 U11274 ( .ip(n11238), .op(n11820) );
  fulladder U11275 ( .a(n11241), .b(n11240), .ci(n11239), .co(n11819), .s(
        n11246) );
  fulladder U11276 ( .a(n11244), .b(n11243), .ci(n11242), .co(n11804), .s(
        n11198) );
  fulladder U11277 ( .a(n11247), .b(n11246), .ci(n11245), .co(n11782), .s(
        n11172) );
  fulladder U11278 ( .a(n11250), .b(n11249), .ci(n11248), .co(n11243), .s(
        n11251) );
  inv_1 U11279 ( .ip(n11251), .op(n11338) );
  fulladder U11280 ( .a(n11254), .b(n11253), .ci(n11252), .co(n11245), .s(
        n11255) );
  inv_1 U11281 ( .ip(n11255), .op(n11337) );
  fulladder U11282 ( .a(n11258), .b(n11257), .ci(n11256), .co(n11252), .s(
        n11259) );
  inv_1 U11283 ( .ip(n11259), .op(n11297) );
  nor3_1 U11284 ( .ip1(n11511), .ip2(n14836), .ip3(n11320), .op(n11264) );
  inv_1 U11285 ( .ip(m1Inputs[44]), .op(n11561) );
  inv_1 U11286 ( .ip(n11264), .op(n11263) );
  nand2_1 U11287 ( .ip1(m1Inputs[43]), .ip2(\STAGE_1/weightReg [6]), .op(
        n11261) );
  nand2_1 U11288 ( .ip1(m1Inputs[42]), .ip2(\STAGE_1/weightReg [7]), .op(
        n11260) );
  nand2_1 U11289 ( .ip1(n11261), .ip2(n11260), .op(n11262) );
  nand2_1 U11290 ( .ip1(n11263), .ip2(n11262), .op(n11313) );
  nor3_1 U11291 ( .ip1(n11561), .ip2(n12746), .ip3(n11313), .op(n11314) );
  nor2_1 U11292 ( .ip1(n11264), .ip2(n11314), .op(n11378) );
  nand2_1 U11293 ( .ip1(m1Inputs[45]), .ip2(n11974), .op(n11384) );
  nor2_1 U11294 ( .ip1(n11539), .ip2(n14853), .op(n11383) );
  nand2_1 U11295 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[41]), .op(
        n11382) );
  xor2_1 U11296 ( .ip1(n11266), .ip2(n11265), .op(n11376) );
  inv_1 U11297 ( .ip(n11267), .op(n11296) );
  nor2_1 U11298 ( .ip1(n14902), .ip2(n11283), .op(n11300) );
  nor2_1 U11299 ( .ip1(n14340), .ip2(n11555), .op(n11299) );
  and2_1 U11300 ( .ip1(column[41]), .ip2(n13498), .op(n11310) );
  nand2_1 U11301 ( .ip1(column[40]), .ip2(n13039), .op(n11363) );
  inv_1 U11302 ( .ip(n11363), .op(n11309) );
  nor2_1 U11303 ( .ip1(n12083), .ip2(n11461), .op(n11308) );
  fulladder U11304 ( .a(n11270), .b(n11269), .ci(n11268), .co(n11216), .s(
        n11333) );
  fulladder U11305 ( .a(n11273), .b(n11272), .ci(n11271), .co(n11292), .s(
        n11274) );
  inv_1 U11306 ( .ip(n11274), .op(n11346) );
  fulladder U11307 ( .a(n11277), .b(n11276), .ci(n11275), .co(n11293), .s(
        n11278) );
  inv_1 U11308 ( .ip(n11278), .op(n11345) );
  nor2_1 U11309 ( .ip1(n11280), .ip2(n11279), .op(n11282) );
  xor2_1 U11310 ( .ip1(n11282), .ip2(n11281), .op(n11381) );
  nor2_1 U11311 ( .ip1(n13594), .ip2(n11283), .op(n11327) );
  and3_1 U11312 ( .ip1(\STAGE_1/weightReg [11]), .ip2(m1Inputs[39]), .ip3(
        n11327), .op(n11288) );
  nor2_1 U11313 ( .ip1(n14824), .ip2(n11283), .op(n11284) );
  or2_1 U11314 ( .ip1(m1Inputs[39]), .ip2(n11284), .op(n11286) );
  or2_1 U11315 ( .ip1(n14876), .ip2(n11284), .op(n11285) );
  nand2_1 U11316 ( .ip1(n11286), .ip2(n11285), .op(n11287) );
  nor2_1 U11317 ( .ip1(n11288), .ip2(n11287), .op(n11319) );
  or2_1 U11318 ( .ip1(n11319), .ip2(n11288), .op(n11290) );
  nor2_1 U11319 ( .ip1(n14340), .ip2(n11477), .op(n11318) );
  or2_1 U11320 ( .ip1(n11318), .ip2(n11288), .op(n11289) );
  nand2_1 U11321 ( .ip1(n11290), .ip2(n11289), .op(n11380) );
  nand2_1 U11322 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[46]), .op(
        n11470) );
  nand2_1 U11323 ( .ip1(m1Inputs[35]), .ip2(n14816), .op(n11385) );
  inv_1 U11324 ( .ip(n11291), .op(n11342) );
  fulladder U11325 ( .a(n11294), .b(n11293), .ci(n11292), .co(n11268), .s(
        n11341) );
  fulladder U11326 ( .a(n11297), .b(n11296), .ci(n11295), .co(n11336), .s(
        n11405) );
  fulladder U11327 ( .a(n11300), .b(n11299), .ci(n11298), .co(n11295), .s(
        n11352) );
  nor2_1 U11328 ( .ip1(n11544), .ip2(n14289), .op(n11356) );
  and3_1 U11329 ( .ip1(m1Inputs[42]), .ip2(n4627), .ip3(n11356), .op(n11305)
         );
  nor2_1 U11330 ( .ip1(n11511), .ip2(n14836), .op(n11301) );
  or2_1 U11331 ( .ip1(\STAGE_1/weightReg [7]), .ip2(n11301), .op(n11303) );
  or2_1 U11332 ( .ip1(m1Inputs[41]), .ip2(n11301), .op(n11302) );
  nand2_1 U11333 ( .ip1(n11303), .ip2(n11302), .op(n11304) );
  nor2_1 U11334 ( .ip1(n11305), .ip2(n11304), .op(n11374) );
  or2_1 U11335 ( .ip1(n11374), .ip2(n11305), .op(n11307) );
  nor2_1 U11336 ( .ip1(n11472), .ip2(n12746), .op(n11373) );
  or2_1 U11337 ( .ip1(n11373), .ip2(n11305), .op(n11306) );
  nand2_1 U11338 ( .ip1(n11307), .ip2(n11306), .op(n11415) );
  nand2_1 U11339 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[45]), .op(
        n11509) );
  nand2_1 U11340 ( .ip1(m1Inputs[34]), .ip2(n14816), .op(n11420) );
  fulladder U11341 ( .a(n11310), .b(n11309), .ci(n11308), .co(n11298), .s(
        n11311) );
  inv_1 U11342 ( .ip(n11311), .op(n11413) );
  inv_1 U11343 ( .ip(n11312), .op(n11351) );
  or2_1 U11344 ( .ip1(n11313), .ip2(n11314), .op(n11317) );
  nand2_1 U11345 ( .ip1(m1Inputs[44]), .ip2(n12699), .op(n11315) );
  or2_1 U11346 ( .ip1(n11315), .ip2(n11314), .op(n11316) );
  nand2_1 U11347 ( .ip1(n11317), .ip2(n11316), .op(n11418) );
  xor2_1 U11348 ( .ip1(n11319), .ip2(n11318), .op(n11417) );
  nor2_1 U11349 ( .ip1(n11561), .ip2(n14783), .op(n11424) );
  nand2_1 U11350 ( .ip1(m1Inputs[33]), .ip2(n14976), .op(n11422) );
  fulladder U11351 ( .a(n11322), .b(n11321), .ci(n11320), .co(n11215), .s(
        n11323) );
  inv_1 U11352 ( .ip(n11323), .op(n11349) );
  fulladder U11353 ( .a(n11326), .b(n11325), .ci(n11324), .co(n11271), .s(
        n11348) );
  nor2_1 U11354 ( .ip1(n14188), .ip2(n11555), .op(n11355) );
  or2_1 U11355 ( .ip1(m1Inputs[37]), .ip2(n11327), .op(n11329) );
  or2_1 U11356 ( .ip1(n14847), .ip2(n11327), .op(n11328) );
  nand2_1 U11357 ( .ip1(n11329), .ip2(n11328), .op(n11368) );
  nor3_1 U11358 ( .ip1(n11368), .ip2(n11370), .ip3(n14373), .op(n11330) );
  nor2_1 U11359 ( .ip1(n13594), .ip2(n11555), .op(n11478) );
  and3_1 U11360 ( .ip1(n14847), .ip2(m1Inputs[38]), .ip3(n11478), .op(n11369)
         );
  or2_1 U11361 ( .ip1(n11330), .ip2(n11369), .op(n11354) );
  nor2_1 U11362 ( .ip1(n12083), .ip2(n11534), .op(n11365) );
  nor2_1 U11363 ( .ip1(n13854), .ip2(n11391), .op(n11364) );
  inv_1 U11364 ( .ip(n11331), .op(n11815) );
  fulladder U11365 ( .a(n11334), .b(n11333), .ci(n11332), .co(n11331), .s(
        n11335) );
  inv_1 U11366 ( .ip(n11335), .op(n11741) );
  fulladder U11367 ( .a(n11338), .b(n11337), .ci(n11336), .co(n11334), .s(
        n11339) );
  inv_1 U11368 ( .ip(n11339), .op(n11402) );
  fulladder U11369 ( .a(n11342), .b(n11341), .ci(n11340), .co(n11332), .s(
        n11343) );
  inv_1 U11370 ( .ip(n11343), .op(n11401) );
  fulladder U11371 ( .a(n11346), .b(n11345), .ci(n11344), .co(n11291), .s(
        n11409) );
  fulladder U11372 ( .a(n11349), .b(n11348), .ci(n11347), .co(n11403), .s(
        n11490) );
  fulladder U11373 ( .a(n11352), .b(n11351), .ci(n11350), .co(n11404), .s(
        n11489) );
  fulladder U11374 ( .a(n11355), .b(n11354), .ci(n11353), .co(n11347), .s(
        n11497) );
  nand2_1 U11375 ( .ip1(m1Inputs[41]), .ip2(n11974), .op(n11546) );
  nor3_1 U11376 ( .ip1(n11472), .ip2(n14289), .ip3(n11546), .op(n11360) );
  or2_1 U11377 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n11356), .op(n11358) );
  or2_1 U11378 ( .ip1(m1Inputs[43]), .ip2(n11356), .op(n11357) );
  nand2_1 U11379 ( .ip1(n11358), .ip2(n11357), .op(n11359) );
  nor2_1 U11380 ( .ip1(n11360), .ip2(n11359), .op(n11445) );
  or2_1 U11381 ( .ip1(n11445), .ip2(n11360), .op(n11362) );
  nor2_1 U11382 ( .ip1(n11549), .ip2(n14842), .op(n11444) );
  or2_1 U11383 ( .ip1(n11444), .ip2(n11360), .op(n11361) );
  nand2_1 U11384 ( .ip1(n11362), .ip2(n11361), .op(n11451) );
  nor2_1 U11385 ( .ip1(n13646), .ip2(n11858), .op(n11439) );
  nand2_1 U11386 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[38]), .op(
        n11438) );
  fulladder U11387 ( .a(n11365), .b(n11364), .ci(n11363), .co(n11353), .s(
        n11366) );
  inv_1 U11388 ( .ip(n11366), .op(n11449) );
  inv_1 U11389 ( .ip(n11367), .op(n11496) );
  nor2_1 U11390 ( .ip1(n11369), .ip2(n11368), .op(n11372) );
  nor2_1 U11391 ( .ip1(n11370), .ip2(n14340), .op(n11371) );
  xor2_1 U11392 ( .ip1(n11372), .ip2(n11371), .op(n11448) );
  xor2_1 U11393 ( .ip1(n11374), .ip2(n11373), .op(n11447) );
  nor2_1 U11394 ( .ip1(n11511), .ip2(n12746), .op(n11443) );
  nand2_1 U11395 ( .ip1(m1Inputs[32]), .ip2(n14976), .op(n11442) );
  inv_1 U11396 ( .ip(n11375), .op(n11408) );
  fulladder U11397 ( .a(n11378), .b(n11377), .ci(n11376), .co(n11267), .s(
        n11412) );
  fulladder U11398 ( .a(n11381), .b(n11380), .ci(n11379), .co(n11344), .s(
        n11411) );
  fulladder U11399 ( .a(n11384), .b(n11383), .ci(n11382), .co(n11377), .s(
        n11437) );
  fulladder U11400 ( .a(n11470), .b(n11386), .ci(n11385), .co(n11379), .s(
        n11436) );
  nor2_1 U11401 ( .ip1(n11534), .ip2(n12156), .op(n11462) );
  and2_1 U11402 ( .ip1(n11423), .ip2(n11462), .op(n11467) );
  nor2_1 U11403 ( .ip1(n11461), .ip2(n12156), .op(n11387) );
  or2_1 U11404 ( .ip1(m1Inputs[39]), .ip2(n11387), .op(n11389) );
  or2_1 U11405 ( .ip1(n14838), .ip2(n11387), .op(n11388) );
  nand2_1 U11406 ( .ip1(n11389), .ip2(n11388), .op(n11466) );
  nand2_1 U11407 ( .ip1(m1Inputs[34]), .ip2(n15028), .op(n11468) );
  nor2_1 U11408 ( .ip1(n11466), .ip2(n11468), .op(n11390) );
  nor2_1 U11409 ( .ip1(n11467), .ip2(n11390), .op(n11456) );
  nand2_1 U11410 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[45]), .op(
        n11392) );
  nand2_1 U11411 ( .ip1(n12809), .ip2(m1Inputs[45]), .op(n11428) );
  nor3_1 U11412 ( .ip1(n13709), .ip2(n11391), .ip3(n11428), .op(n11396) );
  or2_1 U11413 ( .ip1(n11392), .ip2(n11396), .op(n11395) );
  nand2_1 U11414 ( .ip1(n12809), .ip2(m1Inputs[46]), .op(n11393) );
  or2_1 U11415 ( .ip1(n11393), .ip2(n11396), .op(n11394) );
  nand2_1 U11416 ( .ip1(n11395), .ip2(n11394), .op(n11484) );
  or2_1 U11417 ( .ip1(n11484), .ip2(n11396), .op(n11399) );
  nand2_1 U11418 ( .ip1(column[39]), .ip2(n13039), .op(n11483) );
  inv_1 U11419 ( .ip(n11483), .op(n11397) );
  or2_1 U11420 ( .ip1(n11397), .ip2(n11396), .op(n11398) );
  nand2_1 U11421 ( .ip1(n11399), .ip2(n11398), .op(n11455) );
  nand2_1 U11422 ( .ip1(n15025), .ip2(m1Inputs[36]), .op(n11454) );
  fulladder U11423 ( .a(n11402), .b(n11401), .ci(n11400), .co(n11740), .s(
        n11745) );
  fulladder U11424 ( .a(n11405), .b(n11404), .ci(n11403), .co(n11340), .s(
        n11406) );
  inv_1 U11425 ( .ip(n11406), .op(n11487) );
  fulladder U11426 ( .a(n11409), .b(n11408), .ci(n11407), .co(n11400), .s(
        n11486) );
  fulladder U11427 ( .a(n11412), .b(n11411), .ci(n11410), .co(n11407), .s(
        n11494) );
  fulladder U11428 ( .a(n11415), .b(n11414), .ci(n11413), .co(n11312), .s(
        n11501) );
  fulladder U11429 ( .a(n11418), .b(n11417), .ci(n11416), .co(n11350), .s(
        n11419) );
  inv_1 U11430 ( .ip(n11419), .op(n11500) );
  fulladder U11431 ( .a(n11421), .b(n11509), .ci(n11420), .co(n11414), .s(
        n11504) );
  fulladder U11432 ( .a(n11424), .b(n11423), .ci(n11422), .co(n11416), .s(
        n11425) );
  inv_1 U11433 ( .ip(n11425), .op(n11503) );
  nand2_1 U11434 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[44]), .op(
        n11427) );
  nand2_1 U11435 ( .ip1(n12809), .ip2(m1Inputs[44]), .op(n11563) );
  nor3_1 U11436 ( .ip1(n13709), .ip2(n11426), .ip3(n11563), .op(n11431) );
  or2_1 U11437 ( .ip1(n11427), .ip2(n11431), .op(n11430) );
  or2_1 U11438 ( .ip1(n11428), .ip2(n11431), .op(n11429) );
  nand2_1 U11439 ( .ip1(n11430), .ip2(n11429), .op(n11554) );
  or2_1 U11440 ( .ip1(n11554), .ip2(n11431), .op(n11434) );
  nand2_1 U11441 ( .ip1(column[38]), .ip2(n13039), .op(n11553) );
  inv_1 U11442 ( .ip(n11553), .op(n11432) );
  or2_1 U11443 ( .ip1(n11432), .ip2(n11431), .op(n11433) );
  nand2_1 U11444 ( .ip1(n11434), .ip2(n11433), .op(n11532) );
  nand2_1 U11445 ( .ip1(m1Inputs[35]), .ip2(n15025), .op(n11531) );
  nand2_1 U11446 ( .ip1(n13718), .ip2(m1Inputs[36]), .op(n11530) );
  fulladder U11447 ( .a(n11437), .b(n11436), .ci(n11435), .co(n11410), .s(
        n11575) );
  fulladder U11448 ( .a(n11440), .b(n11439), .ci(n11438), .co(n11450), .s(
        n11441) );
  inv_1 U11449 ( .ip(n11441), .op(n11588) );
  fulladder U11450 ( .a(n11443), .b(n11478), .ci(n11442), .co(n11446), .s(
        n11587) );
  xor2_1 U11451 ( .ip1(n11445), .ip2(n11444), .op(n11586) );
  fulladder U11452 ( .a(n11448), .b(n11447), .ci(n11446), .co(n11495), .s(
        n11583) );
  fulladder U11453 ( .a(n11451), .b(n11450), .ci(n11449), .co(n11367), .s(
        n11452) );
  inv_1 U11454 ( .ip(n11452), .op(n11582) );
  inv_1 U11455 ( .ip(n11453), .op(n11574) );
  fulladder U11456 ( .a(n11456), .b(n11455), .ci(n11454), .co(n11435), .s(
        n11581) );
  nor3_1 U11457 ( .ip1(n11511), .ip2(n13835), .ip3(n11546), .op(n11604) );
  nor2_1 U11458 ( .ip1(n11544), .ip2(n12746), .op(n11457) );
  or2_1 U11459 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n11457), .op(n11459) );
  or2_1 U11460 ( .ip1(m1Inputs[42]), .ip2(n11457), .op(n11458) );
  nand2_1 U11461 ( .ip1(n11459), .ip2(n11458), .op(n11603) );
  nand2_1 U11462 ( .ip1(n14975), .ip2(m1Inputs[38]), .op(n11605) );
  nor2_1 U11463 ( .ip1(n11603), .ip2(n11605), .op(n11460) );
  nor2_1 U11464 ( .ip1(n11604), .ip2(n11460), .op(n11526) );
  nor3_1 U11465 ( .ip1(n11461), .ip2(n14384), .ip3(n11536), .op(n11506) );
  or2_1 U11466 ( .ip1(n13749), .ip2(n11462), .op(n11464) );
  or2_1 U11467 ( .ip1(m1Inputs[40]), .ip2(n11462), .op(n11463) );
  nand2_1 U11468 ( .ip1(n11464), .ip2(n11463), .op(n11505) );
  nand2_1 U11469 ( .ip1(m1Inputs[33]), .ip2(\STAGE_1/weightReg [13]), .op(
        n11507) );
  nor2_1 U11470 ( .ip1(n11505), .ip2(n11507), .op(n11465) );
  nor2_1 U11471 ( .ip1(n11506), .ip2(n11465), .op(n11525) );
  nor2_1 U11472 ( .ip1(n11467), .ip2(n11466), .op(n11469) );
  xor2_1 U11473 ( .ip1(n11469), .ip2(n11468), .op(n11524) );
  nor2_1 U11474 ( .ip1(n11471), .ip2(n11470), .op(n11608) );
  nor2_1 U11475 ( .ip1(n13801), .ip2(n11472), .op(n11473) );
  or2_1 U11476 ( .ip1(m1Inputs[46]), .ip2(n11473), .op(n11475) );
  or2_1 U11477 ( .ip1(n13803), .ip2(n11473), .op(n11474) );
  nand2_1 U11478 ( .ip1(n11475), .ip2(n11474), .op(n11607) );
  nand2_1 U11479 ( .ip1(m1Inputs[32]), .ip2(n14816), .op(n11609) );
  nor2_1 U11480 ( .ip1(n11607), .ip2(n11609), .op(n11476) );
  nor2_1 U11481 ( .ip1(n11608), .ip2(n11476), .op(n11529) );
  nor2_1 U11482 ( .ip1(n12083), .ip2(n11477), .op(n11556) );
  and2_1 U11483 ( .ip1(n11556), .ip2(n11478), .op(n11521) );
  nor2_1 U11484 ( .ip1(n12083), .ip2(n11555), .op(n11479) );
  or2_1 U11485 ( .ip1(m1Inputs[36]), .ip2(n11479), .op(n11481) );
  or2_1 U11486 ( .ip1(n14876), .ip2(n11479), .op(n11480) );
  nand2_1 U11487 ( .ip1(n11481), .ip2(n11480), .op(n11520) );
  nand2_1 U11488 ( .ip1(m1Inputs[34]), .ip2(n15025), .op(n11522) );
  nor2_1 U11489 ( .ip1(n11520), .ip2(n11522), .op(n11482) );
  nor2_1 U11490 ( .ip1(n11521), .ip2(n11482), .op(n11528) );
  xor2_1 U11491 ( .ip1(n11484), .ip2(n11483), .op(n11527) );
  fulladder U11492 ( .a(n11487), .b(n11486), .ci(n11485), .co(n11744), .s(
        n11749) );
  fulladder U11493 ( .a(n11490), .b(n11489), .ci(n11488), .co(n11375), .s(
        n11491) );
  inv_1 U11494 ( .ip(n11491), .op(n11572) );
  fulladder U11495 ( .a(n11494), .b(n11493), .ci(n11492), .co(n11485), .s(
        n11571) );
  fulladder U11496 ( .a(n11497), .b(n11496), .ci(n11495), .co(n11488), .s(
        n11498) );
  inv_1 U11497 ( .ip(n11498), .op(n11578) );
  fulladder U11498 ( .a(n11501), .b(n11500), .ci(n11499), .co(n11493), .s(
        n11577) );
  fulladder U11499 ( .a(n11504), .b(n11503), .ci(n11502), .co(n11499), .s(
        n11639) );
  nor2_1 U11500 ( .ip1(n11506), .ip2(n11505), .op(n11508) );
  xor2_1 U11501 ( .ip1(n11508), .ip2(n11507), .op(n11651) );
  nor2_1 U11502 ( .ip1(n11510), .ip2(n11509), .op(n11517) );
  nor2_1 U11503 ( .ip1(n13801), .ip2(n11511), .op(n11512) );
  or2_1 U11504 ( .ip1(m1Inputs[45]), .ip2(n11512), .op(n11514) );
  or2_1 U11505 ( .ip1(n13803), .ip2(n11512), .op(n11513) );
  nand2_1 U11506 ( .ip1(n11514), .ip2(n11513), .op(n11515) );
  nor2_1 U11507 ( .ip1(n11517), .ip2(n11515), .op(n11658) );
  or2_1 U11508 ( .ip1(n11658), .ip2(n11517), .op(n11519) );
  nor2_1 U11509 ( .ip1(n11516), .ip2(n14340), .op(n11657) );
  or2_1 U11510 ( .ip1(n11657), .ip2(n11517), .op(n11518) );
  nand2_1 U11511 ( .ip1(n11519), .ip2(n11518), .op(n11650) );
  nor2_1 U11512 ( .ip1(n11521), .ip2(n11520), .op(n11523) );
  xor2_1 U11513 ( .ip1(n11523), .ip2(n11522), .op(n11649) );
  fulladder U11514 ( .a(n11526), .b(n11525), .ci(n11524), .co(n11580), .s(
        n11646) );
  fulladder U11515 ( .a(n11529), .b(n11528), .ci(n11527), .co(n11579), .s(
        n11645) );
  fulladder U11516 ( .a(n11532), .b(n11531), .ci(n11530), .co(n11502), .s(
        n11643) );
  nand2_1 U11517 ( .ip1(m1Inputs[38]), .ip2(n4627), .op(n11535) );
  nor3_1 U11518 ( .ip1(n11534), .ip2(n14384), .ip3(n11533), .op(n11540) );
  or2_1 U11519 ( .ip1(n11535), .ip2(n11540), .op(n11538) );
  or2_1 U11520 ( .ip1(n11536), .ip2(n11540), .op(n11537) );
  nand2_1 U11521 ( .ip1(n11538), .ip2(n11537), .op(n11662) );
  or2_1 U11522 ( .ip1(n11662), .ip2(n11540), .op(n11542) );
  nor2_1 U11523 ( .ip1(n11539), .ip2(n14824), .op(n11661) );
  or2_1 U11524 ( .ip1(n11661), .ip2(n11540), .op(n11541) );
  nand2_1 U11525 ( .ip1(n11542), .ip2(n11541), .op(n11616) );
  nand2_1 U11526 ( .ip1(m1Inputs[40]), .ip2(n12699), .op(n11545) );
  nor3_1 U11527 ( .ip1(n11544), .ip2(n13835), .ip3(n11543), .op(n11550) );
  or2_1 U11528 ( .ip1(n11545), .ip2(n11550), .op(n11548) );
  or2_1 U11529 ( .ip1(n11546), .ip2(n11550), .op(n11547) );
  nand2_1 U11530 ( .ip1(n11548), .ip2(n11547), .op(n11660) );
  or2_1 U11531 ( .ip1(n11660), .ip2(n11550), .op(n11552) );
  nor2_1 U11532 ( .ip1(n11549), .ip2(n14188), .op(n11659) );
  or2_1 U11533 ( .ip1(n11659), .ip2(n11550), .op(n11551) );
  nand2_1 U11534 ( .ip1(n11552), .ip2(n11551), .op(n11615) );
  xor2_1 U11535 ( .ip1(n11554), .ip2(n11553), .op(n11614) );
  nor3_1 U11536 ( .ip1(n12083), .ip2(n11555), .ip3(n11690), .op(n11627) );
  or2_1 U11537 ( .ip1(m1Inputs[37]), .ip2(n11556), .op(n11558) );
  or2_1 U11538 ( .ip1(n14838), .ip2(n11556), .op(n11557) );
  nand2_1 U11539 ( .ip1(n11558), .ip2(n11557), .op(n11626) );
  nand2_1 U11540 ( .ip1(m1Inputs[35]), .ip2(n14876), .op(n11628) );
  nor2_1 U11541 ( .ip1(n11626), .ip2(n11628), .op(n11559) );
  nor2_1 U11542 ( .ip1(n11627), .ip2(n11559), .op(n11613) );
  nand2_1 U11543 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[43]), .op(
        n11562) );
  nor3_1 U11544 ( .ip1(n13709), .ip2(n11561), .ip3(n11560), .op(n11566) );
  or2_1 U11545 ( .ip1(n11562), .ip2(n11566), .op(n11565) );
  or2_1 U11546 ( .ip1(n11563), .ip2(n11566), .op(n11564) );
  nand2_1 U11547 ( .ip1(n11565), .ip2(n11564), .op(n11602) );
  or2_1 U11548 ( .ip1(n11602), .ip2(n11566), .op(n11569) );
  nand2_1 U11549 ( .ip1(column[37]), .ip2(n13039), .op(n11601) );
  inv_1 U11550 ( .ip(n11601), .op(n11567) );
  or2_1 U11551 ( .ip1(n11567), .ip2(n11566), .op(n11568) );
  nand2_1 U11552 ( .ip1(n11569), .ip2(n11568), .op(n11612) );
  nand2_1 U11553 ( .ip1(m1Inputs[35]), .ip2(n14847), .op(n11611) );
  fulladder U11554 ( .a(n11572), .b(n11571), .ci(n11570), .co(n11748), .s(
        n11753) );
  fulladder U11555 ( .a(n11575), .b(n11574), .ci(n11573), .co(n11492), .s(
        n11632) );
  fulladder U11556 ( .a(n11578), .b(n11577), .ci(n11576), .co(n11570), .s(
        n11631) );
  fulladder U11557 ( .a(n11581), .b(n11580), .ci(n11579), .co(n11573), .s(
        n11635) );
  fulladder U11558 ( .a(n11584), .b(n11583), .ci(n11582), .co(n11453), .s(
        n11585) );
  inv_1 U11559 ( .ip(n11585), .op(n11634) );
  fulladder U11560 ( .a(n11588), .b(n11587), .ci(n11586), .co(n11584), .s(
        n11589) );
  inv_1 U11561 ( .ip(n11589), .op(n11670) );
  or2_1 U11562 ( .ip1(n11590), .ip2(n11592), .op(n11595) );
  inv_1 U11563 ( .ip(n11591), .op(n11593) );
  or2_1 U11564 ( .ip1(n11593), .ip2(n11592), .op(n11594) );
  nand2_1 U11565 ( .ip1(n11595), .ip2(n11594), .op(n11687) );
  or2_1 U11566 ( .ip1(n11596), .ip2(n11597), .op(n11600) );
  or2_1 U11567 ( .ip1(n11598), .ip2(n11597), .op(n11599) );
  nand2_1 U11568 ( .ip1(n11600), .ip2(n11599), .op(n11686) );
  xor2_1 U11569 ( .ip1(n11602), .ip2(n11601), .op(n11685) );
  nor2_1 U11570 ( .ip1(n11604), .ip2(n11603), .op(n11606) );
  xor2_1 U11571 ( .ip1(n11606), .ip2(n11605), .op(n11654) );
  nor2_1 U11572 ( .ip1(n11608), .ip2(n11607), .op(n11610) );
  xor2_1 U11573 ( .ip1(n11610), .ip2(n11609), .op(n11653) );
  fulladder U11574 ( .a(n11613), .b(n11612), .ci(n11611), .co(n11641), .s(
        n11677) );
  fulladder U11575 ( .a(n11616), .b(n11615), .ci(n11614), .co(n11642), .s(
        n11676) );
  or2_1 U11576 ( .ip1(n11617), .ip2(n11618), .op(n11621) );
  or2_1 U11577 ( .ip1(n11619), .ip2(n11618), .op(n11620) );
  nand2_1 U11578 ( .ip1(n11621), .ip2(n11620), .op(n11680) );
  nor2_1 U11579 ( .ip1(n11623), .ip2(n11622), .op(n11624) );
  nor2_1 U11580 ( .ip1(n11625), .ip2(n11624), .op(n11679) );
  nor2_1 U11581 ( .ip1(n11627), .ip2(n11626), .op(n11629) );
  xor2_1 U11582 ( .ip1(n11629), .ip2(n11628), .op(n11678) );
  fulladder U11583 ( .a(n11632), .b(n11631), .ci(n11630), .co(n11752), .s(
        n11757) );
  fulladder U11584 ( .a(n11635), .b(n11634), .ci(n11633), .co(n11630), .s(
        n11636) );
  inv_1 U11585 ( .ip(n11636), .op(n11666) );
  fulladder U11586 ( .a(n11639), .b(n11638), .ci(n11637), .co(n11576), .s(
        n11640) );
  inv_1 U11587 ( .ip(n11640), .op(n11665) );
  fulladder U11588 ( .a(n11643), .b(n11642), .ci(n11641), .co(n11637), .s(
        n11644) );
  inv_1 U11589 ( .ip(n11644), .op(n11673) );
  fulladder U11590 ( .a(n11647), .b(n11646), .ci(n11645), .co(n11638), .s(
        n11648) );
  inv_1 U11591 ( .ip(n11648), .op(n11672) );
  fulladder U11592 ( .a(n11651), .b(n11650), .ci(n11649), .co(n11647), .s(
        n11652) );
  inv_1 U11593 ( .ip(n11652), .op(n11702) );
  fulladder U11594 ( .a(n11655), .b(n11654), .ci(n11653), .co(n11669), .s(
        n11656) );
  inv_1 U11595 ( .ip(n11656), .op(n11701) );
  xor2_1 U11596 ( .ip1(n11658), .ip2(n11657), .op(n11683) );
  xor2_1 U11597 ( .ip1(n11660), .ip2(n11659), .op(n11682) );
  xor2_1 U11598 ( .ip1(n11662), .ip2(n11661), .op(n11681) );
  inv_1 U11599 ( .ip(n11663), .op(n11756) );
  fulladder U11600 ( .a(n11666), .b(n11665), .ci(n11664), .co(n11663), .s(
        n11667) );
  inv_1 U11601 ( .ip(n11667), .op(n11761) );
  fulladder U11602 ( .a(n11670), .b(n11669), .ci(n11668), .co(n11633), .s(
        n11699) );
  fulladder U11603 ( .a(n11673), .b(n11672), .ci(n11671), .co(n11664), .s(
        n11674) );
  inv_1 U11604 ( .ip(n11674), .op(n11698) );
  fulladder U11605 ( .a(n11677), .b(n11676), .ci(n11675), .co(n11668), .s(
        n11706) );
  fulladder U11606 ( .a(n11680), .b(n11679), .ci(n11678), .co(n11675), .s(
        n11721) );
  fulladder U11607 ( .a(n11683), .b(n11682), .ci(n11681), .co(n11700), .s(
        n11684) );
  inv_1 U11608 ( .ip(n11684), .op(n11720) );
  fulladder U11609 ( .a(n11687), .b(n11686), .ci(n11685), .co(n11655), .s(
        n11719) );
  fulladder U11610 ( .a(n11690), .b(n11689), .ci(n11688), .co(n11709), .s(
        n11711) );
  fulladder U11611 ( .a(n11693), .b(n11692), .ci(n11691), .co(n11708), .s(
        n11715) );
  fulladder U11612 ( .a(n11696), .b(n11695), .ci(n11694), .co(n11707), .s(
        n11727) );
  fulladder U11613 ( .a(n11699), .b(n11698), .ci(n11697), .co(n11760), .s(
        n11765) );
  fulladder U11614 ( .a(n11702), .b(n11701), .ci(n11700), .co(n11671), .s(
        n11703) );
  inv_1 U11615 ( .ip(n11703), .op(n11718) );
  fulladder U11616 ( .a(n11706), .b(n11705), .ci(n11704), .co(n11697), .s(
        n11717) );
  fulladder U11617 ( .a(n11709), .b(n11708), .ci(n11707), .co(n11704), .s(
        n11724) );
  fulladder U11618 ( .a(n11712), .b(n11711), .ci(n11710), .co(n11723), .s(
        n11726) );
  fulladder U11619 ( .a(n11715), .b(n11714), .ci(n11713), .co(n11722), .s(
        n11737) );
  fulladder U11620 ( .a(n11718), .b(n11717), .ci(n11716), .co(n11764), .s(
        n11769) );
  fulladder U11621 ( .a(n11721), .b(n11720), .ci(n11719), .co(n11705), .s(
        n11730) );
  fulladder U11622 ( .a(n11724), .b(n11723), .ci(n11722), .co(n11716), .s(
        n11729) );
  fulladder U11623 ( .a(n11727), .b(n11726), .ci(n11725), .co(n11728), .s(
        n11736) );
  fulladder U11624 ( .a(n11730), .b(n11729), .ci(n11728), .co(n11768), .s(
        n11773) );
  fulladder U11625 ( .a(n11733), .b(n11732), .ci(n11731), .co(n11734), .s(
        \STAGE_1/M3/sum [4]) );
  inv_1 U11626 ( .ip(n11734), .op(n11772) );
  fulladder U11627 ( .a(n11737), .b(n11736), .ci(n11735), .co(n11771), .s(
        n11140) );
  inv_1 U11628 ( .ip(n11738), .op(\STAGE_1/M3/sum [14]) );
  fulladder U11629 ( .a(n11741), .b(n11740), .ci(n11739), .co(n11814), .s(
        n11742) );
  inv_1 U11630 ( .ip(n11742), .op(\STAGE_1/M3/sum [13]) );
  fulladder U11631 ( .a(n11745), .b(n11744), .ci(n11743), .co(n11739), .s(
        n11746) );
  inv_1 U11632 ( .ip(n11746), .op(\STAGE_1/M3/sum [12]) );
  fulladder U11633 ( .a(n11749), .b(n11748), .ci(n11747), .co(n11743), .s(
        n11750) );
  inv_1 U11634 ( .ip(n11750), .op(\STAGE_1/M3/sum [11]) );
  fulladder U11635 ( .a(n11753), .b(n11752), .ci(n11751), .co(n11747), .s(
        n11754) );
  inv_1 U11636 ( .ip(n11754), .op(\STAGE_1/M3/sum [10]) );
  fulladder U11637 ( .a(n11757), .b(n11756), .ci(n11755), .co(n11751), .s(
        n11758) );
  inv_1 U11638 ( .ip(n11758), .op(\STAGE_1/M3/sum [9]) );
  fulladder U11639 ( .a(n11761), .b(n11760), .ci(n11759), .co(n11755), .s(
        n11762) );
  inv_1 U11640 ( .ip(n11762), .op(\STAGE_1/M3/sum [8]) );
  fulladder U11641 ( .a(n11765), .b(n11764), .ci(n11763), .co(n11759), .s(
        n11766) );
  inv_1 U11642 ( .ip(n11766), .op(\STAGE_1/M3/sum [7]) );
  fulladder U11643 ( .a(n11769), .b(n11768), .ci(n11767), .co(n11763), .s(
        n11770) );
  inv_1 U11644 ( .ip(n11770), .op(\STAGE_1/M3/sum [6]) );
  fulladder U11645 ( .a(n11773), .b(n11772), .ci(n11771), .co(n11767), .s(
        n11774) );
  inv_1 U11646 ( .ip(n11774), .op(\STAGE_1/M3/sum [5]) );
  nand2_1 U11647 ( .ip1(column[47]), .ip2(n13039), .op(n11779) );
  nand3_1 U11648 ( .ip1(column[46]), .ip2(n15042), .ip3(n11775), .op(n11777)
         );
  nand2_1 U11649 ( .ip1(n11777), .ip2(n11776), .op(n11778) );
  xor2_1 U11650 ( .ip1(n11779), .ip2(n11778), .op(n11840) );
  nand2_1 U11651 ( .ip1(m1Inputs[42]), .ip2(n15028), .op(n11781) );
  nand2_1 U11652 ( .ip1(m1Inputs[40]), .ip2(n14976), .op(n11780) );
  xor2_1 U11653 ( .ip1(n11781), .ip2(n11780), .op(n11786) );
  fulladder U11654 ( .a(n11784), .b(n11783), .ci(n11782), .co(n11785), .s(
        n11816) );
  xor2_1 U11655 ( .ip1(n11786), .ip2(n11785), .op(n11796) );
  fulladder U11656 ( .a(n11789), .b(n11788), .ci(n11787), .co(n11794), .s(
        n11812) );
  fulladder U11657 ( .a(n11792), .b(n11791), .ci(n11790), .co(n11793), .s(
        n11823) );
  xor2_1 U11658 ( .ip1(n11794), .ip2(n11793), .op(n11795) );
  xor2_1 U11659 ( .ip1(n11796), .ip2(n11795), .op(n11798) );
  nand2_1 U11660 ( .ip1(m1Inputs[46]), .ip2(n14994), .op(n11797) );
  xor2_1 U11661 ( .ip1(n11798), .ip2(n11797), .op(n11838) );
  nand2_1 U11662 ( .ip1(m1Inputs[43]), .ip2(n15025), .op(n11800) );
  nand2_1 U11663 ( .ip1(m1Inputs[45]), .ip2(n14629), .op(n11799) );
  xor2_1 U11664 ( .ip1(n11800), .ip2(n11799), .op(n11836) );
  fulladder U11665 ( .a(n11803), .b(n11802), .ci(n11801), .co(n11808), .s(
        n11238) );
  fulladder U11666 ( .a(n11806), .b(n11805), .ci(n11804), .co(n11807), .s(
        n11783) );
  xor2_1 U11667 ( .ip1(n11808), .ip2(n11807), .op(n11809) );
  xor2_1 U11668 ( .ip1(n11810), .ip2(n11809), .op(n11834) );
  fulladder U11669 ( .a(n11813), .b(n11812), .ci(n11811), .co(n11818), .s(
        n11806) );
  fulladder U11670 ( .a(n11816), .b(n11815), .ci(n11814), .co(n11817), .s(
        n11738) );
  xor2_1 U11671 ( .ip1(n11818), .ip2(n11817), .op(n11828) );
  fulladder U11672 ( .a(n11821), .b(n11820), .ci(n11819), .co(n11826), .s(
        n11805) );
  fulladder U11673 ( .a(n11824), .b(n11823), .ci(n11822), .co(n11825), .s(
        n11813) );
  xor2_1 U11674 ( .ip1(n11826), .ip2(n11825), .op(n11827) );
  xor2_1 U11675 ( .ip1(n11828), .ip2(n11827), .op(n11832) );
  nand2_1 U11676 ( .ip1(m1Inputs[41]), .ip2(n14816), .op(n11829) );
  xnor2_1 U11677 ( .ip1(n11830), .ip2(n11829), .op(n11831) );
  xor2_1 U11678 ( .ip1(n11832), .ip2(n11831), .op(n11833) );
  xor2_1 U11679 ( .ip1(n11834), .ip2(n11833), .op(n11835) );
  xor2_1 U11680 ( .ip1(n11836), .ip2(n11835), .op(n11837) );
  xor2_1 U11681 ( .ip1(n11838), .ip2(n11837), .op(n11839) );
  xor2_1 U11682 ( .ip1(n11840), .ip2(n11839), .op(\STAGE_1/M3/sum [15]) );
  or2_1 U11683 ( .ip1(n11841), .ip2(n11842), .op(n11845) );
  or2_1 U11684 ( .ip1(n11843), .ip2(n11842), .op(n11844) );
  nand2_1 U11685 ( .ip1(n11845), .ip2(n11844), .op(n12365) );
  nor2_1 U11686 ( .ip1(n11847), .ip2(n11846), .op(n11848) );
  nor2_1 U11687 ( .ip1(n11849), .ip2(n11848), .op(n12364) );
  nor3_1 U11688 ( .ip1(n12083), .ip2(n12255), .ip3(n11885), .op(n12319) );
  inv_1 U11689 ( .ip(\STAGE_1/weightReg [9]), .op(n13766) );
  nor2_1 U11690 ( .ip1(n13766), .ip2(n12066), .op(n12254) );
  or2_1 U11691 ( .ip1(m1Inputs[53]), .ip2(n12254), .op(n11851) );
  or2_1 U11692 ( .ip1(n14838), .ip2(n12254), .op(n11850) );
  nand2_1 U11693 ( .ip1(n11851), .ip2(n11850), .op(n12317) );
  nor2_1 U11694 ( .ip1(n12319), .ip2(n12317), .op(n11852) );
  nand2_1 U11695 ( .ip1(m1Inputs[51]), .ip2(n14629), .op(n12316) );
  xor2_1 U11696 ( .ip1(n11852), .ip2(n12316), .op(n12363) );
  nand2_1 U11697 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[61]), .op(
        n12192) );
  nor2_1 U11698 ( .ip1(n11853), .ip2(n12192), .op(n12287) );
  nor2_1 U11699 ( .ip1(n13082), .ip2(n12230), .op(n11854) );
  or2_1 U11700 ( .ip1(m1Inputs[61]), .ip2(n11854), .op(n11856) );
  or2_1 U11701 ( .ip1(n13803), .ip2(n11854), .op(n11855) );
  nand2_1 U11702 ( .ip1(n11856), .ip2(n11855), .op(n11857) );
  nor2_1 U11703 ( .ip1(n12287), .ip2(n11857), .op(n12286) );
  nor2_1 U11704 ( .ip1(n11858), .ip2(n14340), .op(n12288) );
  xor2_1 U11705 ( .ip1(n12286), .ip2(n12288), .op(n12395) );
  nand2_1 U11706 ( .ip1(m1Inputs[56]), .ip2(n12699), .op(n11860) );
  nor3_1 U11707 ( .ip1(n12231), .ip2(n13835), .ip3(n11859), .op(n12310) );
  or2_1 U11708 ( .ip1(n11860), .ip2(n12310), .op(n11862) );
  nand2_1 U11709 ( .ip1(m1Inputs[57]), .ip2(n11974), .op(n12229) );
  or2_1 U11710 ( .ip1(n12229), .ip2(n12310), .op(n11861) );
  nand2_1 U11711 ( .ip1(n11862), .ip2(n11861), .op(n12309) );
  nor2_1 U11712 ( .ip1(n12126), .ip2(n14188), .op(n12311) );
  xor2_1 U11713 ( .ip1(n12309), .ip2(n12311), .op(n12394) );
  nand2_1 U11714 ( .ip1(m1Inputs[54]), .ip2(n4627), .op(n11864) );
  nor3_1 U11715 ( .ip1(n12155), .ip2(n14384), .ip3(n11863), .op(n12305) );
  or2_1 U11716 ( .ip1(n11864), .ip2(n12305), .op(n11866) );
  nand2_1 U11717 ( .ip1(m1Inputs[55]), .ip2(n12981), .op(n12236) );
  or2_1 U11718 ( .ip1(n12236), .ip2(n12305), .op(n11865) );
  nand2_1 U11719 ( .ip1(n11866), .ip2(n11865), .op(n12304) );
  nor2_1 U11720 ( .ip1(n12032), .ip2(n13579), .op(n12306) );
  xor2_1 U11721 ( .ip1(n12304), .ip2(n12306), .op(n12393) );
  inv_1 U11722 ( .ip(n11867), .op(n12412) );
  or2_1 U11723 ( .ip1(n11868), .ip2(n11870), .op(n11873) );
  inv_1 U11724 ( .ip(n11869), .op(n11871) );
  or2_1 U11725 ( .ip1(n11871), .ip2(n11870), .op(n11872) );
  nand2_1 U11726 ( .ip1(n11873), .ip2(n11872), .op(n12348) );
  or2_1 U11727 ( .ip1(n11874), .ip2(n11875), .op(n11878) );
  or2_1 U11728 ( .ip1(n11876), .ip2(n11875), .op(n11877) );
  nand2_1 U11729 ( .ip1(n11878), .ip2(n11877), .op(n12347) );
  nand2_1 U11730 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[59]), .op(
        n11880) );
  inv_1 U11731 ( .ip(m1Inputs[60]), .op(n12071) );
  nor3_1 U11732 ( .ip1(n13709), .ip2(n12071), .ip3(n11879), .op(n12322) );
  or2_1 U11733 ( .ip1(n11880), .ip2(n12322), .op(n11882) );
  nand2_1 U11734 ( .ip1(n12809), .ip2(m1Inputs[60]), .op(n12197) );
  or2_1 U11735 ( .ip1(n12197), .ip2(n12322), .op(n11881) );
  nand2_1 U11736 ( .ip1(n11882), .ip2(n11881), .op(n12320) );
  nand2_1 U11737 ( .ip1(column[53]), .ip2(n14768), .op(n12321) );
  xor2_1 U11738 ( .ip1(n12320), .ip2(n12321), .op(n12346) );
  fulladder U11739 ( .a(n11885), .b(n11884), .ci(n11883), .co(n12416), .s(
        n11893) );
  fulladder U11740 ( .a(n11888), .b(n11887), .ci(n11886), .co(n12415), .s(
        n11897) );
  fulladder U11741 ( .a(n11891), .b(n11890), .ci(n11889), .co(n12414), .s(
        n11900) );
  fulladder U11742 ( .a(n11894), .b(n11893), .ci(n11892), .co(n12428), .s(
        n11899) );
  fulladder U11743 ( .a(n11897), .b(n11896), .ci(n11895), .co(n12427), .s(
        n6872) );
  fulladder U11744 ( .a(n11900), .b(n11899), .ci(n11898), .co(n12437), .s(
        n6834) );
  inv_1 U11745 ( .ip(n11901), .op(n12435) );
  fulladder U11746 ( .a(n11904), .b(n11903), .ci(n11902), .co(n12434), .s(
        n11907) );
  fulladder U11747 ( .a(n11907), .b(n11906), .ci(n11905), .co(n12433), .s(
        \STAGE_1/M4/sum [4]) );
  nand2_1 U11748 ( .ip1(m1Inputs[62]), .ip2(\STAGE_1/weightReg [7]), .op(
        n11992) );
  nor2_1 U11749 ( .ip1(n14853), .ip2(n12063), .op(n11991) );
  nand2_1 U11750 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[60]), .op(
        n11990) );
  nand2_1 U11751 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[61]), .op(
        n11979) );
  inv_1 U11752 ( .ip(m1Inputs[63]), .op(n12130) );
  nor2_1 U11753 ( .ip1(n12130), .ip2(n14836), .op(n11978) );
  nand2_1 U11754 ( .ip1(n15025), .ip2(m1Inputs[57]), .op(n11977) );
  nor2_1 U11755 ( .ip1(n12130), .ip2(n12746), .op(n11921) );
  nand2_1 U11756 ( .ip1(m1Inputs[62]), .ip2(\STAGE_1/weightReg [6]), .op(
        n11920) );
  nand2_1 U11757 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[60]), .op(
        n11919) );
  nand2_1 U11758 ( .ip1(m1Inputs[55]), .ip2(\STAGE_1/weightReg [13]), .op(
        n11909) );
  nand2_1 U11759 ( .ip1(m1Inputs[57]), .ip2(n14847), .op(n11908) );
  xor2_1 U11760 ( .ip1(n11909), .ip2(n11908), .op(n11945) );
  nor2_1 U11761 ( .ip1(n13579), .ip2(n12155), .op(n12064) );
  inv_1 U11762 ( .ip(n12064), .op(n11940) );
  nand2_1 U11763 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[57]), .op(
        n12496) );
  nor2_1 U11764 ( .ip1(n11940), .ip2(n12496), .op(n11910) );
  or2_1 U11765 ( .ip1(n11945), .ip2(n11910), .op(n11912) );
  nor2_1 U11766 ( .ip1(n14842), .ip2(n12063), .op(n11944) );
  or2_1 U11767 ( .ip1(n11944), .ip2(n11910), .op(n11911) );
  nand2_1 U11768 ( .ip1(n11912), .ip2(n11911), .op(n12002) );
  nand2_1 U11769 ( .ip1(n14629), .ip2(m1Inputs[59]), .op(n11932) );
  nand2_1 U11770 ( .ip1(n13718), .ip2(m1Inputs[59]), .op(n11980) );
  nand2_1 U11771 ( .ip1(n14629), .ip2(m1Inputs[58]), .op(n11933) );
  nor2_1 U11772 ( .ip1(n11980), .ip2(n11933), .op(n11989) );
  or2_1 U11773 ( .ip1(n11932), .ip2(n11989), .op(n11915) );
  nand2_1 U11774 ( .ip1(n13718), .ip2(m1Inputs[58]), .op(n11913) );
  or2_1 U11775 ( .ip1(n11913), .ip2(n11989), .op(n11914) );
  nand2_1 U11776 ( .ip1(n11915), .ip2(n11914), .op(n11987) );
  nand2_1 U11777 ( .ip1(column[61]), .ip2(n14768), .op(n11916) );
  xor2_1 U11778 ( .ip1(n11987), .ip2(n11916), .op(n12001) );
  nor2_1 U11779 ( .ip1(n14853), .ip2(n12255), .op(n11918) );
  nand2_1 U11780 ( .ip1(n15025), .ip2(m1Inputs[56]), .op(n11939) );
  nand2_1 U11781 ( .ip1(m1Inputs[61]), .ip2(\STAGE_1/weightReg [7]), .op(
        n11917) );
  fulladder U11782 ( .a(n11918), .b(n11939), .ci(n11917), .co(n12000), .s(
        n12015) );
  fulladder U11783 ( .a(n11921), .b(n11920), .ci(n11919), .co(n11993), .s(
        n12014) );
  nand2_1 U11784 ( .ip1(n13718), .ip2(m1Inputs[60]), .op(n12501) );
  nor2_1 U11785 ( .ip1(n12501), .ip2(n12236), .op(n12094) );
  or2_1 U11786 ( .ip1(n13749), .ip2(n12064), .op(n11923) );
  or2_1 U11787 ( .ip1(m1Inputs[60]), .ip2(n12064), .op(n11922) );
  nand2_1 U11788 ( .ip1(n11923), .ip2(n11922), .op(n12093) );
  nand2_1 U11789 ( .ip1(n14816), .ip2(m1Inputs[52]), .op(n12095) );
  nor2_1 U11790 ( .ip1(n12093), .ip2(n12095), .op(n11924) );
  nor2_1 U11791 ( .ip1(n12094), .ip2(n11924), .op(n12023) );
  nand2_1 U11792 ( .ip1(m1Inputs[58]), .ip2(n14975), .op(n11926) );
  nand2_1 U11793 ( .ip1(m1Inputs[56]), .ip2(\STAGE_1/weightReg [10]), .op(
        n11925) );
  xor2_1 U11794 ( .ip1(n11926), .ip2(n11925), .op(n12034) );
  nor2_1 U11795 ( .ip1(n6503), .ip2(n12237), .op(n12194) );
  and3_1 U11796 ( .ip1(n14629), .ip2(m1Inputs[58]), .ip3(n12194), .op(n11927)
         );
  or2_1 U11797 ( .ip1(n12034), .ip2(n11927), .op(n11930) );
  nand2_1 U11798 ( .ip1(column[58]), .ip2(n13039), .op(n12033) );
  inv_1 U11799 ( .ip(n12033), .op(n11928) );
  or2_1 U11800 ( .ip1(n11928), .ip2(n11927), .op(n11929) );
  nand2_1 U11801 ( .ip1(n11930), .ip2(n11929), .op(n12022) );
  nand2_1 U11802 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[54]), .op(
        n12021) );
  inv_1 U11803 ( .ip(n11931), .op(n12011) );
  nand2_1 U11804 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[56]), .op(
        n11998) );
  nand2_1 U11805 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[58]), .op(
        n11951) );
  nor2_1 U11806 ( .ip1(n11932), .ip2(n11951), .op(n11947) );
  inv_1 U11807 ( .ip(n11933), .op(n11950) );
  or2_1 U11808 ( .ip1(m1Inputs[59]), .ip2(n11950), .op(n11935) );
  or2_1 U11809 ( .ip1(\STAGE_1/weightReg [9]), .ip2(n11950), .op(n11934) );
  nand2_1 U11810 ( .ip1(n11935), .ip2(n11934), .op(n11946) );
  nand2_1 U11811 ( .ip1(column[60]), .ip2(n13039), .op(n11948) );
  nor2_1 U11812 ( .ip1(n11946), .ip2(n11948), .op(n11936) );
  nor2_1 U11813 ( .ip1(n11947), .ip2(n11936), .op(n11997) );
  nand2_1 U11814 ( .ip1(n14816), .ip2(m1Inputs[55]), .op(n11996) );
  nand2_1 U11815 ( .ip1(m1Inputs[55]), .ip2(n15025), .op(n11938) );
  nand2_1 U11816 ( .ip1(m1Inputs[56]), .ip2(n14847), .op(n11937) );
  xor2_1 U11817 ( .ip1(n11938), .ip2(n11937), .op(n11963) );
  nor2_1 U11818 ( .ip1(n11940), .ip2(n11939), .op(n11941) );
  or2_1 U11819 ( .ip1(n11963), .ip2(n11941), .op(n11943) );
  nor2_1 U11820 ( .ip1(n14842), .ip2(n12255), .op(n11962) );
  or2_1 U11821 ( .ip1(n11962), .ip2(n11941), .op(n11942) );
  nand2_1 U11822 ( .ip1(n11943), .ip2(n11942), .op(n12019) );
  nand2_1 U11823 ( .ip1(m1Inputs[60]), .ip2(\STAGE_1/weightReg [7]), .op(
        n11966) );
  nor2_1 U11824 ( .ip1(n12130), .ip2(n14783), .op(n11965) );
  nand2_1 U11825 ( .ip1(m1Inputs[62]), .ip2(n12699), .op(n11964) );
  xnor2_1 U11826 ( .ip1(n11945), .ip2(n11944), .op(n12017) );
  nor2_1 U11827 ( .ip1(n11947), .ip2(n11946), .op(n11949) );
  xor2_1 U11828 ( .ip1(n11949), .ip2(n11948), .op(n11960) );
  nor2_1 U11829 ( .ip1(n12083), .ip2(n12231), .op(n12077) );
  nand2_1 U11830 ( .ip1(n11950), .ip2(n12077), .op(n11953) );
  inv_1 U11831 ( .ip(n11953), .op(n11956) );
  nand2_1 U11832 ( .ip1(m1Inputs[57]), .ip2(n14629), .op(n11952) );
  nand2_1 U11833 ( .ip1(n11952), .ip2(n11951), .op(n11954) );
  nand2_1 U11834 ( .ip1(n11954), .ip2(n11953), .op(n11973) );
  nand2_1 U11835 ( .ip1(column[59]), .ip2(n13039), .op(n11972) );
  nor2_1 U11836 ( .ip1(n11973), .ip2(n11972), .op(n11955) );
  nor2_1 U11837 ( .ip1(n11956), .ip2(n11955), .op(n11959) );
  nor2_1 U11838 ( .ip1(n14853), .ip2(n12066), .op(n11970) );
  nand2_1 U11839 ( .ip1(m1Inputs[61]), .ip2(n12981), .op(n11969) );
  nand2_1 U11840 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[59]), .op(
        n11968) );
  inv_1 U11841 ( .ip(n11957), .op(n12010) );
  fulladder U11842 ( .a(n11960), .b(n11959), .ci(n11958), .co(n12003), .s(
        n11961) );
  inv_1 U11843 ( .ip(n11961), .op(n12039) );
  xor2_1 U11844 ( .ip1(n11963), .ip2(n11962), .op(n12091) );
  fulladder U11845 ( .a(n11966), .b(n11965), .ci(n11964), .co(n12018), .s(
        n11967) );
  inv_1 U11846 ( .ip(n11967), .op(n12090) );
  fulladder U11847 ( .a(n11970), .b(n11969), .ci(n11968), .co(n11958), .s(
        n11971) );
  inv_1 U11848 ( .ip(n11971), .op(n12089) );
  xor2_1 U11849 ( .ip1(n11973), .ip2(n11972), .op(n12087) );
  nand2_1 U11850 ( .ip1(m1Inputs[62]), .ip2(n11974), .op(n12074) );
  nor2_1 U11851 ( .ip1(n13801), .ip2(n12130), .op(n12073) );
  nand2_1 U11852 ( .ip1(m1Inputs[59]), .ip2(\STAGE_1/weightReg [7]), .op(
        n12072) );
  inv_1 U11853 ( .ip(n11975), .op(n12086) );
  inv_1 U11854 ( .ip(m1Inputs[61]), .op(n12198) );
  nor2_1 U11855 ( .ip1(n12198), .ip2(n12746), .op(n12078) );
  nand2_1 U11856 ( .ip1(m1Inputs[51]), .ip2(n14976), .op(n12076) );
  inv_1 U11857 ( .ip(n11976), .op(n12485) );
  fulladder U11858 ( .a(n11979), .b(n11978), .ci(n11977), .co(n12477), .s(
        n11994) );
  nand4_1 U11859 ( .ip1(\STAGE_1/weightReg [11]), .ip2(\STAGE_1/weightReg [10]), .ip3(m1Inputs[60]), .ip4(m1Inputs[59]), .op(n12536) );
  inv_1 U11860 ( .ip(n12536), .op(n11981) );
  or2_1 U11861 ( .ip1(n11980), .ip2(n11981), .op(n11984) );
  nand2_1 U11862 ( .ip1(n14629), .ip2(m1Inputs[60]), .op(n11982) );
  or2_1 U11863 ( .ip1(n11982), .ip2(n11981), .op(n11983) );
  nand2_1 U11864 ( .ip1(n11984), .ip2(n11983), .op(n12534) );
  nand2_1 U11865 ( .ip1(column[62]), .ip2(n14768), .op(n11985) );
  xor2_1 U11866 ( .ip1(n12534), .ip2(n11985), .op(n12476) );
  nor2_1 U11867 ( .ip1(n14842), .ip2(n12237), .op(n12515) );
  nor2_1 U11868 ( .ip1(n13766), .ip2(n12198), .op(n12514) );
  nand2_1 U11869 ( .ip1(m1Inputs[63]), .ip2(\STAGE_1/weightReg [7]), .op(
        n12513) );
  inv_1 U11870 ( .ip(n11986), .op(n12475) );
  and3_1 U11871 ( .ip1(column[61]), .ip2(n15042), .ip3(n11987), .op(n11988) );
  nor2_1 U11872 ( .ip1(n11989), .ip2(n11988), .op(n12497) );
  fulladder U11873 ( .a(n11992), .b(n11991), .ci(n11990), .co(n12495), .s(
        n11995) );
  fulladder U11874 ( .a(n11995), .b(n11994), .ci(n11993), .co(n12492), .s(
        n12008) );
  fulladder U11875 ( .a(n11998), .b(n11997), .ci(n11996), .co(n12507), .s(
        n12005) );
  nor2_1 U11876 ( .ip1(n14902), .ip2(n12230), .op(n12512) );
  inv_1 U11877 ( .ip(m1Inputs[62]), .op(n12161) );
  nor2_1 U11878 ( .ip1(n6503), .ip2(n12161), .op(n12511) );
  nand2_1 U11879 ( .ip1(n14976), .ip2(m1Inputs[55]), .op(n12510) );
  inv_1 U11880 ( .ip(n11999), .op(n12506) );
  fulladder U11881 ( .a(n12002), .b(n12001), .ci(n12000), .co(n12505), .s(
        n12007) );
  fulladder U11882 ( .a(n12005), .b(n12004), .ci(n12003), .co(n12480), .s(
        n11957) );
  fulladder U11883 ( .a(n12008), .b(n12007), .ci(n12006), .co(n12483), .s(
        n11931) );
  fulladder U11884 ( .a(n12011), .b(n12010), .ci(n12009), .co(n11976), .s(
        n12012) );
  inv_1 U11885 ( .ip(n12012), .op(n12102) );
  fulladder U11886 ( .a(n12015), .b(n12014), .ci(n12013), .co(n12006), .s(
        n12016) );
  inv_1 U11887 ( .ip(n12016), .op(n12108) );
  fulladder U11888 ( .a(n12019), .b(n12018), .ci(n12017), .co(n12004), .s(
        n12020) );
  inv_1 U11889 ( .ip(n12020), .op(n12107) );
  fulladder U11890 ( .a(n12023), .b(n12022), .ci(n12021), .co(n12013), .s(
        n12024) );
  inv_1 U11891 ( .ip(n12024), .op(n12043) );
  nand2_1 U11892 ( .ip1(m1Inputs[59]), .ip2(n12981), .op(n12025) );
  nor3_1 U11893 ( .ip1(n12230), .ip2(n14836), .ip3(n12072), .op(n12029) );
  or2_1 U11894 ( .ip1(n12025), .ip2(n12029), .op(n12028) );
  nand2_1 U11895 ( .ip1(m1Inputs[58]), .ip2(\STAGE_1/weightReg [7]), .op(
        n12026) );
  or2_1 U11896 ( .ip1(n12026), .ip2(n12029), .op(n12027) );
  nand2_1 U11897 ( .ip1(n12028), .ip2(n12027), .op(n12060) );
  or2_1 U11898 ( .ip1(n12060), .ip2(n12029), .op(n12031) );
  nor2_1 U11899 ( .ip1(n12071), .ip2(n12746), .op(n12059) );
  or2_1 U11900 ( .ip1(n12059), .ip2(n12029), .op(n12030) );
  nand2_1 U11901 ( .ip1(n12031), .ip2(n12030), .op(n12146) );
  nand2_1 U11902 ( .ip1(m1Inputs[61]), .ip2(\STAGE_1/weightReg [4]), .op(
        n12152) );
  nor2_1 U11903 ( .ip1(n12032), .ip2(n14853), .op(n12151) );
  nand2_1 U11904 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[57]), .op(
        n12150) );
  xor2_1 U11905 ( .ip1(n12034), .ip2(n12033), .op(n12144) );
  inv_1 U11906 ( .ip(n12035), .op(n12042) );
  nor2_1 U11907 ( .ip1(n14340), .ip2(n12255), .op(n12046) );
  nor2_1 U11908 ( .ip1(n14902), .ip2(n12063), .op(n12045) );
  nor2_1 U11909 ( .ip1(n12083), .ip2(n12237), .op(n12056) );
  and2_1 U11910 ( .ip1(column[57]), .ip2(n13498), .op(n12055) );
  nand2_1 U11911 ( .ip1(column[56]), .ip2(n13039), .op(n12132) );
  inv_1 U11912 ( .ip(n12132), .op(n12054) );
  inv_1 U11913 ( .ip(n12036), .op(n12101) );
  fulladder U11914 ( .a(n12039), .b(n12038), .ci(n12037), .co(n12009), .s(
        n12040) );
  inv_1 U11915 ( .ip(n12040), .op(n12105) );
  fulladder U11916 ( .a(n12043), .b(n12042), .ci(n12041), .co(n12106), .s(
        n12175) );
  fulladder U11917 ( .a(n12046), .b(n12045), .ci(n12044), .co(n12041), .s(
        n12118) );
  nor2_1 U11918 ( .ip1(n12231), .ip2(n14836), .op(n12122) );
  and3_1 U11919 ( .ip1(m1Inputs[58]), .ip2(n4627), .ip3(n12122), .op(n12051)
         );
  nor2_1 U11920 ( .ip1(n12230), .ip2(n14289), .op(n12047) );
  or2_1 U11921 ( .ip1(\STAGE_1/weightReg [7]), .ip2(n12047), .op(n12049) );
  or2_1 U11922 ( .ip1(m1Inputs[57]), .ip2(n12047), .op(n12048) );
  nand2_1 U11923 ( .ip1(n12049), .ip2(n12048), .op(n12050) );
  nor2_1 U11924 ( .ip1(n12051), .ip2(n12050), .op(n12142) );
  or2_1 U11925 ( .ip1(n12142), .ip2(n12051), .op(n12053) );
  nor2_1 U11926 ( .ip1(n12248), .ip2(n12746), .op(n12141) );
  or2_1 U11927 ( .ip1(n12141), .ip2(n12051), .op(n12052) );
  nand2_1 U11928 ( .ip1(n12053), .ip2(n12052), .op(n12185) );
  nor2_1 U11929 ( .ip1(n13570), .ip2(n12130), .op(n12191) );
  nand2_1 U11930 ( .ip1(m1Inputs[50]), .ip2(n14816), .op(n12190) );
  fulladder U11931 ( .a(n12056), .b(n12055), .ci(n12054), .co(n12044), .s(
        n12057) );
  inv_1 U11932 ( .ip(n12057), .op(n12183) );
  inv_1 U11933 ( .ip(n12058), .op(n12117) );
  xor2_1 U11934 ( .ip1(n12060), .ip2(n12059), .op(n12188) );
  nand2_1 U11935 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[52]), .op(
        n12067) );
  nand2_1 U11936 ( .ip1(m1Inputs[55]), .ip2(\STAGE_1/weightReg [10]), .op(
        n12062) );
  nand2_1 U11937 ( .ip1(n13718), .ip2(m1Inputs[54]), .op(n12061) );
  nand2_1 U11938 ( .ip1(n12062), .ip2(n12061), .op(n12065) );
  nor2_1 U11939 ( .ip1(n13594), .ip2(n12063), .op(n12079) );
  nand2_1 U11940 ( .ip1(n12079), .ip2(n12064), .op(n12097) );
  nand2_1 U11941 ( .ip1(n12065), .ip2(n12097), .op(n12068) );
  nor3_1 U11942 ( .ip1(n14340), .ip2(n12066), .ip3(n12068), .op(n12098) );
  or2_1 U11943 ( .ip1(n12067), .ip2(n12098), .op(n12070) );
  or2_1 U11944 ( .ip1(n12068), .ip2(n12098), .op(n12069) );
  nand2_1 U11945 ( .ip1(n12070), .ip2(n12069), .op(n12187) );
  nor2_1 U11946 ( .ip1(n12071), .ip2(n14783), .op(n12195) );
  nand2_1 U11947 ( .ip1(m1Inputs[49]), .ip2(n14976), .op(n12193) );
  fulladder U11948 ( .a(n12074), .b(n12073), .ci(n12072), .co(n11975), .s(
        n12075) );
  inv_1 U11949 ( .ip(n12075), .op(n12115) );
  fulladder U11950 ( .a(n12078), .b(n12077), .ci(n12076), .co(n12085), .s(
        n12114) );
  nor2_1 U11951 ( .ip1(n14902), .ip2(n12255), .op(n12121) );
  or2_1 U11952 ( .ip1(m1Inputs[53]), .ip2(n12079), .op(n12081) );
  or2_1 U11953 ( .ip1(n14847), .ip2(n12079), .op(n12080) );
  nand2_1 U11954 ( .ip1(n12081), .ip2(n12080), .op(n12136) );
  nor3_1 U11955 ( .ip1(n12136), .ip2(n12138), .ip3(n14340), .op(n12082) );
  nor2_1 U11956 ( .ip1(n13594), .ip2(n12255), .op(n12253) );
  and3_1 U11957 ( .ip1(\STAGE_1/weightReg [11]), .ip2(m1Inputs[54]), .ip3(
        n12253), .op(n12137) );
  or2_1 U11958 ( .ip1(n12082), .ip2(n12137), .op(n12120) );
  nor2_1 U11959 ( .ip1(n13854), .ip2(n12161), .op(n12133) );
  nor2_1 U11960 ( .ip1(n12083), .ip2(n12155), .op(n12131) );
  inv_1 U11961 ( .ip(n12084), .op(n12104) );
  fulladder U11962 ( .a(n12087), .b(n12086), .ci(n12085), .co(n12037), .s(
        n12088) );
  inv_1 U11963 ( .ip(n12088), .op(n12112) );
  fulladder U11964 ( .a(n12091), .b(n12090), .ci(n12089), .co(n12038), .s(
        n12092) );
  inv_1 U11965 ( .ip(n12092), .op(n12111) );
  nor2_1 U11966 ( .ip1(n12094), .ip2(n12093), .op(n12096) );
  xor2_1 U11967 ( .ip1(n12096), .ip2(n12095), .op(n12149) );
  inv_1 U11968 ( .ip(n12097), .op(n12099) );
  nor2_1 U11969 ( .ip1(n12099), .ip2(n12098), .op(n12148) );
  nor2_1 U11970 ( .ip1(n13854), .ip2(n12130), .op(n12154) );
  nand2_1 U11971 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[62]), .op(
        n12246) );
  nand2_1 U11972 ( .ip1(m1Inputs[51]), .ip2(n14816), .op(n12153) );
  fulladder U11973 ( .a(n12102), .b(n12101), .ci(n12100), .co(n12503), .s(
        n12443) );
  fulladder U11974 ( .a(n12105), .b(n12104), .ci(n12103), .co(n12100), .s(
        n12172) );
  fulladder U11975 ( .a(n12108), .b(n12107), .ci(n12106), .co(n12036), .s(
        n12109) );
  inv_1 U11976 ( .ip(n12109), .op(n12171) );
  fulladder U11977 ( .a(n12112), .b(n12111), .ci(n12110), .co(n12103), .s(
        n12179) );
  fulladder U11978 ( .a(n12115), .b(n12114), .ci(n12113), .co(n12173), .s(
        n12270) );
  fulladder U11979 ( .a(n12118), .b(n12117), .ci(n12116), .co(n12174), .s(
        n12269) );
  fulladder U11980 ( .a(n12121), .b(n12120), .ci(n12119), .co(n12113), .s(
        n12274) );
  nor3_1 U11981 ( .ip1(n12248), .ip2(n14289), .ip3(n12229), .op(n12127) );
  or2_1 U11982 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n12122), .op(n12124) );
  or2_1 U11983 ( .ip1(m1Inputs[59]), .ip2(n12122), .op(n12123) );
  nand2_1 U11984 ( .ip1(n12124), .ip2(n12123), .op(n12125) );
  nor2_1 U11985 ( .ip1(n12127), .ip2(n12125), .op(n12217) );
  or2_1 U11986 ( .ip1(n12217), .ip2(n12127), .op(n12129) );
  nor2_1 U11987 ( .ip1(n12126), .ip2(n14842), .op(n12216) );
  or2_1 U11988 ( .ip1(n12216), .ip2(n12127), .op(n12128) );
  nand2_1 U11989 ( .ip1(n12129), .ip2(n12128), .op(n12223) );
  nor2_1 U11990 ( .ip1(n13646), .ip2(n12130), .op(n12211) );
  nand2_1 U11991 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[54]), .op(
        n12210) );
  fulladder U11992 ( .a(n12133), .b(n12132), .ci(n12131), .co(n12119), .s(
        n12134) );
  inv_1 U11993 ( .ip(n12134), .op(n12221) );
  inv_1 U11994 ( .ip(n12135), .op(n12273) );
  nor2_1 U11995 ( .ip1(n12137), .ip2(n12136), .op(n12140) );
  nor2_1 U11996 ( .ip1(n12138), .ip2(n14340), .op(n12139) );
  xor2_1 U11997 ( .ip1(n12140), .ip2(n12139), .op(n12220) );
  xor2_1 U11998 ( .ip1(n12142), .ip2(n12141), .op(n12219) );
  nor2_1 U11999 ( .ip1(n12230), .ip2(n12746), .op(n12215) );
  nand2_1 U12000 ( .ip1(m1Inputs[48]), .ip2(n14976), .op(n12214) );
  inv_1 U12001 ( .ip(n12143), .op(n12178) );
  fulladder U12002 ( .a(n12146), .b(n12145), .ci(n12144), .co(n12035), .s(
        n12182) );
  fulladder U12003 ( .a(n12149), .b(n12148), .ci(n12147), .co(n12110), .s(
        n12181) );
  fulladder U12004 ( .a(n12152), .b(n12151), .ci(n12150), .co(n12145), .s(
        n12209) );
  fulladder U12005 ( .a(n12154), .b(n12246), .ci(n12153), .co(n12147), .s(
        n12208) );
  nor2_1 U12006 ( .ip1(n12155), .ip2(n12156), .op(n12238) );
  and2_1 U12007 ( .ip1(n12194), .ip2(n12238), .op(n12243) );
  nor2_1 U12008 ( .ip1(n12237), .ip2(n12156), .op(n12157) );
  or2_1 U12009 ( .ip1(m1Inputs[55]), .ip2(n12157), .op(n12159) );
  or2_1 U12010 ( .ip1(n14838), .ip2(n12157), .op(n12158) );
  nand2_1 U12011 ( .ip1(n12159), .ip2(n12158), .op(n12242) );
  nand2_1 U12012 ( .ip1(m1Inputs[50]), .ip2(n15028), .op(n12244) );
  nor2_1 U12013 ( .ip1(n12242), .ip2(n12244), .op(n12160) );
  nor2_1 U12014 ( .ip1(n12243), .ip2(n12160), .op(n12228) );
  nand2_1 U12015 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[61]), .op(
        n12162) );
  nand2_1 U12016 ( .ip1(n12809), .ip2(m1Inputs[61]), .op(n12200) );
  nor3_1 U12017 ( .ip1(n13709), .ip2(n12161), .ip3(n12200), .op(n12166) );
  or2_1 U12018 ( .ip1(n12162), .ip2(n12166), .op(n12165) );
  nand2_1 U12019 ( .ip1(n12809), .ip2(m1Inputs[62]), .op(n12163) );
  or2_1 U12020 ( .ip1(n12163), .ip2(n12166), .op(n12164) );
  nand2_1 U12021 ( .ip1(n12165), .ip2(n12164), .op(n12261) );
  or2_1 U12022 ( .ip1(n12261), .ip2(n12166), .op(n12169) );
  nand2_1 U12023 ( .ip1(column[55]), .ip2(n13039), .op(n12260) );
  inv_1 U12024 ( .ip(n12260), .op(n12167) );
  or2_1 U12025 ( .ip1(n12167), .ip2(n12166), .op(n12168) );
  nand2_1 U12026 ( .ip1(n12169), .ip2(n12168), .op(n12227) );
  nand2_1 U12027 ( .ip1(n15025), .ip2(m1Inputs[52]), .op(n12226) );
  fulladder U12028 ( .a(n12172), .b(n12171), .ci(n12170), .co(n12442), .s(
        n12447) );
  fulladder U12029 ( .a(n12175), .b(n12174), .ci(n12173), .co(n12084), .s(
        n12176) );
  inv_1 U12030 ( .ip(n12176), .op(n12264) );
  fulladder U12031 ( .a(n12179), .b(n12178), .ci(n12177), .co(n12170), .s(
        n12263) );
  fulladder U12032 ( .a(n12182), .b(n12181), .ci(n12180), .co(n12177), .s(
        n12267) );
  fulladder U12033 ( .a(n12185), .b(n12184), .ci(n12183), .co(n12058), .s(
        n12278) );
  fulladder U12034 ( .a(n12188), .b(n12187), .ci(n12186), .co(n12116), .s(
        n12189) );
  inv_1 U12035 ( .ip(n12189), .op(n12277) );
  fulladder U12036 ( .a(n12192), .b(n12191), .ci(n12190), .co(n12184), .s(
        n12281) );
  fulladder U12037 ( .a(n12195), .b(n12194), .ci(n12193), .co(n12186), .s(
        n12196) );
  inv_1 U12038 ( .ip(n12196), .op(n12280) );
  nand2_1 U12039 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[60]), .op(
        n12199) );
  nor3_1 U12040 ( .ip1(n13709), .ip2(n12198), .ip3(n12197), .op(n12203) );
  or2_1 U12041 ( .ip1(n12199), .ip2(n12203), .op(n12202) );
  or2_1 U12042 ( .ip1(n12200), .ip2(n12203), .op(n12201) );
  nand2_1 U12043 ( .ip1(n12202), .ip2(n12201), .op(n12315) );
  or2_1 U12044 ( .ip1(n12315), .ip2(n12203), .op(n12206) );
  nand2_1 U12045 ( .ip1(column[54]), .ip2(n13039), .op(n12314) );
  inv_1 U12046 ( .ip(n12314), .op(n12204) );
  or2_1 U12047 ( .ip1(n12204), .ip2(n12203), .op(n12205) );
  nand2_1 U12048 ( .ip1(n12206), .ip2(n12205), .op(n12303) );
  nand2_1 U12049 ( .ip1(m1Inputs[51]), .ip2(n15025), .op(n12302) );
  nand2_1 U12050 ( .ip1(n13718), .ip2(m1Inputs[52]), .op(n12301) );
  fulladder U12051 ( .a(n12209), .b(n12208), .ci(n12207), .co(n12180), .s(
        n12331) );
  fulladder U12052 ( .a(n12212), .b(n12211), .ci(n12210), .co(n12222), .s(
        n12213) );
  inv_1 U12053 ( .ip(n12213), .op(n12344) );
  fulladder U12054 ( .a(n12215), .b(n12253), .ci(n12214), .co(n12218), .s(
        n12343) );
  xor2_1 U12055 ( .ip1(n12217), .ip2(n12216), .op(n12342) );
  fulladder U12056 ( .a(n12220), .b(n12219), .ci(n12218), .co(n12272), .s(
        n12339) );
  fulladder U12057 ( .a(n12223), .b(n12222), .ci(n12221), .co(n12135), .s(
        n12224) );
  inv_1 U12058 ( .ip(n12224), .op(n12338) );
  inv_1 U12059 ( .ip(n12225), .op(n12330) );
  fulladder U12060 ( .a(n12228), .b(n12227), .ci(n12226), .co(n12207), .s(
        n12337) );
  nor3_1 U12061 ( .ip1(n12230), .ip2(n4624), .ip3(n12229), .op(n12350) );
  nor2_1 U12062 ( .ip1(n12231), .ip2(n12746), .op(n12232) );
  or2_1 U12063 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n12232), .op(n12234) );
  or2_1 U12064 ( .ip1(m1Inputs[58]), .ip2(n12232), .op(n12233) );
  nand2_1 U12065 ( .ip1(n12234), .ip2(n12233), .op(n12349) );
  nand2_1 U12066 ( .ip1(n14975), .ip2(m1Inputs[54]), .op(n12351) );
  nor2_1 U12067 ( .ip1(n12349), .ip2(n12351), .op(n12235) );
  nor2_1 U12068 ( .ip1(n12350), .ip2(n12235), .op(n12297) );
  nor3_1 U12069 ( .ip1(n12237), .ip2(n14368), .ip3(n12236), .op(n12283) );
  or2_1 U12070 ( .ip1(n13749), .ip2(n12238), .op(n12240) );
  or2_1 U12071 ( .ip1(m1Inputs[56]), .ip2(n12238), .op(n12239) );
  nand2_1 U12072 ( .ip1(n12240), .ip2(n12239), .op(n12282) );
  nand2_1 U12073 ( .ip1(m1Inputs[49]), .ip2(\STAGE_1/weightReg [13]), .op(
        n12284) );
  nor2_1 U12074 ( .ip1(n12282), .ip2(n12284), .op(n12241) );
  nor2_1 U12075 ( .ip1(n12283), .ip2(n12241), .op(n12296) );
  nor2_1 U12076 ( .ip1(n12243), .ip2(n12242), .op(n12245) );
  xor2_1 U12077 ( .ip1(n12245), .ip2(n12244), .op(n12295) );
  nor2_1 U12078 ( .ip1(n12247), .ip2(n12246), .op(n12354) );
  nor2_1 U12079 ( .ip1(n13082), .ip2(n12248), .op(n12249) );
  or2_1 U12080 ( .ip1(m1Inputs[62]), .ip2(n12249), .op(n12251) );
  or2_1 U12081 ( .ip1(n13803), .ip2(n12249), .op(n12250) );
  nand2_1 U12082 ( .ip1(n12251), .ip2(n12250), .op(n12353) );
  nand2_1 U12083 ( .ip1(m1Inputs[48]), .ip2(n14816), .op(n12355) );
  nor2_1 U12084 ( .ip1(n12353), .ip2(n12355), .op(n12252) );
  nor2_1 U12085 ( .ip1(n12354), .ip2(n12252), .op(n12300) );
  and2_1 U12086 ( .ip1(n12254), .ip2(n12253), .op(n12292) );
  nor2_1 U12087 ( .ip1(n13766), .ip2(n12255), .op(n12256) );
  or2_1 U12088 ( .ip1(m1Inputs[52]), .ip2(n12256), .op(n12258) );
  or2_1 U12089 ( .ip1(n14876), .ip2(n12256), .op(n12257) );
  nand2_1 U12090 ( .ip1(n12258), .ip2(n12257), .op(n12291) );
  nand2_1 U12091 ( .ip1(m1Inputs[50]), .ip2(n15025), .op(n12293) );
  nor2_1 U12092 ( .ip1(n12291), .ip2(n12293), .op(n12259) );
  nor2_1 U12093 ( .ip1(n12292), .ip2(n12259), .op(n12299) );
  xor2_1 U12094 ( .ip1(n12261), .ip2(n12260), .op(n12298) );
  fulladder U12095 ( .a(n12264), .b(n12263), .ci(n12262), .co(n12446), .s(
        n12451) );
  fulladder U12096 ( .a(n12267), .b(n12266), .ci(n12265), .co(n12262), .s(
        n12328) );
  fulladder U12097 ( .a(n12270), .b(n12269), .ci(n12268), .co(n12143), .s(
        n12271) );
  inv_1 U12098 ( .ip(n12271), .op(n12327) );
  fulladder U12099 ( .a(n12274), .b(n12273), .ci(n12272), .co(n12268), .s(
        n12275) );
  inv_1 U12100 ( .ip(n12275), .op(n12334) );
  fulladder U12101 ( .a(n12278), .b(n12277), .ci(n12276), .co(n12266), .s(
        n12333) );
  fulladder U12102 ( .a(n12281), .b(n12280), .ci(n12279), .co(n12276), .s(
        n12371) );
  nor2_1 U12103 ( .ip1(n12283), .ip2(n12282), .op(n12285) );
  xor2_1 U12104 ( .ip1(n12285), .ip2(n12284), .op(n12387) );
  or2_1 U12105 ( .ip1(n12286), .ip2(n12287), .op(n12290) );
  or2_1 U12106 ( .ip1(n12288), .ip2(n12287), .op(n12289) );
  nand2_1 U12107 ( .ip1(n12290), .ip2(n12289), .op(n12386) );
  nor2_1 U12108 ( .ip1(n12292), .ip2(n12291), .op(n12294) );
  xor2_1 U12109 ( .ip1(n12294), .ip2(n12293), .op(n12385) );
  fulladder U12110 ( .a(n12297), .b(n12296), .ci(n12295), .co(n12336), .s(
        n12382) );
  fulladder U12111 ( .a(n12300), .b(n12299), .ci(n12298), .co(n12335), .s(
        n12381) );
  fulladder U12112 ( .a(n12303), .b(n12302), .ci(n12301), .co(n12279), .s(
        n12379) );
  or2_1 U12113 ( .ip1(n12304), .ip2(n12305), .op(n12308) );
  or2_1 U12114 ( .ip1(n12306), .ip2(n12305), .op(n12307) );
  nand2_1 U12115 ( .ip1(n12308), .ip2(n12307), .op(n12362) );
  or2_1 U12116 ( .ip1(n12309), .ip2(n12310), .op(n12313) );
  or2_1 U12117 ( .ip1(n12311), .ip2(n12310), .op(n12312) );
  nand2_1 U12118 ( .ip1(n12313), .ip2(n12312), .op(n12361) );
  xor2_1 U12119 ( .ip1(n12315), .ip2(n12314), .op(n12360) );
  nor2_1 U12120 ( .ip1(n12317), .ip2(n12316), .op(n12318) );
  nor2_1 U12121 ( .ip1(n12319), .ip2(n12318), .op(n12359) );
  or2_1 U12122 ( .ip1(n12320), .ip2(n12322), .op(n12325) );
  inv_1 U12123 ( .ip(n12321), .op(n12323) );
  or2_1 U12124 ( .ip1(n12323), .ip2(n12322), .op(n12324) );
  nand2_1 U12125 ( .ip1(n12325), .ip2(n12324), .op(n12358) );
  nand2_1 U12126 ( .ip1(m1Inputs[51]), .ip2(n13718), .op(n12357) );
  fulladder U12127 ( .a(n12328), .b(n12327), .ci(n12326), .co(n12450), .s(
        n12455) );
  fulladder U12128 ( .a(n12331), .b(n12330), .ci(n12329), .co(n12265), .s(
        n12368) );
  fulladder U12129 ( .a(n12334), .b(n12333), .ci(n12332), .co(n12326), .s(
        n12367) );
  fulladder U12130 ( .a(n12337), .b(n12336), .ci(n12335), .co(n12329), .s(
        n12375) );
  fulladder U12131 ( .a(n12340), .b(n12339), .ci(n12338), .co(n12225), .s(
        n12341) );
  inv_1 U12132 ( .ip(n12341), .op(n12374) );
  fulladder U12133 ( .a(n12344), .b(n12343), .ci(n12342), .co(n12340), .s(
        n12345) );
  inv_1 U12134 ( .ip(n12345), .op(n12403) );
  fulladder U12135 ( .a(n12348), .b(n12347), .ci(n12346), .co(n12391), .s(
        n12411) );
  nor2_1 U12136 ( .ip1(n12350), .ip2(n12349), .op(n12352) );
  xor2_1 U12137 ( .ip1(n12352), .ip2(n12351), .op(n12390) );
  nor2_1 U12138 ( .ip1(n12354), .ip2(n12353), .op(n12356) );
  xor2_1 U12139 ( .ip1(n12356), .ip2(n12355), .op(n12389) );
  fulladder U12140 ( .a(n12359), .b(n12358), .ci(n12357), .co(n12377), .s(
        n12410) );
  fulladder U12141 ( .a(n12362), .b(n12361), .ci(n12360), .co(n12378), .s(
        n12409) );
  fulladder U12142 ( .a(n12365), .b(n12364), .ci(n12363), .co(n12408), .s(
        n12413) );
  fulladder U12143 ( .a(n12368), .b(n12367), .ci(n12366), .co(n12454), .s(
        n12459) );
  fulladder U12144 ( .a(n12371), .b(n12370), .ci(n12369), .co(n12332), .s(
        n12372) );
  inv_1 U12145 ( .ip(n12372), .op(n12399) );
  fulladder U12146 ( .a(n12375), .b(n12374), .ci(n12373), .co(n12366), .s(
        n12376) );
  inv_1 U12147 ( .ip(n12376), .op(n12398) );
  fulladder U12148 ( .a(n12379), .b(n12378), .ci(n12377), .co(n12369), .s(
        n12380) );
  inv_1 U12149 ( .ip(n12380), .op(n12406) );
  fulladder U12150 ( .a(n12383), .b(n12382), .ci(n12381), .co(n12370), .s(
        n12384) );
  inv_1 U12151 ( .ip(n12384), .op(n12405) );
  fulladder U12152 ( .a(n12387), .b(n12386), .ci(n12385), .co(n12383), .s(
        n12388) );
  inv_1 U12153 ( .ip(n12388), .op(n12422) );
  fulladder U12154 ( .a(n12391), .b(n12390), .ci(n12389), .co(n12402), .s(
        n12392) );
  inv_1 U12155 ( .ip(n12392), .op(n12421) );
  fulladder U12156 ( .a(n12395), .b(n12394), .ci(n12393), .co(n12420), .s(
        n11867) );
  inv_1 U12157 ( .ip(n12396), .op(n12458) );
  fulladder U12158 ( .a(n12399), .b(n12398), .ci(n12397), .co(n12396), .s(
        n12400) );
  inv_1 U12159 ( .ip(n12400), .op(n12463) );
  fulladder U12160 ( .a(n12403), .b(n12402), .ci(n12401), .co(n12373), .s(
        n12419) );
  fulladder U12161 ( .a(n12406), .b(n12405), .ci(n12404), .co(n12397), .s(
        n12407) );
  inv_1 U12162 ( .ip(n12407), .op(n12418) );
  fulladder U12163 ( .a(n12410), .b(n12409), .ci(n12408), .co(n12401), .s(
        n12426) );
  fulladder U12164 ( .a(n12413), .b(n12412), .ci(n12411), .co(n12425), .s(
        n12439) );
  fulladder U12165 ( .a(n12416), .b(n12415), .ci(n12414), .co(n12424), .s(
        n12429) );
  fulladder U12166 ( .a(n12419), .b(n12418), .ci(n12417), .co(n12462), .s(
        n12467) );
  fulladder U12167 ( .a(n12422), .b(n12421), .ci(n12420), .co(n12404), .s(
        n12423) );
  inv_1 U12168 ( .ip(n12423), .op(n12432) );
  fulladder U12169 ( .a(n12426), .b(n12425), .ci(n12424), .co(n12417), .s(
        n12431) );
  fulladder U12170 ( .a(n12429), .b(n12428), .ci(n12427), .co(n12430), .s(
        n12438) );
  fulladder U12171 ( .a(n12432), .b(n12431), .ci(n12430), .co(n12466), .s(
        n12471) );
  fulladder U12172 ( .a(n12435), .b(n12434), .ci(n12433), .co(n12436), .s(
        \STAGE_1/M4/sum [5]) );
  inv_1 U12173 ( .ip(n12436), .op(n12470) );
  fulladder U12174 ( .a(n12439), .b(n12438), .ci(n12437), .co(n12469), .s(
        n11901) );
  inv_1 U12175 ( .ip(n12440), .op(\STAGE_1/M4/sum [14]) );
  fulladder U12176 ( .a(n12443), .b(n12442), .ci(n12441), .co(n12502), .s(
        n12444) );
  inv_1 U12177 ( .ip(n12444), .op(\STAGE_1/M4/sum [13]) );
  fulladder U12178 ( .a(n12447), .b(n12446), .ci(n12445), .co(n12441), .s(
        n12448) );
  inv_1 U12179 ( .ip(n12448), .op(\STAGE_1/M4/sum [12]) );
  fulladder U12180 ( .a(n12451), .b(n12450), .ci(n12449), .co(n12445), .s(
        n12452) );
  inv_1 U12181 ( .ip(n12452), .op(\STAGE_1/M4/sum [11]) );
  fulladder U12182 ( .a(n12455), .b(n12454), .ci(n12453), .co(n12449), .s(
        n12456) );
  inv_1 U12183 ( .ip(n12456), .op(\STAGE_1/M4/sum [10]) );
  fulladder U12184 ( .a(n12459), .b(n12458), .ci(n12457), .co(n12453), .s(
        n12460) );
  inv_1 U12185 ( .ip(n12460), .op(\STAGE_1/M4/sum [9]) );
  fulladder U12186 ( .a(n12463), .b(n12462), .ci(n12461), .co(n12457), .s(
        n12464) );
  inv_1 U12187 ( .ip(n12464), .op(\STAGE_1/M4/sum [8]) );
  fulladder U12188 ( .a(n12467), .b(n12466), .ci(n12465), .co(n12461), .s(
        n12468) );
  inv_1 U12189 ( .ip(n12468), .op(\STAGE_1/M4/sum [7]) );
  fulladder U12190 ( .a(n12471), .b(n12470), .ci(n12469), .co(n12465), .s(
        n12472) );
  inv_1 U12191 ( .ip(n12472), .op(\STAGE_1/M4/sum [6]) );
  nand2_1 U12192 ( .ip1(m1Inputs[63]), .ip2(n14975), .op(n12474) );
  nand2_1 U12193 ( .ip1(m1Inputs[57]), .ip2(\STAGE_1/weightReg [14]), .op(
        n12473) );
  xor2_1 U12194 ( .ip1(n12474), .ip2(n12473), .op(n12479) );
  fulladder U12195 ( .a(n12477), .b(n12476), .ci(n12475), .co(n12478), .s(
        n12494) );
  xor2_1 U12196 ( .ip1(n12479), .ip2(n12478), .op(n12489) );
  fulladder U12197 ( .a(n12482), .b(n12481), .ci(n12480), .co(n12487), .s(
        n12484) );
  fulladder U12198 ( .a(n12485), .b(n12484), .ci(n12483), .co(n12486), .s(
        n12504) );
  xor2_1 U12199 ( .ip1(n12487), .ip2(n12486), .op(n12488) );
  xor2_1 U12200 ( .ip1(n12489), .ip2(n12488), .op(n12491) );
  nand2_1 U12201 ( .ip1(m1Inputs[59]), .ip2(n15025), .op(n12490) );
  xor2_1 U12202 ( .ip1(n12491), .ip2(n12490), .op(n12533) );
  fulladder U12203 ( .a(n12494), .b(n12493), .ci(n12492), .co(n12499), .s(
        n12482) );
  fulladder U12204 ( .a(n12497), .b(n12496), .ci(n12495), .co(n12498), .s(
        n12493) );
  xor2_1 U12205 ( .ip1(n12499), .ip2(n12498), .op(n12500) );
  xor2_1 U12206 ( .ip1(n12501), .ip2(n12500), .op(n12529) );
  fulladder U12207 ( .a(n12504), .b(n12503), .ci(n12502), .co(n12509), .s(
        n12440) );
  fulladder U12208 ( .a(n12507), .b(n12506), .ci(n12505), .co(n12508), .s(
        n12481) );
  xor2_1 U12209 ( .ip1(n12509), .ip2(n12508), .op(n12519) );
  fulladder U12210 ( .a(n12512), .b(n12511), .ci(n12510), .co(n12517), .s(
        n11999) );
  fulladder U12211 ( .a(n12515), .b(n12514), .ci(n12513), .co(n12516), .s(
        n11986) );
  xor2_1 U12212 ( .ip1(n12517), .ip2(n12516), .op(n12518) );
  xor2_1 U12213 ( .ip1(n12519), .ip2(n12518), .op(n12527) );
  nand2_1 U12214 ( .ip1(m1Inputs[62]), .ip2(n14994), .op(n12521) );
  nand2_1 U12215 ( .ip1(m1Inputs[56]), .ip2(n14976), .op(n12520) );
  xor2_1 U12216 ( .ip1(n12521), .ip2(n12520), .op(n12525) );
  nand2_1 U12217 ( .ip1(m1Inputs[58]), .ip2(n15028), .op(n12523) );
  nand2_1 U12218 ( .ip1(m1Inputs[61]), .ip2(n14629), .op(n12522) );
  xor2_1 U12219 ( .ip1(n12523), .ip2(n12522), .op(n12524) );
  xor2_1 U12220 ( .ip1(n12525), .ip2(n12524), .op(n12526) );
  xor2_1 U12221 ( .ip1(n12527), .ip2(n12526), .op(n12528) );
  xor2_1 U12222 ( .ip1(n12529), .ip2(n12528), .op(n12531) );
  nand2_1 U12223 ( .ip1(n15042), .ip2(column[63]), .op(n12530) );
  xor2_1 U12224 ( .ip1(n12531), .ip2(n12530), .op(n12532) );
  xor2_1 U12225 ( .ip1(n12533), .ip2(n12532), .op(n12538) );
  nand3_1 U12226 ( .ip1(column[62]), .ip2(n15042), .ip3(n12534), .op(n12535)
         );
  nand2_1 U12227 ( .ip1(n12536), .ip2(n12535), .op(n12537) );
  xor2_1 U12228 ( .ip1(n12538), .ip2(n12537), .op(\STAGE_1/M4/sum [15]) );
  or2_1 U12229 ( .ip1(n12539), .ip2(n12541), .op(n12544) );
  inv_1 U12230 ( .ip(n12540), .op(n12542) );
  or2_1 U12231 ( .ip1(n12542), .ip2(n12541), .op(n12543) );
  nand2_1 U12232 ( .ip1(n12544), .ip2(n12543), .op(n13191) );
  or2_1 U12233 ( .ip1(n12545), .ip2(n12546), .op(n12549) );
  or2_1 U12234 ( .ip1(n12547), .ip2(n12546), .op(n12548) );
  nand2_1 U12235 ( .ip1(n12549), .ip2(n12548), .op(n13190) );
  nand2_1 U12236 ( .ip1(m1Inputs[67]), .ip2(n14975), .op(n13189) );
  fulladder U12237 ( .a(n12552), .b(n12551), .ci(n12550), .co(n13225), .s(
        n12587) );
  fulladder U12238 ( .a(n12555), .b(n12554), .ci(n12553), .co(n13224), .s(
        n12588) );
  nor2_1 U12239 ( .ip1(n12557), .ip2(n12556), .op(n12558) );
  nor2_1 U12240 ( .ip1(n12559), .ip2(n12558), .op(n13208) );
  or2_1 U12241 ( .ip1(n12560), .ip2(n12561), .op(n12564) );
  or2_1 U12242 ( .ip1(n12562), .ip2(n12561), .op(n12563) );
  nand2_1 U12243 ( .ip1(n12564), .ip2(n12563), .op(n13207) );
  nand2_1 U12244 ( .ip1(n4672), .ip2(m1Inputs[73]), .op(n12566) );
  nor3_1 U12245 ( .ip1(n13854), .ip2(n12959), .ip3(n12565), .op(n13151) );
  or2_1 U12246 ( .ip1(n12566), .ip2(n13151), .op(n12568) );
  nand2_1 U12247 ( .ip1(n13707), .ip2(m1Inputs[74]), .op(n13033) );
  or2_1 U12248 ( .ip1(n13033), .ip2(n13151), .op(n12567) );
  nand2_1 U12249 ( .ip1(n12568), .ip2(n12567), .op(n13149) );
  nand2_1 U12250 ( .ip1(column[67]), .ip2(n13039), .op(n13150) );
  xor2_1 U12251 ( .ip1(n13149), .ip2(n13150), .op(n13206) );
  nand2_1 U12252 ( .ip1(m1Inputs[68]), .ip2(\STAGE_1/weightReg [7]), .op(
        n12570) );
  and3_1 U12253 ( .ip1(n4627), .ip2(m1Inputs[69]), .ip3(n12569), .op(n13161)
         );
  or2_1 U12254 ( .ip1(n12570), .ip2(n13161), .op(n12572) );
  nand2_1 U12255 ( .ip1(n13749), .ip2(m1Inputs[69]), .op(n13044) );
  or2_1 U12256 ( .ip1(n13044), .ip2(n13161), .op(n12571) );
  nand2_1 U12257 ( .ip1(n12572), .ip2(n12571), .op(n13160) );
  nor2_1 U12258 ( .ip1(n13050), .ip2(n13766), .op(n13162) );
  xor2_1 U12259 ( .ip1(n13160), .ip2(n13162), .op(n13204) );
  nand2_1 U12260 ( .ip1(m1Inputs[70]), .ip2(\STAGE_1/weightReg [5]), .op(
        n12574) );
  inv_1 U12261 ( .ip(m1Inputs[71]), .op(n12982) );
  nor3_1 U12262 ( .ip1(n12982), .ip2(n13835), .ip3(n12573), .op(n13168) );
  or2_1 U12263 ( .ip1(n12574), .ip2(n13168), .op(n12576) );
  nand2_1 U12264 ( .ip1(m1Inputs[71]), .ip2(\STAGE_1/weightReg [4]), .op(
        n13070) );
  or2_1 U12265 ( .ip1(n13070), .ip2(n13168), .op(n12575) );
  nand2_1 U12266 ( .ip1(n12576), .ip2(n12575), .op(n13167) );
  nor2_1 U12267 ( .ip1(n13076), .ip2(n13594), .op(n13169) );
  xor2_1 U12268 ( .ip1(n13167), .ip2(n13169), .op(n13203) );
  nand2_1 U12269 ( .ip1(n13614), .ip2(m1Inputs[72]), .op(n12579) );
  and3_1 U12270 ( .ip1(n12578), .ip2(m1Inputs[75]), .ip3(n12577), .op(n13156)
         );
  or2_1 U12271 ( .ip1(n12579), .ip2(n13156), .op(n12581) );
  nand2_1 U12272 ( .ip1(\STAGE_1/weightReg [0]), .ip2(m1Inputs[75]), .op(
        n12920) );
  or2_1 U12273 ( .ip1(n12920), .ip2(n13156), .op(n12580) );
  nand2_1 U12274 ( .ip1(n12581), .ip2(n12580), .op(n13155) );
  nor2_1 U12275 ( .ip1(n12964), .ip2(n13579), .op(n13157) );
  xor2_1 U12276 ( .ip1(n13155), .ip2(n13157), .op(n13202) );
  inv_1 U12277 ( .ip(n12582), .op(n13237) );
  fulladder U12278 ( .a(n12585), .b(n12584), .ci(n12583), .co(n13236), .s(
        n5995) );
  fulladder U12279 ( .a(n12588), .b(n12587), .ci(n12586), .co(n13246), .s(
        n6026) );
  inv_1 U12280 ( .ip(n12589), .op(n13244) );
  fulladder U12281 ( .a(n12592), .b(n12591), .ci(n12590), .co(n13243), .s(
        n12595) );
  fulladder U12282 ( .a(n12595), .b(n12594), .ci(n12593), .co(n13242), .s(
        \STAGE_1/M5/sum [2]) );
  inv_1 U12283 ( .ip(m1Inputs[76]), .op(n13004) );
  nor2_1 U12284 ( .ip1(n13766), .ip2(n13004), .op(n12637) );
  inv_1 U12285 ( .ip(m1Inputs[78]), .op(n12810) );
  nor2_1 U12286 ( .ip1(n12810), .ip2(n14368), .op(n12636) );
  nand2_1 U12287 ( .ip1(n14976), .ip2(m1Inputs[70]), .op(n12635) );
  inv_1 U12288 ( .ip(n12596), .op(n12645) );
  nor2_1 U12289 ( .ip1(n14902), .ip2(n13081), .op(n12633) );
  inv_1 U12290 ( .ip(m1Inputs[77]), .op(n12874) );
  nor2_1 U12291 ( .ip1(n6503), .ip2(n12874), .op(n12632) );
  nand2_1 U12292 ( .ip1(m1Inputs[79]), .ip2(n12981), .op(n12631) );
  inv_1 U12293 ( .ip(n12597), .op(n12644) );
  inv_1 U12294 ( .ip(m1Inputs[79]), .op(n12837) );
  nor2_1 U12295 ( .ip1(n12837), .ip2(n12746), .op(n12614) );
  nand2_1 U12296 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[76]), .op(
        n12613) );
  nand2_1 U12297 ( .ip1(m1Inputs[78]), .ip2(n12981), .op(n12612) );
  nand2_1 U12298 ( .ip1(n14629), .ip2(m1Inputs[75]), .op(n12598) );
  nand2_1 U12299 ( .ip1(n13718), .ip2(m1Inputs[75]), .op(n12624) );
  nand2_1 U12300 ( .ip1(\STAGE_1/weightReg [10]), .ip2(m1Inputs[74]), .op(
        n12659) );
  nor2_1 U12301 ( .ip1(n12624), .ip2(n12659), .op(n12638) );
  or2_1 U12302 ( .ip1(n12598), .ip2(n12638), .op(n12601) );
  nand2_1 U12303 ( .ip1(n13718), .ip2(m1Inputs[74]), .op(n12599) );
  or2_1 U12304 ( .ip1(n12599), .ip2(n12638), .op(n12600) );
  nand2_1 U12305 ( .ip1(n12601), .ip2(n12600), .op(n12639) );
  inv_1 U12306 ( .ip(n12639), .op(n12603) );
  nand2_1 U12307 ( .ip1(column[77]), .ip2(n15042), .op(n12602) );
  mux2_1 U12308 ( .ip1(n12603), .ip2(n12639), .s(n12602), .op(n12655) );
  nor2_1 U12309 ( .ip1(n14373), .ip2(n13081), .op(n13321) );
  nand3_1 U12310 ( .ip1(n14847), .ip2(m1Inputs[71]), .ip3(n13321), .op(n12607)
         );
  nand2_1 U12311 ( .ip1(m1Inputs[71]), .ip2(\STAGE_1/weightReg [13]), .op(
        n12605) );
  nand2_1 U12312 ( .ip1(m1Inputs[73]), .ip2(n14847), .op(n12604) );
  xor2_1 U12313 ( .ip1(n12605), .ip2(n12604), .op(n12669) );
  nand3_1 U12314 ( .ip1(n14816), .ip2(m1Inputs[70]), .ip3(n12669), .op(n12606)
         );
  nand2_1 U12315 ( .ip1(n12607), .ip2(n12606), .op(n12654) );
  nor2_1 U12316 ( .ip1(n12874), .ip2(n14368), .op(n12610) );
  nor2_1 U12317 ( .ip1(n14902), .ip2(n13071), .op(n12671) );
  nand2_1 U12318 ( .ip1(n14976), .ip2(m1Inputs[69]), .op(n12609) );
  inv_1 U12319 ( .ip(n12608), .op(n12682) );
  fulladder U12320 ( .a(n12610), .b(n12671), .ci(n12609), .co(n12653), .s(
        n12611) );
  inv_1 U12321 ( .ip(n12611), .op(n12705) );
  fulladder U12322 ( .a(n12614), .b(n12613), .ci(n12612), .co(n12643), .s(
        n12704) );
  nand2_1 U12323 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[72]), .op(
        n12871) );
  nor2_1 U12324 ( .ip1(n12659), .ip2(n12871), .op(n12618) );
  nand2_1 U12325 ( .ip1(m1Inputs[74]), .ip2(n14975), .op(n12616) );
  nand2_1 U12326 ( .ip1(m1Inputs[72]), .ip2(\STAGE_1/weightReg [10]), .op(
        n12615) );
  xor2_1 U12327 ( .ip1(n12616), .ip2(n12615), .op(n12714) );
  and3_1 U12328 ( .ip1(column[74]), .ip2(n13498), .ip3(n12714), .op(n12617) );
  nor2_1 U12329 ( .ip1(n12618), .ip2(n12617), .op(n12718) );
  nand2_1 U12330 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[70]), .op(
        n12717) );
  nand2_1 U12331 ( .ip1(n13718), .ip2(m1Inputs[76]), .op(n13318) );
  nand2_1 U12332 ( .ip1(m1Inputs[71]), .ip2(n12981), .op(n12984) );
  nor2_1 U12333 ( .ip1(n13318), .ip2(n12984), .op(n12623) );
  nor2_1 U12334 ( .ip1(n14824), .ip2(n12982), .op(n12733) );
  or2_1 U12335 ( .ip1(n13749), .ip2(n12733), .op(n12620) );
  or2_1 U12336 ( .ip1(m1Inputs[76]), .ip2(n12733), .op(n12619) );
  nand2_1 U12337 ( .ip1(n12620), .ip2(n12619), .op(n12621) );
  or2_1 U12338 ( .ip1(n12623), .ip2(n12621), .op(n12774) );
  nor3_1 U12339 ( .ip1(n14842), .ip2(n12925), .ip3(n12774), .op(n12622) );
  nor2_1 U12340 ( .ip1(n12623), .ip2(n12622), .op(n12716) );
  nand4_1 U12341 ( .ip1(\STAGE_1/weightReg [11]), .ip2(\STAGE_1/weightReg [10]), .ip3(m1Inputs[76]), .ip4(m1Inputs[75]), .op(n13353) );
  inv_1 U12342 ( .ip(n13353), .op(n12625) );
  or2_1 U12343 ( .ip1(n12624), .ip2(n12625), .op(n12628) );
  nand2_1 U12344 ( .ip1(n14629), .ip2(m1Inputs[76]), .op(n12626) );
  or2_1 U12345 ( .ip1(n12626), .ip2(n12625), .op(n12627) );
  nand2_1 U12346 ( .ip1(n12628), .ip2(n12627), .op(n13351) );
  inv_1 U12347 ( .ip(n13351), .op(n12630) );
  nand2_1 U12348 ( .ip1(column[78]), .ip2(n13859), .op(n12629) );
  mux2_1 U12349 ( .ip1(n12630), .ip2(n13351), .s(n12629), .op(n13329) );
  nor2_1 U12350 ( .ip1(n14883), .ip2(n13071), .op(n13324) );
  nor2_1 U12351 ( .ip1(n13766), .ip2(n12874), .op(n13323) );
  nand2_1 U12352 ( .ip1(m1Inputs[79]), .ip2(\STAGE_1/weightReg [7]), .op(
        n13322) );
  fulladder U12353 ( .a(n12633), .b(n12632), .ci(n12631), .co(n13327), .s(
        n12597) );
  inv_1 U12354 ( .ip(n12634), .op(n13302) );
  fulladder U12355 ( .a(n12637), .b(n12636), .ci(n12635), .co(n13320), .s(
        n12596) );
  inv_1 U12356 ( .ip(n12638), .op(n12641) );
  nand3_1 U12357 ( .ip1(column[77]), .ip2(n15042), .ip3(n12639), .op(n12640)
         );
  nand2_1 U12358 ( .ip1(n12641), .ip2(n12640), .op(n13319) );
  inv_1 U12359 ( .ip(n12642), .op(n13301) );
  fulladder U12360 ( .a(n12645), .b(n12644), .ci(n12643), .co(n13300), .s(
        n12683) );
  inv_1 U12361 ( .ip(n12646), .op(n13299) );
  nor2_1 U12362 ( .ip1(n14842), .ip2(n12982), .op(n12658) );
  nor2_1 U12363 ( .ip1(n14340), .ip2(n13071), .op(n12657) );
  nand4_1 U12364 ( .ip1(\STAGE_1/weightReg [10]), .ip2(n14994), .ip3(
        m1Inputs[75]), .ip4(m1Inputs[74]), .op(n12652) );
  inv_1 U12365 ( .ip(n12652), .op(n12647) );
  or2_1 U12366 ( .ip1(n12659), .ip2(n12647), .op(n12650) );
  nand2_1 U12367 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[75]), .op(
        n12648) );
  or2_1 U12368 ( .ip1(n12648), .ip2(n12647), .op(n12649) );
  nand2_1 U12369 ( .ip1(n12650), .ip2(n12649), .op(n12667) );
  nand3_1 U12370 ( .ip1(column[76]), .ip2(n15042), .ip3(n12667), .op(n12651)
         );
  nand2_1 U12371 ( .ip1(n12652), .ip2(n12651), .op(n12656) );
  nor2_1 U12372 ( .ip1(n14902), .ip2(n12959), .op(n13332) );
  nor2_1 U12373 ( .ip1(n6504), .ip2(n12810), .op(n13331) );
  nand2_1 U12374 ( .ip1(n14976), .ip2(m1Inputs[71]), .op(n13330) );
  fulladder U12375 ( .a(n12655), .b(n12654), .ci(n12653), .co(n13309), .s(
        n12608) );
  fulladder U12376 ( .a(n12658), .b(n12657), .ci(n12656), .co(n13311), .s(
        n12679) );
  nand2_1 U12377 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[73]), .op(
        n12755) );
  nor2_1 U12378 ( .ip1(n12659), .ip2(n12755), .op(n12665) );
  nand2_1 U12379 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[74]), .op(
        n12660) );
  or2_1 U12380 ( .ip1(n12660), .ip2(n12665), .op(n12663) );
  nand2_1 U12381 ( .ip1(n14629), .ip2(m1Inputs[73]), .op(n12661) );
  or2_1 U12382 ( .ip1(n12661), .ip2(n12665), .op(n12662) );
  nand2_1 U12383 ( .ip1(n12663), .ip2(n12662), .op(n12698) );
  and3_1 U12384 ( .ip1(column[75]), .ip2(n15042), .ip3(n12698), .op(n12664) );
  nor2_1 U12385 ( .ip1(n12665), .ip2(n12664), .op(n12686) );
  nand2_1 U12386 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[75]), .op(
        n12694) );
  nor2_1 U12387 ( .ip1(n14853), .ip2(n12925), .op(n12693) );
  nand2_1 U12388 ( .ip1(m1Inputs[77]), .ip2(n12981), .op(n12692) );
  nand2_1 U12389 ( .ip1(column[76]), .ip2(n13039), .op(n12666) );
  xor2_1 U12390 ( .ip1(n12667), .ip2(n12666), .op(n12684) );
  inv_1 U12391 ( .ip(n12668), .op(n12678) );
  nor2_1 U12392 ( .ip1(n14842), .ip2(n13045), .op(n12670) );
  xor2_1 U12393 ( .ip1(n12670), .ip2(n12669), .op(n12702) );
  nand3_1 U12394 ( .ip1(n14847), .ip2(m1Inputs[71]), .ip3(n12671), .op(n12675)
         );
  nand2_1 U12395 ( .ip1(m1Inputs[71]), .ip2(n15025), .op(n12673) );
  nand2_1 U12396 ( .ip1(m1Inputs[72]), .ip2(n14847), .op(n12672) );
  xor2_1 U12397 ( .ip1(n12673), .ip2(n12672), .op(n12688) );
  nand3_1 U12398 ( .ip1(n14816), .ip2(n12688), .ip3(m1Inputs[69]), .op(n12674)
         );
  nand2_1 U12399 ( .ip1(n12675), .ip2(n12674), .op(n12701) );
  nor2_1 U12400 ( .ip1(n13004), .ip2(n14384), .op(n12691) );
  nor2_1 U12401 ( .ip1(n12810), .ip2(n12746), .op(n12690) );
  nand2_1 U12402 ( .ip1(m1Inputs[79]), .ip2(\STAGE_1/weightReg [4]), .op(
        n12689) );
  inv_1 U12403 ( .ip(n12676), .op(n13293) );
  fulladder U12404 ( .a(n12679), .b(n12678), .ci(n12677), .co(n13297), .s(
        n12680) );
  inv_1 U12405 ( .ip(n12680), .op(n12723) );
  fulladder U12406 ( .a(n12683), .b(n12682), .ci(n12681), .co(n13294), .s(
        n12722) );
  fulladder U12407 ( .a(n12686), .b(n12685), .ci(n12684), .co(n12668), .s(
        n12766) );
  nor2_1 U12408 ( .ip1(n14842), .ip2(n12999), .op(n12687) );
  xor2_1 U12409 ( .ip1(n12688), .ip2(n12687), .op(n12772) );
  fulladder U12410 ( .a(n12691), .b(n12690), .ci(n12689), .co(n12700), .s(
        n12771) );
  fulladder U12411 ( .a(n12694), .b(n12693), .ci(n12692), .co(n12685), .s(
        n12695) );
  inv_1 U12412 ( .ip(n12695), .op(n12770) );
  inv_1 U12413 ( .ip(n12696), .op(n12765) );
  nand2_1 U12414 ( .ip1(column[75]), .ip2(n14768), .op(n12697) );
  xor2_1 U12415 ( .ip1(n12698), .ip2(n12697), .op(n12769) );
  nand2_1 U12416 ( .ip1(m1Inputs[77]), .ip2(n12699), .op(n12757) );
  nor2_1 U12417 ( .ip1(n12845), .ip2(n14853), .op(n12756) );
  nor2_1 U12418 ( .ip1(n13082), .ip2(n12837), .op(n12753) );
  nand2_1 U12419 ( .ip1(m1Inputs[78]), .ip2(\STAGE_1/weightReg [4]), .op(
        n12752) );
  nand2_1 U12420 ( .ip1(m1Inputs[75]), .ip2(\STAGE_1/weightReg [7]), .op(
        n12751) );
  fulladder U12421 ( .a(n12702), .b(n12701), .ci(n12700), .co(n12677), .s(
        n12785) );
  fulladder U12422 ( .a(n12705), .b(n12704), .ci(n12703), .co(n12681), .s(
        n12706) );
  inv_1 U12423 ( .ip(n12706), .op(n12784) );
  nor3_1 U12424 ( .ip1(n12959), .ip2(n14289), .ip3(n12751), .op(n12712) );
  inv_1 U12425 ( .ip(n12712), .op(n12710) );
  nand2_1 U12426 ( .ip1(m1Inputs[75]), .ip2(n12981), .op(n12708) );
  nand2_1 U12427 ( .ip1(m1Inputs[74]), .ip2(\STAGE_1/weightReg [7]), .op(
        n12707) );
  nand2_1 U12428 ( .ip1(n12708), .ip2(n12707), .op(n12709) );
  nand2_1 U12429 ( .ip1(n12710), .ip2(n12709), .op(n12736) );
  nor3_1 U12430 ( .ip1(n13004), .ip2(n13835), .ip3(n12736), .op(n12711) );
  nor2_1 U12431 ( .ip1(n12712), .ip2(n12711), .op(n12796) );
  nand2_1 U12432 ( .ip1(m1Inputs[77]), .ip2(\STAGE_1/weightReg [4]), .op(
        n12802) );
  nor2_1 U12433 ( .ip1(n13050), .ip2(n14853), .op(n12801) );
  nand2_1 U12434 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[73]), .op(
        n12800) );
  nand2_1 U12435 ( .ip1(column[74]), .ip2(n13039), .op(n12713) );
  xor2_1 U12436 ( .ip1(n12714), .ip2(n12713), .op(n12794) );
  inv_1 U12437 ( .ip(n12715), .op(n12726) );
  fulladder U12438 ( .a(n12718), .b(n12717), .ci(n12716), .co(n12703), .s(
        n12719) );
  inv_1 U12439 ( .ip(n12719), .op(n12725) );
  nor2_1 U12440 ( .ip1(n14902), .ip2(n13045), .op(n12729) );
  nor2_1 U12441 ( .ip1(n14340), .ip2(n12999), .op(n12728) );
  and2_1 U12442 ( .ip1(column[73]), .ip2(n13498), .op(n12740) );
  nand2_1 U12443 ( .ip1(column[72]), .ip2(n14768), .op(n12838) );
  inv_1 U12444 ( .ip(n12838), .op(n12739) );
  nor2_1 U12445 ( .ip1(n13766), .ip2(n13071), .op(n12738) );
  inv_1 U12446 ( .ip(n12720), .op(n12782) );
  fulladder U12447 ( .a(n12723), .b(n12722), .ci(n12721), .co(n13292), .s(
        n12781) );
  fulladder U12448 ( .a(n12726), .b(n12725), .ci(n12724), .co(n12783), .s(
        n12861) );
  fulladder U12449 ( .a(n12729), .b(n12728), .ci(n12727), .co(n12724), .s(
        n12730) );
  inv_1 U12450 ( .ip(n12730), .op(n12825) );
  nor2_1 U12451 ( .ip1(n14340), .ip2(n12925), .op(n12735) );
  nand2_1 U12452 ( .ip1(m1Inputs[71]), .ip2(\STAGE_1/weightReg [10]), .op(
        n12732) );
  nand2_1 U12453 ( .ip1(n13718), .ip2(m1Inputs[70]), .op(n12731) );
  nand2_1 U12454 ( .ip1(n12732), .ip2(n12731), .op(n12734) );
  nor2_1 U12455 ( .ip1(n13594), .ip2(n13045), .op(n12759) );
  nand2_1 U12456 ( .ip1(n12733), .ip2(n12759), .op(n12776) );
  nand2_1 U12457 ( .ip1(n12734), .ip2(n12776), .op(n12777) );
  xor2_1 U12458 ( .ip1(n12735), .ip2(n12777), .op(n12868) );
  nand2_1 U12459 ( .ip1(m1Inputs[76]), .ip2(\STAGE_1/weightReg [4]), .op(
        n12873) );
  nor2_1 U12460 ( .ip1(n13076), .ip2(n14853), .op(n12872) );
  nor2_1 U12461 ( .ip1(n13004), .ip2(n12746), .op(n12737) );
  xor2_1 U12462 ( .ip1(n12737), .ip2(n12736), .op(n12866) );
  fulladder U12463 ( .a(n12740), .b(n12739), .ci(n12738), .co(n12727), .s(
        n12741) );
  inv_1 U12464 ( .ip(n12741), .op(n12865) );
  nor2_1 U12465 ( .ip1(n13081), .ip2(n14836), .op(n12830) );
  and3_1 U12466 ( .ip1(m1Inputs[74]), .ip2(n14835), .ip3(n12830), .op(n12747)
         );
  nor2_1 U12467 ( .ip1(n12959), .ip2(n14289), .op(n12742) );
  or2_1 U12468 ( .ip1(\STAGE_1/weightReg [7]), .ip2(n12742), .op(n12744) );
  or2_1 U12469 ( .ip1(m1Inputs[73]), .ip2(n12742), .op(n12743) );
  nand2_1 U12470 ( .ip1(n12744), .ip2(n12743), .op(n12745) );
  nor2_1 U12471 ( .ip1(n12747), .ip2(n12745), .op(n12849) );
  or2_1 U12472 ( .ip1(n12849), .ip2(n12747), .op(n12749) );
  inv_1 U12473 ( .ip(m1Inputs[75]), .op(n13034) );
  nor2_1 U12474 ( .ip1(n13034), .ip2(n12746), .op(n12848) );
  or2_1 U12475 ( .ip1(n12848), .ip2(n12747), .op(n12748) );
  nand2_1 U12476 ( .ip1(n12749), .ip2(n12748), .op(n12864) );
  nor2_1 U12477 ( .ip1(n13570), .ip2(n12837), .op(n12870) );
  nand2_1 U12478 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[77]), .op(
        n12957) );
  nand2_1 U12479 ( .ip1(m1Inputs[66]), .ip2(\STAGE_1/weightReg [14]), .op(
        n12869) );
  inv_1 U12480 ( .ip(n12750), .op(n12860) );
  fulladder U12481 ( .a(n12753), .b(n12752), .ci(n12751), .co(n12767), .s(
        n12754) );
  inv_1 U12482 ( .ip(n12754), .op(n12822) );
  fulladder U12483 ( .a(n12757), .b(n12756), .ci(n12755), .co(n12768), .s(
        n12758) );
  inv_1 U12484 ( .ip(n12758), .op(n12821) );
  nor2_1 U12485 ( .ip1(n14902), .ip2(n12999), .op(n12829) );
  or2_1 U12486 ( .ip1(m1Inputs[69]), .ip2(n12759), .op(n12761) );
  or2_1 U12487 ( .ip1(\STAGE_1/weightReg [11]), .ip2(n12759), .op(n12760) );
  nand2_1 U12488 ( .ip1(n12761), .ip2(n12760), .op(n12843) );
  nor3_1 U12489 ( .ip1(n12843), .ip2(n12845), .ip3(n14340), .op(n12762) );
  nor2_1 U12490 ( .ip1(n13594), .ip2(n12999), .op(n12926) );
  and3_1 U12491 ( .ip1(\STAGE_1/weightReg [11]), .ip2(m1Inputs[70]), .ip3(
        n12926), .op(n12844) );
  or2_1 U12492 ( .ip1(n12762), .ip2(n12844), .op(n12828) );
  nor2_1 U12493 ( .ip1(n13766), .ip2(n12982), .op(n12840) );
  nor2_1 U12494 ( .ip1(n13854), .ip2(n12810), .op(n12839) );
  inv_1 U12495 ( .ip(n12763), .op(n12788) );
  fulladder U12496 ( .a(n12766), .b(n12765), .ci(n12764), .co(n12721), .s(
        n12787) );
  fulladder U12497 ( .a(n12769), .b(n12768), .ci(n12767), .co(n12764), .s(
        n12792) );
  fulladder U12498 ( .a(n12772), .b(n12771), .ci(n12770), .co(n12696), .s(
        n12773) );
  inv_1 U12499 ( .ip(n12773), .op(n12791) );
  nor2_1 U12500 ( .ip1(n14842), .ip2(n12925), .op(n12775) );
  xor2_1 U12501 ( .ip1(n12775), .ip2(n12774), .op(n12799) );
  inv_1 U12502 ( .ip(n12776), .op(n12779) );
  nor3_1 U12503 ( .ip1(n14340), .ip2(n12925), .ip3(n12777), .op(n12778) );
  nor2_1 U12504 ( .ip1(n12779), .ip2(n12778), .op(n12798) );
  nor2_1 U12505 ( .ip1(n13854), .ip2(n12837), .op(n12804) );
  nand2_1 U12506 ( .ip1(n13614), .ip2(m1Inputs[78]), .op(n12919) );
  nand2_1 U12507 ( .ip1(m1Inputs[67]), .ip2(\STAGE_1/weightReg [14]), .op(
        n12803) );
  fulladder U12508 ( .a(n12782), .b(n12781), .ci(n12780), .co(n13313), .s(
        n13252) );
  fulladder U12509 ( .a(n12785), .b(n12784), .ci(n12783), .co(n12720), .s(
        n12853) );
  fulladder U12510 ( .a(n12788), .b(n12787), .ci(n12786), .co(n12780), .s(
        n12789) );
  inv_1 U12511 ( .ip(n12789), .op(n12852) );
  fulladder U12512 ( .a(n12792), .b(n12791), .ci(n12790), .co(n12786), .s(
        n12793) );
  inv_1 U12513 ( .ip(n12793), .op(n12857) );
  fulladder U12514 ( .a(n12796), .b(n12795), .ci(n12794), .co(n12715), .s(
        n12885) );
  fulladder U12515 ( .a(n12799), .b(n12798), .ci(n12797), .co(n12790), .s(
        n12884) );
  fulladder U12516 ( .a(n12802), .b(n12801), .ci(n12800), .co(n12795), .s(
        n12888) );
  fulladder U12517 ( .a(n12804), .b(n12919), .ci(n12803), .co(n12797), .s(
        n12887) );
  nor3_1 U12518 ( .ip1(n12982), .ip2(n12871), .ip3(n14368), .op(n12916) );
  nor2_1 U12519 ( .ip1(n13071), .ip2(n14368), .op(n12805) );
  or2_1 U12520 ( .ip1(m1Inputs[71]), .ip2(n12805), .op(n12807) );
  or2_1 U12521 ( .ip1(n14838), .ip2(n12805), .op(n12806) );
  nand2_1 U12522 ( .ip1(n12807), .ip2(n12806), .op(n12915) );
  nand2_1 U12523 ( .ip1(m1Inputs[66]), .ip2(\STAGE_1/weightReg [13]), .op(
        n12917) );
  nor2_1 U12524 ( .ip1(n12915), .ip2(n12917), .op(n12808) );
  nor2_1 U12525 ( .ip1(n12916), .ip2(n12808), .op(n12906) );
  nand2_1 U12526 ( .ip1(n4672), .ip2(m1Inputs[77]), .op(n12811) );
  nand2_1 U12527 ( .ip1(n12809), .ip2(m1Inputs[77]), .op(n12876) );
  nor3_1 U12528 ( .ip1(n13709), .ip2(n12810), .ip3(n12876), .op(n12815) );
  or2_1 U12529 ( .ip1(n12811), .ip2(n12815), .op(n12814) );
  nand2_1 U12530 ( .ip1(n13707), .ip2(m1Inputs[78]), .op(n12812) );
  or2_1 U12531 ( .ip1(n12812), .ip2(n12815), .op(n12813) );
  nand2_1 U12532 ( .ip1(n12814), .ip2(n12813), .op(n12932) );
  or2_1 U12533 ( .ip1(n12932), .ip2(n12815), .op(n12818) );
  nand2_1 U12534 ( .ip1(column[71]), .ip2(n13039), .op(n12931) );
  inv_1 U12535 ( .ip(n12931), .op(n12816) );
  or2_1 U12536 ( .ip1(n12816), .ip2(n12815), .op(n12817) );
  nand2_1 U12537 ( .ip1(n12818), .ip2(n12817), .op(n12905) );
  nand2_1 U12538 ( .ip1(n15025), .ip2(m1Inputs[68]), .op(n12904) );
  inv_1 U12539 ( .ip(n12819), .op(n12856) );
  fulladder U12540 ( .a(n12822), .b(n12821), .ci(n12820), .co(n12859), .s(
        n12938) );
  fulladder U12541 ( .a(n12825), .b(n12824), .ci(n12823), .co(n12750), .s(
        n12826) );
  inv_1 U12542 ( .ip(n12826), .op(n12937) );
  fulladder U12543 ( .a(n12829), .b(n12828), .ci(n12827), .co(n12820), .s(
        n12945) );
  nand2_1 U12544 ( .ip1(m1Inputs[73]), .ip2(\STAGE_1/weightReg [4]), .op(
        n12991) );
  nor3_1 U12545 ( .ip1(n13034), .ip2(n14289), .ip3(n12991), .op(n12834) );
  or2_1 U12546 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n12830), .op(n12832) );
  or2_1 U12547 ( .ip1(m1Inputs[75]), .ip2(n12830), .op(n12831) );
  nand2_1 U12548 ( .ip1(n12832), .ip2(n12831), .op(n12833) );
  nor2_1 U12549 ( .ip1(n12834), .ip2(n12833), .op(n12895) );
  or2_1 U12550 ( .ip1(n12895), .ip2(n12834), .op(n12836) );
  nor2_1 U12551 ( .ip1(n13076), .ip2(n14842), .op(n12894) );
  or2_1 U12552 ( .ip1(n12894), .ip2(n12834), .op(n12835) );
  nand2_1 U12553 ( .ip1(n12836), .ip2(n12835), .op(n12901) );
  nand2_1 U12554 ( .ip1(\STAGE_1/weightReg [3]), .ip2(m1Inputs[76]), .op(
        n13080) );
  nor2_1 U12555 ( .ip1(n13646), .ip2(n12837), .op(n12892) );
  nand2_1 U12556 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[70]), .op(
        n12891) );
  fulladder U12557 ( .a(n12840), .b(n12839), .ci(n12838), .co(n12827), .s(
        n12841) );
  inv_1 U12558 ( .ip(n12841), .op(n12899) );
  inv_1 U12559 ( .ip(n12842), .op(n12944) );
  nor2_1 U12560 ( .ip1(n12844), .ip2(n12843), .op(n12847) );
  nor2_1 U12561 ( .ip1(n12845), .ip2(n14340), .op(n12846) );
  xor2_1 U12562 ( .ip1(n12847), .ip2(n12846), .op(n12898) );
  xor2_1 U12563 ( .ip1(n12849), .ip2(n12848), .op(n12897) );
  nor2_1 U12564 ( .ip1(n12959), .ip2(n4624), .op(n12890) );
  nand2_1 U12565 ( .ip1(m1Inputs[64]), .ip2(n14976), .op(n12889) );
  inv_1 U12566 ( .ip(n12850), .op(n13251) );
  fulladder U12567 ( .a(n12853), .b(n12852), .ci(n12851), .co(n12850), .s(
        n12854) );
  inv_1 U12568 ( .ip(n12854), .op(n13256) );
  fulladder U12569 ( .a(n12857), .b(n12856), .ci(n12855), .co(n12851), .s(
        n12858) );
  inv_1 U12570 ( .ip(n12858), .op(n12935) );
  fulladder U12571 ( .a(n12861), .b(n12860), .ci(n12859), .co(n12763), .s(
        n12862) );
  inv_1 U12572 ( .ip(n12862), .op(n12934) );
  fulladder U12573 ( .a(n12865), .b(n12864), .ci(n12863), .co(n12823), .s(
        n12949) );
  fulladder U12574 ( .a(n12868), .b(n12867), .ci(n12866), .co(n12824), .s(
        n12948) );
  fulladder U12575 ( .a(n12870), .b(n12957), .ci(n12869), .co(n12863), .s(
        n12952) );
  fulladder U12576 ( .a(n12873), .b(n12872), .ci(n12871), .co(n12867), .s(
        n12951) );
  nand2_1 U12577 ( .ip1(n4672), .ip2(m1Inputs[76]), .op(n12875) );
  nand2_1 U12578 ( .ip1(n13707), .ip2(m1Inputs[76]), .op(n13006) );
  nor3_1 U12579 ( .ip1(n13709), .ip2(n12874), .ip3(n13006), .op(n12879) );
  or2_1 U12580 ( .ip1(n12875), .ip2(n12879), .op(n12878) );
  or2_1 U12581 ( .ip1(n12876), .ip2(n12879), .op(n12877) );
  nand2_1 U12582 ( .ip1(n12878), .ip2(n12877), .op(n12998) );
  or2_1 U12583 ( .ip1(n12998), .ip2(n12879), .op(n12882) );
  nand2_1 U12584 ( .ip1(column[70]), .ip2(n13039), .op(n12997) );
  inv_1 U12585 ( .ip(n12997), .op(n12880) );
  or2_1 U12586 ( .ip1(n12880), .ip2(n12879), .op(n12881) );
  nand2_1 U12587 ( .ip1(n12882), .ip2(n12881), .op(n12980) );
  nand2_1 U12588 ( .ip1(m1Inputs[67]), .ip2(\STAGE_1/weightReg [12]), .op(
        n12979) );
  nand2_1 U12589 ( .ip1(n13718), .ip2(m1Inputs[68]), .op(n12978) );
  fulladder U12590 ( .a(n12885), .b(n12884), .ci(n12883), .co(n12819), .s(
        n12941) );
  fulladder U12591 ( .a(n12888), .b(n12887), .ci(n12886), .co(n12883), .s(
        n13018) );
  fulladder U12592 ( .a(n12890), .b(n12926), .ci(n12889), .co(n12896), .s(
        n13031) );
  fulladder U12593 ( .a(n13080), .b(n12892), .ci(n12891), .co(n12900), .s(
        n12893) );
  inv_1 U12594 ( .ip(n12893), .op(n13030) );
  xor2_1 U12595 ( .ip1(n12895), .ip2(n12894), .op(n13029) );
  fulladder U12596 ( .a(n12898), .b(n12897), .ci(n12896), .co(n12943), .s(
        n13026) );
  fulladder U12597 ( .a(n12901), .b(n12900), .ci(n12899), .co(n12842), .s(
        n12902) );
  inv_1 U12598 ( .ip(n12902), .op(n13025) );
  inv_1 U12599 ( .ip(n12903), .op(n13017) );
  fulladder U12600 ( .a(n12906), .b(n12905), .ci(n12904), .co(n12886), .s(
        n13024) );
  nor3_1 U12601 ( .ip1(n12959), .ip2(n13835), .ip3(n12991), .op(n13057) );
  nor2_1 U12602 ( .ip1(n13081), .ip2(n4624), .op(n12907) );
  or2_1 U12603 ( .ip1(n11974), .ip2(n12907), .op(n12909) );
  or2_1 U12604 ( .ip1(m1Inputs[74]), .ip2(n12907), .op(n12908) );
  nand2_1 U12605 ( .ip1(n12909), .ip2(n12908), .op(n13056) );
  nand2_1 U12606 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[70]), .op(
        n13058) );
  nor2_1 U12607 ( .ip1(n13056), .ip2(n13058), .op(n12910) );
  nor2_1 U12608 ( .ip1(n13057), .ip2(n12910), .op(n12974) );
  nor3_1 U12609 ( .ip1(n13071), .ip2(n14368), .ip3(n12984), .op(n12954) );
  nor2_1 U12610 ( .ip1(n12982), .ip2(n14384), .op(n12911) );
  or2_1 U12611 ( .ip1(n13749), .ip2(n12911), .op(n12913) );
  or2_1 U12612 ( .ip1(m1Inputs[72]), .ip2(n12911), .op(n12912) );
  nand2_1 U12613 ( .ip1(n12913), .ip2(n12912), .op(n12953) );
  nand2_1 U12614 ( .ip1(m1Inputs[65]), .ip2(\STAGE_1/weightReg [13]), .op(
        n12955) );
  nor2_1 U12615 ( .ip1(n12953), .ip2(n12955), .op(n12914) );
  nor2_1 U12616 ( .ip1(n12954), .ip2(n12914), .op(n12973) );
  nor2_1 U12617 ( .ip1(n12916), .ip2(n12915), .op(n12918) );
  xor2_1 U12618 ( .ip1(n12918), .ip2(n12917), .op(n12972) );
  nor2_1 U12619 ( .ip1(n12920), .ip2(n12919), .op(n13061) );
  nor2_1 U12620 ( .ip1(n13082), .ip2(n13034), .op(n12921) );
  or2_1 U12621 ( .ip1(m1Inputs[78]), .ip2(n12921), .op(n12923) );
  or2_1 U12622 ( .ip1(n13803), .ip2(n12921), .op(n12922) );
  nand2_1 U12623 ( .ip1(n12923), .ip2(n12922), .op(n13060) );
  nand2_1 U12624 ( .ip1(m1Inputs[64]), .ip2(n14816), .op(n13062) );
  nor2_1 U12625 ( .ip1(n13060), .ip2(n13062), .op(n12924) );
  nor2_1 U12626 ( .ip1(n13061), .ip2(n12924), .op(n12977) );
  nor2_1 U12627 ( .ip1(n13766), .ip2(n12925), .op(n13000) );
  and2_1 U12628 ( .ip1(n13000), .ip2(n12926), .op(n12969) );
  nor2_1 U12629 ( .ip1(n13766), .ip2(n12999), .op(n12927) );
  or2_1 U12630 ( .ip1(m1Inputs[68]), .ip2(n12927), .op(n12929) );
  or2_1 U12631 ( .ip1(n14876), .ip2(n12927), .op(n12928) );
  nand2_1 U12632 ( .ip1(n12929), .ip2(n12928), .op(n12968) );
  nand2_1 U12633 ( .ip1(m1Inputs[66]), .ip2(\STAGE_1/weightReg [12]), .op(
        n12970) );
  nor2_1 U12634 ( .ip1(n12968), .ip2(n12970), .op(n12930) );
  nor2_1 U12635 ( .ip1(n12969), .ip2(n12930), .op(n12976) );
  xor2_1 U12636 ( .ip1(n12932), .ip2(n12931), .op(n12975) );
  fulladder U12637 ( .a(n12935), .b(n12934), .ci(n12933), .co(n13255), .s(
        n13260) );
  fulladder U12638 ( .a(n12938), .b(n12937), .ci(n12936), .co(n12855), .s(
        n12939) );
  inv_1 U12639 ( .ip(n12939), .op(n13015) );
  fulladder U12640 ( .a(n12942), .b(n12941), .ci(n12940), .co(n12933), .s(
        n13014) );
  fulladder U12641 ( .a(n12945), .b(n12944), .ci(n12943), .co(n12936), .s(
        n12946) );
  inv_1 U12642 ( .ip(n12946), .op(n13021) );
  fulladder U12643 ( .a(n12949), .b(n12948), .ci(n12947), .co(n12942), .s(
        n13020) );
  fulladder U12644 ( .a(n12952), .b(n12951), .ci(n12950), .co(n12947), .s(
        n13100) );
  nor2_1 U12645 ( .ip1(n12954), .ip2(n12953), .op(n12956) );
  xor2_1 U12646 ( .ip1(n12956), .ip2(n12955), .op(n13112) );
  nor2_1 U12647 ( .ip1(n12958), .ip2(n12957), .op(n12965) );
  nor2_1 U12648 ( .ip1(n13801), .ip2(n12959), .op(n12960) );
  or2_1 U12649 ( .ip1(m1Inputs[77]), .ip2(n12960), .op(n12962) );
  or2_1 U12650 ( .ip1(n13803), .ip2(n12960), .op(n12961) );
  nand2_1 U12651 ( .ip1(n12962), .ip2(n12961), .op(n12963) );
  nor2_1 U12652 ( .ip1(n12965), .ip2(n12963), .op(n13119) );
  or2_1 U12653 ( .ip1(n13119), .ip2(n12965), .op(n12967) );
  nor2_1 U12654 ( .ip1(n12964), .ip2(n14340), .op(n13118) );
  or2_1 U12655 ( .ip1(n13118), .ip2(n12965), .op(n12966) );
  nand2_1 U12656 ( .ip1(n12967), .ip2(n12966), .op(n13111) );
  nor2_1 U12657 ( .ip1(n12969), .ip2(n12968), .op(n12971) );
  xor2_1 U12658 ( .ip1(n12971), .ip2(n12970), .op(n13110) );
  fulladder U12659 ( .a(n12974), .b(n12973), .ci(n12972), .co(n13023), .s(
        n13107) );
  fulladder U12660 ( .a(n12977), .b(n12976), .ci(n12975), .co(n13022), .s(
        n13106) );
  fulladder U12661 ( .a(n12980), .b(n12979), .ci(n12978), .co(n12950), .s(
        n13104) );
  nand2_1 U12662 ( .ip1(m1Inputs[70]), .ip2(n4627), .op(n12983) );
  nand2_1 U12663 ( .ip1(m1Inputs[70]), .ip2(n12981), .op(n13047) );
  nor3_1 U12664 ( .ip1(n12982), .ip2(n14368), .ip3(n13047), .op(n12987) );
  or2_1 U12665 ( .ip1(n12983), .ip2(n12987), .op(n12986) );
  or2_1 U12666 ( .ip1(n12984), .ip2(n12987), .op(n12985) );
  nand2_1 U12667 ( .ip1(n12986), .ip2(n12985), .op(n13123) );
  or2_1 U12668 ( .ip1(n13123), .ip2(n12987), .op(n12989) );
  nor2_1 U12669 ( .ip1(n13050), .ip2(n14824), .op(n13122) );
  or2_1 U12670 ( .ip1(n13122), .ip2(n12987), .op(n12988) );
  nand2_1 U12671 ( .ip1(n12989), .ip2(n12988), .op(n13069) );
  nand2_1 U12672 ( .ip1(m1Inputs[72]), .ip2(\STAGE_1/weightReg [5]), .op(
        n12990) );
  nand2_1 U12673 ( .ip1(m1Inputs[72]), .ip2(\STAGE_1/weightReg [4]), .op(
        n13073) );
  nor3_1 U12674 ( .ip1(n13081), .ip2(n13835), .ip3(n13073), .op(n12994) );
  or2_1 U12675 ( .ip1(n12990), .ip2(n12994), .op(n12993) );
  or2_1 U12676 ( .ip1(n12991), .ip2(n12994), .op(n12992) );
  nand2_1 U12677 ( .ip1(n12993), .ip2(n12992), .op(n13121) );
  or2_1 U12678 ( .ip1(n13121), .ip2(n12994), .op(n12996) );
  nor2_1 U12679 ( .ip1(n13076), .ip2(n14188), .op(n13120) );
  or2_1 U12680 ( .ip1(n13120), .ip2(n12994), .op(n12995) );
  nand2_1 U12681 ( .ip1(n12996), .ip2(n12995), .op(n13068) );
  xor2_1 U12682 ( .ip1(n12998), .ip2(n12997), .op(n13067) );
  nand2_1 U12683 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[68]), .op(
        n13194) );
  nor3_1 U12684 ( .ip1(n13766), .ip2(n12999), .ip3(n13194), .op(n13088) );
  or2_1 U12685 ( .ip1(m1Inputs[69]), .ip2(n13000), .op(n13002) );
  or2_1 U12686 ( .ip1(n14838), .ip2(n13000), .op(n13001) );
  nand2_1 U12687 ( .ip1(n13002), .ip2(n13001), .op(n13087) );
  nand2_1 U12688 ( .ip1(m1Inputs[67]), .ip2(\STAGE_1/weightReg [10]), .op(
        n13089) );
  nor2_1 U12689 ( .ip1(n13087), .ip2(n13089), .op(n13003) );
  nor2_1 U12690 ( .ip1(n13088), .ip2(n13003), .op(n13066) );
  nand2_1 U12691 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[75]), .op(
        n13005) );
  nand2_1 U12692 ( .ip1(n13707), .ip2(m1Inputs[75]), .op(n13036) );
  nor3_1 U12693 ( .ip1(n13854), .ip2(n13004), .ip3(n13036), .op(n13009) );
  or2_1 U12694 ( .ip1(n13005), .ip2(n13009), .op(n13008) );
  or2_1 U12695 ( .ip1(n13006), .ip2(n13009), .op(n13007) );
  nand2_1 U12696 ( .ip1(n13008), .ip2(n13007), .op(n13055) );
  or2_1 U12697 ( .ip1(n13055), .ip2(n13009), .op(n13012) );
  nand2_1 U12698 ( .ip1(column[69]), .ip2(n15042), .op(n13054) );
  inv_1 U12699 ( .ip(n13054), .op(n13010) );
  or2_1 U12700 ( .ip1(n13010), .ip2(n13009), .op(n13011) );
  nand2_1 U12701 ( .ip1(n13012), .ip2(n13011), .op(n13065) );
  nand2_1 U12702 ( .ip1(m1Inputs[67]), .ip2(n13718), .op(n13064) );
  fulladder U12703 ( .a(n13015), .b(n13014), .ci(n13013), .co(n13259), .s(
        n13264) );
  fulladder U12704 ( .a(n13018), .b(n13017), .ci(n13016), .co(n12940), .s(
        n13093) );
  fulladder U12705 ( .a(n13021), .b(n13020), .ci(n13019), .co(n13013), .s(
        n13092) );
  fulladder U12706 ( .a(n13024), .b(n13023), .ci(n13022), .co(n13016), .s(
        n13096) );
  fulladder U12707 ( .a(n13027), .b(n13026), .ci(n13025), .co(n12903), .s(
        n13028) );
  inv_1 U12708 ( .ip(n13028), .op(n13095) );
  fulladder U12709 ( .a(n13031), .b(n13030), .ci(n13029), .co(n13027), .s(
        n13032) );
  inv_1 U12710 ( .ip(n13032), .op(n13131) );
  nand2_1 U12711 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[74]), .op(
        n13035) );
  nor3_1 U12712 ( .ip1(n13854), .ip2(n13034), .ip3(n13033), .op(n13040) );
  or2_1 U12713 ( .ip1(n13035), .ip2(n13040), .op(n13038) );
  or2_1 U12714 ( .ip1(n13036), .ip2(n13040), .op(n13037) );
  nand2_1 U12715 ( .ip1(n13038), .ip2(n13037), .op(n13166) );
  or2_1 U12716 ( .ip1(n13166), .ip2(n13040), .op(n13043) );
  nand2_1 U12717 ( .ip1(column[68]), .ip2(n13039), .op(n13165) );
  inv_1 U12718 ( .ip(n13165), .op(n13041) );
  or2_1 U12719 ( .ip1(n13041), .ip2(n13040), .op(n13042) );
  nand2_1 U12720 ( .ip1(n13043), .ip2(n13042), .op(n13148) );
  nand2_1 U12721 ( .ip1(n14835), .ip2(m1Inputs[69]), .op(n13046) );
  nor3_1 U12722 ( .ip1(n13045), .ip2(n14384), .ip3(n13044), .op(n13051) );
  or2_1 U12723 ( .ip1(n13046), .ip2(n13051), .op(n13049) );
  or2_1 U12724 ( .ip1(n13047), .ip2(n13051), .op(n13048) );
  nand2_1 U12725 ( .ip1(n13049), .ip2(n13048), .op(n13175) );
  or2_1 U12726 ( .ip1(n13175), .ip2(n13051), .op(n13053) );
  nor2_1 U12727 ( .ip1(n13050), .ip2(n13594), .op(n13174) );
  or2_1 U12728 ( .ip1(n13174), .ip2(n13051), .op(n13052) );
  nand2_1 U12729 ( .ip1(n13053), .ip2(n13052), .op(n13147) );
  xor2_1 U12730 ( .ip1(n13055), .ip2(n13054), .op(n13146) );
  nor2_1 U12731 ( .ip1(n13057), .ip2(n13056), .op(n13059) );
  xor2_1 U12732 ( .ip1(n13059), .ip2(n13058), .op(n13115) );
  nor2_1 U12733 ( .ip1(n13061), .ip2(n13060), .op(n13063) );
  xor2_1 U12734 ( .ip1(n13063), .ip2(n13062), .op(n13114) );
  fulladder U12735 ( .a(n13066), .b(n13065), .ci(n13064), .co(n13102), .s(
        n13138) );
  fulladder U12736 ( .a(n13069), .b(n13068), .ci(n13067), .co(n13103), .s(
        n13137) );
  nand2_1 U12737 ( .ip1(m1Inputs[71]), .ip2(\STAGE_1/weightReg [5]), .op(
        n13072) );
  nor3_1 U12738 ( .ip1(n13071), .ip2(n13835), .ip3(n13070), .op(n13077) );
  or2_1 U12739 ( .ip1(n13072), .ip2(n13077), .op(n13075) );
  or2_1 U12740 ( .ip1(n13073), .ip2(n13077), .op(n13074) );
  nand2_1 U12741 ( .ip1(n13075), .ip2(n13074), .op(n13173) );
  or2_1 U12742 ( .ip1(n13173), .ip2(n13077), .op(n13079) );
  nor2_1 U12743 ( .ip1(n13076), .ip2(n14824), .op(n13172) );
  or2_1 U12744 ( .ip1(n13172), .ip2(n13077), .op(n13078) );
  nand2_1 U12745 ( .ip1(n13079), .ip2(n13078), .op(n13141) );
  nor3_1 U12746 ( .ip1(n10476), .ip2(n13081), .ip3(n13080), .op(n13196) );
  nor2_1 U12747 ( .ip1(n13082), .ip2(n13081), .op(n13083) );
  or2_1 U12748 ( .ip1(m1Inputs[76]), .ip2(n13083), .op(n13085) );
  or2_1 U12749 ( .ip1(n13803), .ip2(n13083), .op(n13084) );
  nand2_1 U12750 ( .ip1(n13085), .ip2(n13084), .op(n13195) );
  nand2_1 U12751 ( .ip1(m1Inputs[64]), .ip2(\STAGE_1/weightReg [12]), .op(
        n13197) );
  nor2_1 U12752 ( .ip1(n13195), .ip2(n13197), .op(n13086) );
  nor2_1 U12753 ( .ip1(n13196), .ip2(n13086), .op(n13140) );
  nor2_1 U12754 ( .ip1(n13088), .ip2(n13087), .op(n13090) );
  xor2_1 U12755 ( .ip1(n13090), .ip2(n13089), .op(n13139) );
  fulladder U12756 ( .a(n13093), .b(n13092), .ci(n13091), .co(n13263), .s(
        n13268) );
  fulladder U12757 ( .a(n13096), .b(n13095), .ci(n13094), .co(n13091), .s(
        n13097) );
  inv_1 U12758 ( .ip(n13097), .op(n13127) );
  fulladder U12759 ( .a(n13100), .b(n13099), .ci(n13098), .co(n13019), .s(
        n13101) );
  inv_1 U12760 ( .ip(n13101), .op(n13126) );
  fulladder U12761 ( .a(n13104), .b(n13103), .ci(n13102), .co(n13098), .s(
        n13105) );
  inv_1 U12762 ( .ip(n13105), .op(n13134) );
  fulladder U12763 ( .a(n13108), .b(n13107), .ci(n13106), .co(n13099), .s(
        n13109) );
  inv_1 U12764 ( .ip(n13109), .op(n13133) );
  fulladder U12765 ( .a(n13112), .b(n13111), .ci(n13110), .co(n13108), .s(
        n13113) );
  inv_1 U12766 ( .ip(n13113), .op(n13181) );
  fulladder U12767 ( .a(n13116), .b(n13115), .ci(n13114), .co(n13130), .s(
        n13117) );
  inv_1 U12768 ( .ip(n13117), .op(n13180) );
  xor2_1 U12769 ( .ip1(n13119), .ip2(n13118), .op(n13144) );
  xor2_1 U12770 ( .ip1(n13121), .ip2(n13120), .op(n13143) );
  xor2_1 U12771 ( .ip1(n13123), .ip2(n13122), .op(n13142) );
  inv_1 U12772 ( .ip(n13124), .op(n13267) );
  fulladder U12773 ( .a(n13127), .b(n13126), .ci(n13125), .co(n13124), .s(
        n13128) );
  inv_1 U12774 ( .ip(n13128), .op(n13272) );
  fulladder U12775 ( .a(n13131), .b(n13130), .ci(n13129), .co(n13094), .s(
        n13178) );
  fulladder U12776 ( .a(n13134), .b(n13133), .ci(n13132), .co(n13125), .s(
        n13135) );
  inv_1 U12777 ( .ip(n13135), .op(n13177) );
  fulladder U12778 ( .a(n13138), .b(n13137), .ci(n13136), .co(n13129), .s(
        n13185) );
  fulladder U12779 ( .a(n13141), .b(n13140), .ci(n13139), .co(n13136), .s(
        n13214) );
  fulladder U12780 ( .a(n13144), .b(n13143), .ci(n13142), .co(n13179), .s(
        n13145) );
  inv_1 U12781 ( .ip(n13145), .op(n13213) );
  fulladder U12782 ( .a(n13148), .b(n13147), .ci(n13146), .co(n13116), .s(
        n13212) );
  or2_1 U12783 ( .ip1(n13149), .ip2(n13151), .op(n13154) );
  inv_1 U12784 ( .ip(n13150), .op(n13152) );
  or2_1 U12785 ( .ip1(n13152), .ip2(n13151), .op(n13153) );
  nand2_1 U12786 ( .ip1(n13154), .ip2(n13153), .op(n13193) );
  nand2_1 U12787 ( .ip1(m1Inputs[67]), .ip2(n14994), .op(n13192) );
  or2_1 U12788 ( .ip1(n13155), .ip2(n13156), .op(n13159) );
  or2_1 U12789 ( .ip1(n13157), .ip2(n13156), .op(n13158) );
  nand2_1 U12790 ( .ip1(n13159), .ip2(n13158), .op(n13201) );
  or2_1 U12791 ( .ip1(n13160), .ip2(n13161), .op(n13164) );
  or2_1 U12792 ( .ip1(n13162), .ip2(n13161), .op(n13163) );
  nand2_1 U12793 ( .ip1(n13164), .ip2(n13163), .op(n13200) );
  xor2_1 U12794 ( .ip1(n13166), .ip2(n13165), .op(n13199) );
  or2_1 U12795 ( .ip1(n13167), .ip2(n13168), .op(n13171) );
  or2_1 U12796 ( .ip1(n13169), .ip2(n13168), .op(n13170) );
  nand2_1 U12797 ( .ip1(n13171), .ip2(n13170), .op(n13220) );
  xnor2_1 U12798 ( .ip1(n13173), .ip2(n13172), .op(n13219) );
  xnor2_1 U12799 ( .ip1(n13175), .ip2(n13174), .op(n13218) );
  fulladder U12800 ( .a(n13178), .b(n13177), .ci(n13176), .co(n13271), .s(
        n13276) );
  fulladder U12801 ( .a(n13181), .b(n13180), .ci(n13179), .co(n13132), .s(
        n13182) );
  inv_1 U12802 ( .ip(n13182), .op(n13211) );
  fulladder U12803 ( .a(n13185), .b(n13184), .ci(n13183), .co(n13176), .s(
        n13210) );
  fulladder U12804 ( .a(n13188), .b(n13187), .ci(n13186), .co(n13183), .s(
        n13217) );
  fulladder U12805 ( .a(n13191), .b(n13190), .ci(n13189), .co(n13223), .s(
        n13226) );
  fulladder U12806 ( .a(n13194), .b(n13193), .ci(n13192), .co(n13188), .s(
        n13222) );
  nor2_1 U12807 ( .ip1(n13196), .ip2(n13195), .op(n13198) );
  xor2_1 U12808 ( .ip1(n13198), .ip2(n13197), .op(n13221) );
  fulladder U12809 ( .a(n13201), .b(n13200), .ci(n13199), .co(n13187), .s(
        n13232) );
  fulladder U12810 ( .a(n13204), .b(n13203), .ci(n13202), .co(n13205), .s(
        n12582) );
  inv_1 U12811 ( .ip(n13205), .op(n13231) );
  fulladder U12812 ( .a(n13208), .b(n13207), .ci(n13206), .co(n13230), .s(
        n13238) );
  fulladder U12813 ( .a(n13211), .b(n13210), .ci(n13209), .co(n13275), .s(
        n13280) );
  fulladder U12814 ( .a(n13214), .b(n13213), .ci(n13212), .co(n13184), .s(
        n13229) );
  fulladder U12815 ( .a(n13217), .b(n13216), .ci(n13215), .co(n13209), .s(
        n13228) );
  fulladder U12816 ( .a(n13220), .b(n13219), .ci(n13218), .co(n13186), .s(
        n13235) );
  fulladder U12817 ( .a(n13223), .b(n13222), .ci(n13221), .co(n13216), .s(
        n13234) );
  fulladder U12818 ( .a(n13226), .b(n13225), .ci(n13224), .co(n13233), .s(
        n13248) );
  fulladder U12819 ( .a(n13229), .b(n13228), .ci(n13227), .co(n13279), .s(
        n13284) );
  fulladder U12820 ( .a(n13232), .b(n13231), .ci(n13230), .co(n13215), .s(
        n13241) );
  fulladder U12821 ( .a(n13235), .b(n13234), .ci(n13233), .co(n13227), .s(
        n13240) );
  fulladder U12822 ( .a(n13238), .b(n13237), .ci(n13236), .co(n13239), .s(
        n13247) );
  fulladder U12823 ( .a(n13241), .b(n13240), .ci(n13239), .co(n13283), .s(
        n13288) );
  fulladder U12824 ( .a(n13244), .b(n13243), .ci(n13242), .co(n13245), .s(
        \STAGE_1/M5/sum [3]) );
  inv_1 U12825 ( .ip(n13245), .op(n13287) );
  fulladder U12826 ( .a(n13248), .b(n13247), .ci(n13246), .co(n13286), .s(
        n12589) );
  inv_1 U12827 ( .ip(n13249), .op(\STAGE_1/M5/sum [14]) );
  fulladder U12828 ( .a(n13252), .b(n13251), .ci(n13250), .co(n13312), .s(
        n13253) );
  inv_1 U12829 ( .ip(n13253), .op(\STAGE_1/M5/sum [13]) );
  fulladder U12830 ( .a(n13256), .b(n13255), .ci(n13254), .co(n13250), .s(
        n13257) );
  inv_1 U12831 ( .ip(n13257), .op(\STAGE_1/M5/sum [12]) );
  fulladder U12832 ( .a(n13260), .b(n13259), .ci(n13258), .co(n13254), .s(
        n13261) );
  inv_1 U12833 ( .ip(n13261), .op(\STAGE_1/M5/sum [11]) );
  fulladder U12834 ( .a(n13264), .b(n13263), .ci(n13262), .co(n13258), .s(
        n13265) );
  inv_1 U12835 ( .ip(n13265), .op(\STAGE_1/M5/sum [10]) );
  fulladder U12836 ( .a(n13268), .b(n13267), .ci(n13266), .co(n13262), .s(
        n13269) );
  inv_1 U12837 ( .ip(n13269), .op(\STAGE_1/M5/sum [9]) );
  fulladder U12838 ( .a(n13272), .b(n13271), .ci(n13270), .co(n13266), .s(
        n13273) );
  inv_1 U12839 ( .ip(n13273), .op(\STAGE_1/M5/sum [8]) );
  fulladder U12840 ( .a(n13276), .b(n13275), .ci(n13274), .co(n13270), .s(
        n13277) );
  inv_1 U12841 ( .ip(n13277), .op(\STAGE_1/M5/sum [7]) );
  fulladder U12842 ( .a(n13280), .b(n13279), .ci(n13278), .co(n13274), .s(
        n13281) );
  inv_1 U12843 ( .ip(n13281), .op(\STAGE_1/M5/sum [6]) );
  fulladder U12844 ( .a(n13284), .b(n13283), .ci(n13282), .co(n13278), .s(
        n13285) );
  inv_1 U12845 ( .ip(n13285), .op(\STAGE_1/M5/sum [5]) );
  fulladder U12846 ( .a(n13288), .b(n13287), .ci(n13286), .co(n13282), .s(
        n13289) );
  inv_1 U12847 ( .ip(n13289), .op(\STAGE_1/M5/sum [4]) );
  nand2_1 U12848 ( .ip1(m1Inputs[72]), .ip2(n14976), .op(n13291) );
  nand2_1 U12849 ( .ip1(m1Inputs[73]), .ip2(\STAGE_1/weightReg [14]), .op(
        n13290) );
  xor2_1 U12850 ( .ip1(n13291), .ip2(n13290), .op(n13296) );
  fulladder U12851 ( .a(n13294), .b(n13293), .ci(n13292), .co(n13295), .s(
        n13314) );
  xor2_1 U12852 ( .ip1(n13296), .ip2(n13295), .op(n13306) );
  fulladder U12853 ( .a(n13299), .b(n13298), .ci(n13297), .co(n13304), .s(
        n12676) );
  fulladder U12854 ( .a(n13302), .b(n13301), .ci(n13300), .co(n13303), .s(
        n12646) );
  xor2_1 U12855 ( .ip1(n13304), .ip2(n13303), .op(n13305) );
  xor2_1 U12856 ( .ip1(n13306), .ip2(n13305), .op(n13308) );
  nand2_1 U12857 ( .ip1(m1Inputs[79]), .ip2(n14975), .op(n13307) );
  xor2_1 U12858 ( .ip1(n13308), .ip2(n13307), .op(n13350) );
  fulladder U12859 ( .a(n13311), .b(n13310), .ci(n13309), .co(n13316), .s(
        n13298) );
  fulladder U12860 ( .a(n13314), .b(n13313), .ci(n13312), .co(n13315), .s(
        n13249) );
  xor2_1 U12861 ( .ip1(n13316), .ip2(n13315), .op(n13317) );
  xor2_1 U12862 ( .ip1(n13318), .ip2(n13317), .op(n13346) );
  fulladder U12863 ( .a(n13321), .b(n13320), .ci(n13319), .co(n13326), .s(
        n12642) );
  fulladder U12864 ( .a(n13324), .b(n13323), .ci(n13322), .co(n13325), .s(
        n13328) );
  xor2_1 U12865 ( .ip1(n13326), .ip2(n13325), .op(n13336) );
  fulladder U12866 ( .a(n13329), .b(n13328), .ci(n13327), .co(n13334), .s(
        n12634) );
  fulladder U12867 ( .a(n13332), .b(n13331), .ci(n13330), .co(n13333), .s(
        n13310) );
  xor2_1 U12868 ( .ip1(n13334), .ip2(n13333), .op(n13335) );
  xor2_1 U12869 ( .ip1(n13336), .ip2(n13335), .op(n13344) );
  nand2_1 U12870 ( .ip1(m1Inputs[78]), .ip2(n14994), .op(n13338) );
  nand2_1 U12871 ( .ip1(m1Inputs[77]), .ip2(\STAGE_1/weightReg [10]), .op(
        n13337) );
  xor2_1 U12872 ( .ip1(n13338), .ip2(n13337), .op(n13342) );
  nand2_1 U12873 ( .ip1(m1Inputs[74]), .ip2(\STAGE_1/weightReg [13]), .op(
        n13340) );
  nand2_1 U12874 ( .ip1(m1Inputs[75]), .ip2(\STAGE_1/weightReg [12]), .op(
        n13339) );
  xor2_1 U12875 ( .ip1(n13340), .ip2(n13339), .op(n13341) );
  xor2_1 U12876 ( .ip1(n13342), .ip2(n13341), .op(n13343) );
  xor2_1 U12877 ( .ip1(n13344), .ip2(n13343), .op(n13345) );
  xor2_1 U12878 ( .ip1(n13346), .ip2(n13345), .op(n13348) );
  nand2_1 U12879 ( .ip1(n15042), .ip2(column[79]), .op(n13347) );
  xor2_1 U12880 ( .ip1(n13348), .ip2(n13347), .op(n13349) );
  xor2_1 U12881 ( .ip1(n13350), .ip2(n13349), .op(n13355) );
  nand3_1 U12882 ( .ip1(column[78]), .ip2(n15042), .ip3(n13351), .op(n13352)
         );
  nand2_1 U12883 ( .ip1(n13353), .ip2(n13352), .op(n13354) );
  xor2_1 U12884 ( .ip1(n13355), .ip2(n13354), .op(\STAGE_1/M5/sum [15]) );
  or2_1 U12885 ( .ip1(n13356), .ip2(n13357), .op(n13360) );
  or2_1 U12886 ( .ip1(n13358), .ip2(n13357), .op(n13359) );
  nand2_1 U12887 ( .ip1(n13360), .ip2(n13359), .op(n13987) );
  or2_1 U12888 ( .ip1(n13361), .ip2(n13362), .op(n13365) );
  or2_1 U12889 ( .ip1(n13363), .ip2(n13362), .op(n13364) );
  nand2_1 U12890 ( .ip1(n13365), .ip2(n13364), .op(n13986) );
  nand2_1 U12891 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[90]), .op(
        n13367) );
  inv_1 U12892 ( .ip(m1Inputs[91]), .op(n13760) );
  nor3_1 U12893 ( .ip1(n13854), .ip2(n13760), .ip3(n13366), .op(n13886) );
  or2_1 U12894 ( .ip1(n13367), .ip2(n13886), .op(n13369) );
  nand2_1 U12895 ( .ip1(n13707), .ip2(m1Inputs[91]), .op(n13852) );
  or2_1 U12896 ( .ip1(n13852), .ip2(n13886), .op(n13368) );
  nand2_1 U12897 ( .ip1(n13369), .ip2(n13368), .op(n13884) );
  nand2_1 U12898 ( .ip1(column[84]), .ip2(n13859), .op(n13885) );
  xor2_1 U12899 ( .ip1(n13884), .ip2(n13885), .op(n13985) );
  fulladder U12900 ( .a(n13372), .b(n13371), .ci(n13370), .co(n13373), .s(
        n6451) );
  inv_1 U12901 ( .ip(n13373), .op(n14008) );
  fulladder U12902 ( .a(n13376), .b(n13375), .ci(n13374), .co(n14007), .s(
        n13409) );
  or2_1 U12903 ( .ip1(n13377), .ip2(n13378), .op(n13381) );
  or2_1 U12904 ( .ip1(n13379), .ip2(n13378), .op(n13380) );
  nand2_1 U12905 ( .ip1(n13381), .ip2(n13380), .op(n13990) );
  nand2_1 U12906 ( .ip1(m1Inputs[87]), .ip2(\STAGE_1/weightReg [5]), .op(
        n13383) );
  nor3_1 U12907 ( .ip1(n13748), .ip2(n13835), .ip3(n13382), .op(n13912) );
  or2_1 U12908 ( .ip1(n13383), .ip2(n13912), .op(n13385) );
  nand2_1 U12909 ( .ip1(m1Inputs[88]), .ip2(n13637), .op(n13834) );
  or2_1 U12910 ( .ip1(n13834), .ip2(n13912), .op(n13384) );
  nand2_1 U12911 ( .ip1(n13385), .ip2(n13384), .op(n13911) );
  nor2_1 U12912 ( .ip1(n13841), .ip2(n13579), .op(n13913) );
  xnor2_1 U12913 ( .ip1(n13911), .ip2(n13913), .op(n13989) );
  nand2_1 U12914 ( .ip1(n14835), .ip2(m1Inputs[85]), .op(n13387) );
  nor3_1 U12915 ( .ip1(n13578), .ip2(n14368), .ip3(n13386), .op(n13891) );
  or2_1 U12916 ( .ip1(n13387), .ip2(n13891), .op(n13389) );
  nand2_1 U12917 ( .ip1(m1Inputs[86]), .ip2(n12981), .op(n13824) );
  or2_1 U12918 ( .ip1(n13824), .ip2(n13891), .op(n13388) );
  nand2_1 U12919 ( .ip1(n13389), .ip2(n13388), .op(n13890) );
  nor2_1 U12920 ( .ip1(n13830), .ip2(n13390), .op(n13892) );
  xnor2_1 U12921 ( .ip1(n13890), .ip2(n13892), .op(n13988) );
  fulladder U12922 ( .a(n13393), .b(n13392), .ci(n13391), .co(n14006), .s(
        n13406) );
  nand2_1 U12923 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[84]), .op(
        n13984) );
  or2_1 U12924 ( .ip1(n13394), .ip2(n13396), .op(n13399) );
  inv_1 U12925 ( .ip(n13395), .op(n13397) );
  or2_1 U12926 ( .ip1(n13397), .ip2(n13396), .op(n13398) );
  nand2_1 U12927 ( .ip1(n13399), .ip2(n13398), .op(n13983) );
  nand2_1 U12928 ( .ip1(m1Inputs[83]), .ip2(n14994), .op(n13982) );
  nand2_1 U12929 ( .ip1(n13614), .ip2(m1Inputs[92]), .op(n13729) );
  nor3_1 U12930 ( .ip1(n13646), .ip2(n13836), .ip3(n13729), .op(n13919) );
  nor2_1 U12931 ( .ip1(n13801), .ip2(n13836), .op(n13400) );
  or2_1 U12932 ( .ip1(m1Inputs[92]), .ip2(n13400), .op(n13402) );
  or2_1 U12933 ( .ip1(n13803), .ip2(n13400), .op(n13401) );
  nand2_1 U12934 ( .ip1(n13402), .ip2(n13401), .op(n13917) );
  nor2_1 U12935 ( .ip1(n13919), .ip2(n13917), .op(n13403) );
  nand2_1 U12936 ( .ip1(m1Inputs[80]), .ip2(\STAGE_1/weightReg [12]), .op(
        n13916) );
  xor2_1 U12937 ( .ip1(n13403), .ip2(n13916), .op(n14004) );
  fulladder U12938 ( .a(n13406), .b(n13405), .ci(n13404), .co(n14019), .s(
        n13413) );
  fulladder U12939 ( .a(n13409), .b(n13408), .ci(n13407), .co(n14029), .s(
        n13412) );
  inv_1 U12940 ( .ip(n13410), .op(n14027) );
  fulladder U12941 ( .a(n13413), .b(n13412), .ci(n13411), .co(n13414), .s(
        n6469) );
  inv_1 U12942 ( .ip(n13414), .op(n14026) );
  fulladder U12943 ( .a(n13417), .b(n13416), .ci(n13415), .co(n14025), .s(
        \STAGE_1/M6/sum [3]) );
  inv_1 U12944 ( .ip(m1Inputs[92]), .op(n13853) );
  nor2_1 U12945 ( .ip1(n13766), .ip2(n13853), .op(n13508) );
  inv_1 U12946 ( .ip(m1Inputs[94]), .op(n13675) );
  nor2_1 U12947 ( .ip1(n13675), .ip2(n14384), .op(n13507) );
  nand2_1 U12948 ( .ip1(n14976), .ip2(m1Inputs[86]), .op(n13506) );
  inv_1 U12949 ( .ip(n13418), .op(n13512) );
  nor2_1 U12950 ( .ip1(n14188), .ip2(n13836), .op(n13492) );
  inv_1 U12951 ( .ip(m1Inputs[93]), .op(n13708) );
  nor2_1 U12952 ( .ip1(n6503), .ip2(n13708), .op(n13491) );
  nand2_1 U12953 ( .ip1(m1Inputs[95]), .ip2(n12981), .op(n13490) );
  inv_1 U12954 ( .ip(n13419), .op(n13511) );
  inv_1 U12955 ( .ip(m1Inputs[95]), .op(n13645) );
  nor2_1 U12956 ( .ip1(n13645), .ip2(n8942), .op(n13433) );
  nand2_1 U12957 ( .ip1(m1Inputs[94]), .ip2(n12981), .op(n13432) );
  nand2_1 U12958 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[92]), .op(
        n13431) );
  nand2_1 U12959 ( .ip1(m1Inputs[87]), .ip2(\STAGE_1/weightReg [13]), .op(
        n13421) );
  nand2_1 U12960 ( .ip1(m1Inputs[89]), .ip2(n14847), .op(n13420) );
  xor2_1 U12961 ( .ip1(n13421), .ip2(n13420), .op(n13461) );
  nor2_1 U12962 ( .ip1(n13579), .ip2(n13825), .op(n13464) );
  nor2_1 U12963 ( .ip1(n14340), .ip2(n13836), .op(n14111) );
  and2_1 U12964 ( .ip1(n13464), .ip2(n14111), .op(n13422) );
  or2_1 U12965 ( .ip1(n13461), .ip2(n13422), .op(n13424) );
  nor2_1 U12966 ( .ip1(n14842), .ip2(n13578), .op(n13460) );
  or2_1 U12967 ( .ip1(n13460), .ip2(n13422), .op(n13423) );
  nand2_1 U12968 ( .ip1(n13424), .ip2(n13423), .op(n13519) );
  nand2_1 U12969 ( .ip1(n14629), .ip2(m1Inputs[91]), .op(n13444) );
  nand2_1 U12970 ( .ip1(n13718), .ip2(m1Inputs[91]), .op(n13493) );
  nand2_1 U12971 ( .ip1(n14629), .ip2(m1Inputs[90]), .op(n13445) );
  nor2_1 U12972 ( .ip1(n13493), .ip2(n13445), .op(n13502) );
  or2_1 U12973 ( .ip1(n13444), .ip2(n13502), .op(n13427) );
  nand2_1 U12974 ( .ip1(n13718), .ip2(m1Inputs[90]), .op(n13425) );
  or2_1 U12975 ( .ip1(n13425), .ip2(n13502), .op(n13426) );
  nand2_1 U12976 ( .ip1(n13427), .ip2(n13426), .op(n13503) );
  nand2_1 U12977 ( .ip1(column[93]), .ip2(n13859), .op(n13428) );
  xor2_1 U12978 ( .ip1(n13503), .ip2(n13428), .op(n13518) );
  nor2_1 U12979 ( .ip1(n14853), .ip2(n13847), .op(n13430) );
  nand2_1 U12980 ( .ip1(n15025), .ip2(m1Inputs[88]), .op(n13465) );
  nand2_1 U12981 ( .ip1(m1Inputs[93]), .ip2(n4627), .op(n13429) );
  fulladder U12982 ( .a(n13430), .b(n13465), .ci(n13429), .co(n13517), .s(
        n13532) );
  fulladder U12983 ( .a(n13433), .b(n13432), .ci(n13431), .co(n13510), .s(
        n13531) );
  nand2_1 U12984 ( .ip1(n13718), .ip2(m1Inputs[92]), .op(n14097) );
  nand2_1 U12985 ( .ip1(m1Inputs[87]), .ip2(n12981), .op(n13827) );
  nor2_1 U12986 ( .ip1(n14097), .ip2(n13827), .op(n13606) );
  or2_1 U12987 ( .ip1(n13749), .ip2(n13464), .op(n13435) );
  or2_1 U12988 ( .ip1(m1Inputs[92]), .ip2(n13464), .op(n13434) );
  nand2_1 U12989 ( .ip1(n13435), .ip2(n13434), .op(n13605) );
  nand2_1 U12990 ( .ip1(n14816), .ip2(m1Inputs[84]), .op(n13607) );
  nor2_1 U12991 ( .ip1(n13605), .ip2(n13607), .op(n13436) );
  nor2_1 U12992 ( .ip1(n13606), .ip2(n13436), .op(n13540) );
  nand2_1 U12993 ( .ip1(m1Inputs[90]), .ip2(n14975), .op(n13438) );
  nand2_1 U12994 ( .ip1(m1Inputs[88]), .ip2(\STAGE_1/weightReg [10]), .op(
        n13437) );
  xor2_1 U12995 ( .ip1(n13438), .ip2(n13437), .op(n13550) );
  nor2_1 U12996 ( .ip1(n6503), .ip2(n13748), .op(n13704) );
  and3_1 U12997 ( .ip1(n14629), .ip2(m1Inputs[90]), .ip3(n13704), .op(n13439)
         );
  or2_1 U12998 ( .ip1(n13550), .ip2(n13439), .op(n13442) );
  nand2_1 U12999 ( .ip1(column[90]), .ip2(n13859), .op(n13549) );
  inv_1 U13000 ( .ip(n13549), .op(n13440) );
  or2_1 U13001 ( .ip1(n13440), .ip2(n13439), .op(n13441) );
  nand2_1 U13002 ( .ip1(n13442), .ip2(n13441), .op(n13539) );
  nand2_1 U13003 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[86]), .op(
        n13538) );
  inv_1 U13004 ( .ip(n13443), .op(n13528) );
  nand2_1 U13005 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[88]), .op(
        n13515) );
  nand2_1 U13006 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[90]), .op(
        n13450) );
  nor2_1 U13007 ( .ip1(n13444), .ip2(n13450), .op(n13457) );
  inv_1 U13008 ( .ip(n13445), .op(n13449) );
  or2_1 U13009 ( .ip1(m1Inputs[91]), .ip2(n13449), .op(n13447) );
  or2_1 U13010 ( .ip1(\STAGE_1/weightReg [9]), .ip2(n13449), .op(n13446) );
  nand2_1 U13011 ( .ip1(n13447), .ip2(n13446), .op(n13456) );
  nand2_1 U13012 ( .ip1(column[92]), .ip2(n13859), .op(n13458) );
  nor2_1 U13013 ( .ip1(n13456), .ip2(n13458), .op(n13448) );
  nor2_1 U13014 ( .ip1(n13457), .ip2(n13448), .op(n13514) );
  nand2_1 U13015 ( .ip1(n14816), .ip2(m1Inputs[87]), .op(n13513) );
  nor2_1 U13016 ( .ip1(n12083), .ip2(n13836), .op(n13589) );
  nand2_1 U13017 ( .ip1(n13449), .ip2(n13589), .op(n13452) );
  inv_1 U13018 ( .ip(n13452), .op(n13455) );
  nand2_1 U13019 ( .ip1(m1Inputs[89]), .ip2(n14629), .op(n13451) );
  nand2_1 U13020 ( .ip1(n13451), .ip2(n13450), .op(n13453) );
  nand2_1 U13021 ( .ip1(n13453), .ip2(n13452), .op(n13486) );
  nand2_1 U13022 ( .ip1(column[91]), .ip2(n13859), .op(n13485) );
  nor2_1 U13023 ( .ip1(n13486), .ip2(n13485), .op(n13454) );
  nor2_1 U13024 ( .ip1(n13455), .ip2(n13454), .op(n13473) );
  nand2_1 U13025 ( .ip1(m1Inputs[93]), .ip2(\STAGE_1/weightReg [6]), .op(
        n13483) );
  nor2_1 U13026 ( .ip1(n14853), .ip2(n13765), .op(n13482) );
  nand2_1 U13027 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[91]), .op(
        n13481) );
  nor2_1 U13028 ( .ip1(n13457), .ip2(n13456), .op(n13459) );
  xor2_1 U13029 ( .ip1(n13459), .ip2(n13458), .op(n13471) );
  xnor2_1 U13030 ( .ip1(n13461), .ip2(n13460), .op(n13536) );
  nand2_1 U13031 ( .ip1(m1Inputs[87]), .ip2(\STAGE_1/weightReg [12]), .op(
        n13463) );
  nand2_1 U13032 ( .ip1(m1Inputs[88]), .ip2(n13718), .op(n13462) );
  xor2_1 U13033 ( .ip1(n13463), .ip2(n13462), .op(n13476) );
  inv_1 U13034 ( .ip(n13464), .op(n13466) );
  nor2_1 U13035 ( .ip1(n13466), .ip2(n13465), .op(n13467) );
  or2_1 U13036 ( .ip1(n13476), .ip2(n13467), .op(n13469) );
  nor2_1 U13037 ( .ip1(n14842), .ip2(n13847), .op(n13475) );
  or2_1 U13038 ( .ip1(n13475), .ip2(n13467), .op(n13468) );
  nand2_1 U13039 ( .ip1(n13469), .ip2(n13468), .op(n13535) );
  nor2_1 U13040 ( .ip1(n13645), .ip2(n14783), .op(n13479) );
  nand2_1 U13041 ( .ip1(m1Inputs[92]), .ip2(n4627), .op(n13478) );
  nand2_1 U13042 ( .ip1(m1Inputs[94]), .ip2(\STAGE_1/weightReg [5]), .op(
        n13477) );
  inv_1 U13043 ( .ip(n13470), .op(n13527) );
  fulladder U13044 ( .a(n13473), .b(n13472), .ci(n13471), .co(n13521), .s(
        n13474) );
  inv_1 U13045 ( .ip(n13474), .op(n13555) );
  xor2_1 U13046 ( .ip1(n13476), .ip2(n13475), .op(n13603) );
  fulladder U13047 ( .a(n13479), .b(n13478), .ci(n13477), .co(n13534), .s(
        n13480) );
  inv_1 U13048 ( .ip(n13480), .op(n13602) );
  fulladder U13049 ( .a(n13483), .b(n13482), .ci(n13481), .co(n13472), .s(
        n13484) );
  inv_1 U13050 ( .ip(n13484), .op(n13601) );
  xor2_1 U13051 ( .ip1(n13486), .ip2(n13485), .op(n13599) );
  nand2_1 U13052 ( .ip1(m1Inputs[94]), .ip2(n13637), .op(n13586) );
  nor2_1 U13053 ( .ip1(n13487), .ip2(n13645), .op(n13585) );
  nand2_1 U13054 ( .ip1(m1Inputs[91]), .ip2(n4627), .op(n13584) );
  inv_1 U13055 ( .ip(n13488), .op(n13598) );
  nor2_1 U13056 ( .ip1(n13708), .ip2(n8942), .op(n13590) );
  nand2_1 U13057 ( .ip1(m1Inputs[83]), .ip2(n14976), .op(n13588) );
  inv_1 U13058 ( .ip(n13489), .op(n14078) );
  fulladder U13059 ( .a(n13492), .b(n13491), .ci(n13490), .co(n14081), .s(
        n13419) );
  nand4_1 U13060 ( .ip1(\STAGE_1/weightReg [11]), .ip2(\STAGE_1/weightReg [10]), .ip3(m1Inputs[92]), .ip4(m1Inputs[91]), .op(n14128) );
  inv_1 U13061 ( .ip(n14128), .op(n13494) );
  or2_1 U13062 ( .ip1(n13493), .ip2(n13494), .op(n13497) );
  nand2_1 U13063 ( .ip1(n14629), .ip2(m1Inputs[92]), .op(n13495) );
  or2_1 U13064 ( .ip1(n13495), .ip2(n13494), .op(n13496) );
  nand2_1 U13065 ( .ip1(n13497), .ip2(n13496), .op(n14126) );
  inv_1 U13066 ( .ip(n14126), .op(n13500) );
  nand2_1 U13067 ( .ip1(column[94]), .ip2(n13498), .op(n13499) );
  mux2_1 U13068 ( .ip1(n13500), .ip2(n14126), .s(n13499), .op(n14080) );
  nor2_1 U13069 ( .ip1(n14842), .ip2(n13748), .op(n14103) );
  nor2_1 U13070 ( .ip1(n12083), .ip2(n13708), .op(n14102) );
  nand2_1 U13071 ( .ip1(m1Inputs[95]), .ip2(n4627), .op(n14101) );
  inv_1 U13072 ( .ip(n13501), .op(n14090) );
  inv_1 U13073 ( .ip(n13502), .op(n13505) );
  nand3_1 U13074 ( .ip1(column[93]), .ip2(n15042), .ip3(n13503), .op(n13504)
         );
  nand2_1 U13075 ( .ip1(n13505), .ip2(n13504), .op(n14110) );
  fulladder U13076 ( .a(n13508), .b(n13507), .ci(n13506), .co(n14109), .s(
        n13418) );
  inv_1 U13077 ( .ip(n13509), .op(n14089) );
  fulladder U13078 ( .a(n13512), .b(n13511), .ci(n13510), .co(n14088), .s(
        n13525) );
  fulladder U13079 ( .a(n13515), .b(n13514), .ci(n13513), .co(n14100), .s(
        n13522) );
  nor2_1 U13080 ( .ip1(n14188), .ip2(n13800), .op(n14093) );
  nor2_1 U13081 ( .ip1(n6503), .ip2(n13675), .op(n14092) );
  nand2_1 U13082 ( .ip1(n14976), .ip2(m1Inputs[87]), .op(n14091) );
  inv_1 U13083 ( .ip(n13516), .op(n14099) );
  fulladder U13084 ( .a(n13519), .b(n13518), .ci(n13517), .co(n14098), .s(
        n13524) );
  fulladder U13085 ( .a(n13522), .b(n13521), .ci(n13520), .co(n14071), .s(
        n13470) );
  fulladder U13086 ( .a(n13525), .b(n13524), .ci(n13523), .co(n14076), .s(
        n13443) );
  fulladder U13087 ( .a(n13528), .b(n13527), .ci(n13526), .co(n13489), .s(
        n13529) );
  inv_1 U13088 ( .ip(n13529), .op(n13617) );
  fulladder U13089 ( .a(n13532), .b(n13531), .ci(n13530), .co(n13523), .s(
        n13533) );
  inv_1 U13090 ( .ip(n13533), .op(n13620) );
  fulladder U13091 ( .a(n13536), .b(n13535), .ci(n13534), .co(n13520), .s(
        n13537) );
  inv_1 U13092 ( .ip(n13537), .op(n13619) );
  fulladder U13093 ( .a(n13540), .b(n13539), .ci(n13538), .co(n13530), .s(
        n13541) );
  inv_1 U13094 ( .ip(n13541), .op(n13559) );
  nand2_1 U13095 ( .ip1(m1Inputs[91]), .ip2(\STAGE_1/weightReg [6]), .op(
        n13542) );
  nor3_1 U13096 ( .ip1(n13800), .ip2(n14289), .ip3(n13584), .op(n13546) );
  or2_1 U13097 ( .ip1(n13542), .ip2(n13546), .op(n13545) );
  nand2_1 U13098 ( .ip1(m1Inputs[90]), .ip2(n4627), .op(n13543) );
  or2_1 U13099 ( .ip1(n13543), .ip2(n13546), .op(n13544) );
  nand2_1 U13100 ( .ip1(n13545), .ip2(n13544), .op(n13577) );
  or2_1 U13101 ( .ip1(n13577), .ip2(n13546), .op(n13548) );
  nor2_1 U13102 ( .ip1(n13853), .ip2(n13835), .op(n13576) );
  or2_1 U13103 ( .ip1(n13576), .ip2(n13546), .op(n13547) );
  nand2_1 U13104 ( .ip1(n13548), .ip2(n13547), .op(n13662) );
  nand2_1 U13105 ( .ip1(m1Inputs[93]), .ip2(n13637), .op(n13668) );
  nor2_1 U13106 ( .ip1(n13830), .ip2(n14853), .op(n13667) );
  nand2_1 U13107 ( .ip1(\STAGE_1/weightReg [8]), .ip2(m1Inputs[89]), .op(
        n13666) );
  xor2_1 U13108 ( .ip1(n13550), .ip2(n13549), .op(n13660) );
  inv_1 U13109 ( .ip(n13551), .op(n13558) );
  nor2_1 U13110 ( .ip1(n14373), .ip2(n13847), .op(n13562) );
  nor2_1 U13111 ( .ip1(n14902), .ip2(n13578), .op(n13561) );
  nor2_1 U13112 ( .ip1(n13766), .ip2(n13748), .op(n13573) );
  and2_1 U13113 ( .ip1(column[89]), .ip2(n13498), .op(n13572) );
  nand2_1 U13114 ( .ip1(column[88]), .ip2(n13859), .op(n13648) );
  inv_1 U13115 ( .ip(n13648), .op(n13571) );
  inv_1 U13116 ( .ip(n13552), .op(n13616) );
  fulladder U13117 ( .a(n13555), .b(n13554), .ci(n13553), .co(n13526), .s(
        n13556) );
  inv_1 U13118 ( .ip(n13556), .op(n13624) );
  fulladder U13119 ( .a(n13559), .b(n13558), .ci(n13557), .co(n13618), .s(
        n13692) );
  fulladder U13120 ( .a(n13562), .b(n13561), .ci(n13560), .co(n13557), .s(
        n13633) );
  nor2_1 U13121 ( .ip1(n13836), .ip2(n14836), .op(n13638) );
  and3_1 U13122 ( .ip1(m1Inputs[90]), .ip2(n14835), .ip3(n13638), .op(n13567)
         );
  nor2_1 U13123 ( .ip1(n13800), .ip2(n14289), .op(n13563) );
  or2_1 U13124 ( .ip1(\STAGE_1/weightReg [7]), .ip2(n13563), .op(n13565) );
  or2_1 U13125 ( .ip1(m1Inputs[89]), .ip2(n13563), .op(n13564) );
  nand2_1 U13126 ( .ip1(n13565), .ip2(n13564), .op(n13566) );
  nor2_1 U13127 ( .ip1(n13567), .ip2(n13566), .op(n13658) );
  or2_1 U13128 ( .ip1(n13658), .ip2(n13567), .op(n13569) );
  nor2_1 U13129 ( .ip1(n13760), .ip2(n4624), .op(n13657) );
  or2_1 U13130 ( .ip1(n13657), .ip2(n13567), .op(n13568) );
  nand2_1 U13131 ( .ip1(n13569), .ip2(n13568), .op(n13696) );
  nand2_1 U13132 ( .ip1(n13614), .ip2(m1Inputs[93]), .op(n13798) );
  nor2_1 U13133 ( .ip1(n13570), .ip2(n13645), .op(n13702) );
  nand2_1 U13134 ( .ip1(m1Inputs[82]), .ip2(\STAGE_1/weightReg [14]), .op(
        n13701) );
  fulladder U13135 ( .a(n13573), .b(n13572), .ci(n13571), .co(n13560), .s(
        n13574) );
  inv_1 U13136 ( .ip(n13574), .op(n13694) );
  inv_1 U13137 ( .ip(n13575), .op(n13632) );
  xor2_1 U13138 ( .ip1(n13577), .ip2(n13576), .op(n13699) );
  nor2_1 U13139 ( .ip1(n13594), .ip2(n13578), .op(n13591) );
  and3_1 U13140 ( .ip1(\STAGE_1/weightReg [11]), .ip2(m1Inputs[87]), .ip3(
        n13591), .op(n13610) );
  nor2_1 U13141 ( .ip1(n13579), .ip2(n13578), .op(n13580) );
  or2_1 U13142 ( .ip1(m1Inputs[87]), .ip2(n13580), .op(n13582) );
  or2_1 U13143 ( .ip1(n14876), .ip2(n13580), .op(n13581) );
  nand2_1 U13144 ( .ip1(n13582), .ip2(n13581), .op(n13583) );
  nor2_1 U13145 ( .ip1(n13610), .ip2(n13583), .op(n13609) );
  nor2_1 U13146 ( .ip1(n14340), .ip2(n13765), .op(n13611) );
  xor2_1 U13147 ( .ip1(n13609), .ip2(n13611), .op(n13698) );
  nor2_1 U13148 ( .ip1(n13853), .ip2(n14783), .op(n13705) );
  nand2_1 U13149 ( .ip1(m1Inputs[81]), .ip2(n14976), .op(n13703) );
  fulladder U13150 ( .a(n13586), .b(n13585), .ci(n13584), .co(n13488), .s(
        n13587) );
  inv_1 U13151 ( .ip(n13587), .op(n13630) );
  fulladder U13152 ( .a(n13590), .b(n13589), .ci(n13588), .co(n13597), .s(
        n13629) );
  nor2_1 U13153 ( .ip1(n14902), .ip2(n13847), .op(n13636) );
  or2_1 U13154 ( .ip1(m1Inputs[85]), .ip2(n13591), .op(n13593) );
  or2_1 U13155 ( .ip1(n13718), .ip2(n13591), .op(n13592) );
  nand2_1 U13156 ( .ip1(n13593), .ip2(n13592), .op(n13652) );
  nor3_1 U13157 ( .ip1(n13652), .ip2(n13654), .ip3(n14373), .op(n13595) );
  nor2_1 U13158 ( .ip1(n13594), .ip2(n13847), .op(n13767) );
  and3_1 U13159 ( .ip1(\STAGE_1/weightReg [11]), .ip2(m1Inputs[86]), .ip3(
        n13767), .op(n13653) );
  or2_1 U13160 ( .ip1(n13595), .ip2(n13653), .op(n13635) );
  nor2_1 U13161 ( .ip1(n13854), .ip2(n13675), .op(n13649) );
  nor2_1 U13162 ( .ip1(n13766), .ip2(n13825), .op(n13647) );
  inv_1 U13163 ( .ip(n13596), .op(n13623) );
  fulladder U13164 ( .a(n13599), .b(n13598), .ci(n13597), .co(n13553), .s(
        n13600) );
  inv_1 U13165 ( .ip(n13600), .op(n13627) );
  fulladder U13166 ( .a(n13603), .b(n13602), .ci(n13601), .co(n13554), .s(
        n13604) );
  inv_1 U13167 ( .ip(n13604), .op(n13626) );
  nor2_1 U13168 ( .ip1(n13606), .ip2(n13605), .op(n13608) );
  xor2_1 U13169 ( .ip1(n13608), .ip2(n13607), .op(n13665) );
  or2_1 U13170 ( .ip1(n13609), .ip2(n13610), .op(n13613) );
  or2_1 U13171 ( .ip1(n13611), .ip2(n13610), .op(n13612) );
  nand2_1 U13172 ( .ip1(n13613), .ip2(n13612), .op(n13664) );
  nor2_1 U13173 ( .ip1(n13854), .ip2(n13645), .op(n13670) );
  nand2_1 U13174 ( .ip1(n13614), .ip2(m1Inputs[94]), .op(n13758) );
  nand2_1 U13175 ( .ip1(m1Inputs[83]), .ip2(\STAGE_1/weightReg [14]), .op(
        n13669) );
  fulladder U13176 ( .a(n13617), .b(n13616), .ci(n13615), .co(n14107), .s(
        n14035) );
  fulladder U13177 ( .a(n13620), .b(n13619), .ci(n13618), .co(n13552), .s(
        n13621) );
  inv_1 U13178 ( .ip(n13621), .op(n13686) );
  fulladder U13179 ( .a(n13624), .b(n13623), .ci(n13622), .co(n13615), .s(
        n13685) );
  fulladder U13180 ( .a(n13627), .b(n13626), .ci(n13625), .co(n13622), .s(
        n13689) );
  fulladder U13181 ( .a(n13630), .b(n13629), .ci(n13628), .co(n13690), .s(
        n13779) );
  fulladder U13182 ( .a(n13633), .b(n13632), .ci(n13631), .co(n13691), .s(
        n13778) );
  fulladder U13183 ( .a(n13636), .b(n13635), .ci(n13634), .co(n13628), .s(
        n13786) );
  nand2_1 U13184 ( .ip1(m1Inputs[89]), .ip2(n13637), .op(n13838) );
  nor3_1 U13185 ( .ip1(n13760), .ip2(n14836), .ip3(n13838), .op(n13642) );
  or2_1 U13186 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n13638), .op(n13640) );
  or2_1 U13187 ( .ip1(m1Inputs[91]), .ip2(n13638), .op(n13639) );
  nand2_1 U13188 ( .ip1(n13640), .ip2(n13639), .op(n13641) );
  nor2_1 U13189 ( .ip1(n13642), .ip2(n13641), .op(n13732) );
  or2_1 U13190 ( .ip1(n13732), .ip2(n13642), .op(n13644) );
  nor2_1 U13191 ( .ip1(n13841), .ip2(n14842), .op(n13731) );
  or2_1 U13192 ( .ip1(n13731), .ip2(n13642), .op(n13643) );
  nand2_1 U13193 ( .ip1(n13644), .ip2(n13643), .op(n13738) );
  nor2_1 U13194 ( .ip1(n13646), .ip2(n13645), .op(n13728) );
  nand2_1 U13195 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[86]), .op(
        n13727) );
  fulladder U13196 ( .a(n13649), .b(n13648), .ci(n13647), .co(n13634), .s(
        n13650) );
  inv_1 U13197 ( .ip(n13650), .op(n13736) );
  inv_1 U13198 ( .ip(n13651), .op(n13785) );
  nor2_1 U13199 ( .ip1(n13653), .ip2(n13652), .op(n13656) );
  nor2_1 U13200 ( .ip1(n13654), .ip2(n14340), .op(n13655) );
  xor2_1 U13201 ( .ip1(n13656), .ip2(n13655), .op(n13735) );
  xor2_1 U13202 ( .ip1(n13658), .ip2(n13657), .op(n13734) );
  nor2_1 U13203 ( .ip1(n13800), .ip2(n13835), .op(n13726) );
  nand2_1 U13204 ( .ip1(m1Inputs[80]), .ip2(n14976), .op(n13725) );
  inv_1 U13205 ( .ip(n13659), .op(n13688) );
  fulladder U13206 ( .a(n13662), .b(n13661), .ci(n13660), .co(n13551), .s(
        n13721) );
  fulladder U13207 ( .a(n13665), .b(n13664), .ci(n13663), .co(n13625), .s(
        n13720) );
  fulladder U13208 ( .a(n13668), .b(n13667), .ci(n13666), .co(n13661), .s(
        n13724) );
  fulladder U13209 ( .a(n13670), .b(n13758), .ci(n13669), .co(n13663), .s(
        n13723) );
  nor2_1 U13210 ( .ip1(n13825), .ip2(n14368), .op(n13750) );
  and2_1 U13211 ( .ip1(n13704), .ip2(n13750), .op(n13755) );
  nor2_1 U13212 ( .ip1(n13748), .ip2(n14384), .op(n13671) );
  or2_1 U13213 ( .ip1(m1Inputs[87]), .ip2(n13671), .op(n13673) );
  or2_1 U13214 ( .ip1(n14838), .ip2(n13671), .op(n13672) );
  nand2_1 U13215 ( .ip1(n13673), .ip2(n13672), .op(n13754) );
  nand2_1 U13216 ( .ip1(m1Inputs[82]), .ip2(n15028), .op(n13756) );
  nor2_1 U13217 ( .ip1(n13754), .ip2(n13756), .op(n13674) );
  nor2_1 U13218 ( .ip1(n13755), .ip2(n13674), .op(n13743) );
  nand2_1 U13219 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[93]), .op(
        n13676) );
  nand2_1 U13220 ( .ip1(n13707), .ip2(m1Inputs[93]), .op(n13711) );
  nor3_1 U13221 ( .ip1(n13854), .ip2(n13675), .ip3(n13711), .op(n13680) );
  or2_1 U13222 ( .ip1(n13676), .ip2(n13680), .op(n13679) );
  nand2_1 U13223 ( .ip1(n13707), .ip2(m1Inputs[94]), .op(n13677) );
  or2_1 U13224 ( .ip1(n13677), .ip2(n13680), .op(n13678) );
  nand2_1 U13225 ( .ip1(n13679), .ip2(n13678), .op(n13773) );
  or2_1 U13226 ( .ip1(n13773), .ip2(n13680), .op(n13683) );
  nand2_1 U13227 ( .ip1(column[87]), .ip2(n13859), .op(n13772) );
  inv_1 U13228 ( .ip(n13772), .op(n13681) );
  or2_1 U13229 ( .ip1(n13681), .ip2(n13680), .op(n13682) );
  nand2_1 U13230 ( .ip1(n13683), .ip2(n13682), .op(n13742) );
  nand2_1 U13231 ( .ip1(n15025), .ip2(m1Inputs[84]), .op(n13741) );
  fulladder U13232 ( .a(n13686), .b(n13685), .ci(n13684), .co(n14034), .s(
        n14039) );
  fulladder U13233 ( .a(n13689), .b(n13688), .ci(n13687), .co(n13684), .s(
        n13776) );
  fulladder U13234 ( .a(n13692), .b(n13691), .ci(n13690), .co(n13596), .s(
        n13693) );
  inv_1 U13235 ( .ip(n13693), .op(n13775) );
  fulladder U13236 ( .a(n13696), .b(n13695), .ci(n13694), .co(n13575), .s(
        n13790) );
  fulladder U13237 ( .a(n13699), .b(n13698), .ci(n13697), .co(n13631), .s(
        n13700) );
  inv_1 U13238 ( .ip(n13700), .op(n13789) );
  fulladder U13239 ( .a(n13798), .b(n13702), .ci(n13701), .co(n13695), .s(
        n13793) );
  fulladder U13240 ( .a(n13705), .b(n13704), .ci(n13703), .co(n13697), .s(
        n13706) );
  inv_1 U13241 ( .ip(n13706), .op(n13792) );
  nand2_1 U13242 ( .ip1(n4672), .ip2(m1Inputs[92]), .op(n13710) );
  nand2_1 U13243 ( .ip1(n13707), .ip2(m1Inputs[92]), .op(n13856) );
  nor3_1 U13244 ( .ip1(n13709), .ip2(n13708), .ip3(n13856), .op(n13714) );
  or2_1 U13245 ( .ip1(n13710), .ip2(n13714), .op(n13713) );
  or2_1 U13246 ( .ip1(n13711), .ip2(n13714), .op(n13712) );
  nand2_1 U13247 ( .ip1(n13713), .ip2(n13712), .op(n13846) );
  or2_1 U13248 ( .ip1(n13846), .ip2(n13714), .op(n13717) );
  nand2_1 U13249 ( .ip1(column[86]), .ip2(n13859), .op(n13845) );
  inv_1 U13250 ( .ip(n13845), .op(n13715) );
  or2_1 U13251 ( .ip1(n13715), .ip2(n13714), .op(n13716) );
  nand2_1 U13252 ( .ip1(n13717), .ip2(n13716), .op(n13823) );
  nand2_1 U13253 ( .ip1(m1Inputs[83]), .ip2(\STAGE_1/weightReg [12]), .op(
        n13822) );
  nand2_1 U13254 ( .ip1(n13718), .ip2(m1Inputs[84]), .op(n13821) );
  fulladder U13255 ( .a(n13721), .b(n13720), .ci(n13719), .co(n13687), .s(
        n13782) );
  fulladder U13256 ( .a(n13724), .b(n13723), .ci(n13722), .co(n13719), .s(
        n13872) );
  fulladder U13257 ( .a(n13726), .b(n13767), .ci(n13725), .co(n13733), .s(
        n13882) );
  fulladder U13258 ( .a(n13729), .b(n13728), .ci(n13727), .co(n13737), .s(
        n13730) );
  inv_1 U13259 ( .ip(n13730), .op(n13881) );
  xor2_1 U13260 ( .ip1(n13732), .ip2(n13731), .op(n13880) );
  fulladder U13261 ( .a(n13735), .b(n13734), .ci(n13733), .co(n13784), .s(
        n13874) );
  fulladder U13262 ( .a(n13738), .b(n13737), .ci(n13736), .co(n13651), .s(
        n13739) );
  inv_1 U13263 ( .ip(n13739), .op(n13873) );
  inv_1 U13264 ( .ip(n13740), .op(n13871) );
  fulladder U13265 ( .a(n13743), .b(n13742), .ci(n13741), .co(n13722), .s(
        n13879) );
  nor3_1 U13266 ( .ip1(n13800), .ip2(n13835), .ip3(n13838), .op(n13898) );
  nor2_1 U13267 ( .ip1(n13836), .ip2(n13835), .op(n13744) );
  or2_1 U13268 ( .ip1(\STAGE_1/weightReg [4]), .ip2(n13744), .op(n13746) );
  or2_1 U13269 ( .ip1(m1Inputs[90]), .ip2(n13744), .op(n13745) );
  nand2_1 U13270 ( .ip1(n13746), .ip2(n13745), .op(n13897) );
  nand2_1 U13271 ( .ip1(n14975), .ip2(m1Inputs[86]), .op(n13899) );
  nor2_1 U13272 ( .ip1(n13897), .ip2(n13899), .op(n13747) );
  nor2_1 U13273 ( .ip1(n13898), .ip2(n13747), .op(n13817) );
  nor3_1 U13274 ( .ip1(n13748), .ip2(n14368), .ip3(n13827), .op(n13795) );
  or2_1 U13275 ( .ip1(n13749), .ip2(n13750), .op(n13752) );
  or2_1 U13276 ( .ip1(m1Inputs[88]), .ip2(n13750), .op(n13751) );
  nand2_1 U13277 ( .ip1(n13752), .ip2(n13751), .op(n13794) );
  nand2_1 U13278 ( .ip1(m1Inputs[81]), .ip2(\STAGE_1/weightReg [13]), .op(
        n13796) );
  nor2_1 U13279 ( .ip1(n13794), .ip2(n13796), .op(n13753) );
  nor2_1 U13280 ( .ip1(n13795), .ip2(n13753), .op(n13816) );
  nor2_1 U13281 ( .ip1(n13755), .ip2(n13754), .op(n13757) );
  xor2_1 U13282 ( .ip1(n13757), .ip2(n13756), .op(n13815) );
  nor2_1 U13283 ( .ip1(n13759), .ip2(n13758), .op(n13902) );
  nor2_1 U13284 ( .ip1(n13801), .ip2(n13760), .op(n13761) );
  or2_1 U13285 ( .ip1(m1Inputs[94]), .ip2(n13761), .op(n13763) );
  or2_1 U13286 ( .ip1(n13803), .ip2(n13761), .op(n13762) );
  nand2_1 U13287 ( .ip1(n13763), .ip2(n13762), .op(n13901) );
  nand2_1 U13288 ( .ip1(m1Inputs[80]), .ip2(n14816), .op(n13903) );
  nor2_1 U13289 ( .ip1(n13901), .ip2(n13903), .op(n13764) );
  nor2_1 U13290 ( .ip1(n13902), .ip2(n13764), .op(n13820) );
  nor2_1 U13291 ( .ip1(n13766), .ip2(n13765), .op(n13848) );
  and2_1 U13292 ( .ip1(n13848), .ip2(n13767), .op(n13812) );
  nor2_1 U13293 ( .ip1(n13766), .ip2(n13847), .op(n13768) );
  or2_1 U13294 ( .ip1(m1Inputs[84]), .ip2(n13768), .op(n13770) );
  or2_1 U13295 ( .ip1(n14876), .ip2(n13768), .op(n13769) );
  nand2_1 U13296 ( .ip1(n13770), .ip2(n13769), .op(n13811) );
  nand2_1 U13297 ( .ip1(m1Inputs[82]), .ip2(n15025), .op(n13813) );
  nor2_1 U13298 ( .ip1(n13811), .ip2(n13813), .op(n13771) );
  nor2_1 U13299 ( .ip1(n13812), .ip2(n13771), .op(n13819) );
  xor2_1 U13300 ( .ip1(n13773), .ip2(n13772), .op(n13818) );
  fulladder U13301 ( .a(n13776), .b(n13775), .ci(n13774), .co(n14038), .s(
        n14043) );
  fulladder U13302 ( .a(n13779), .b(n13778), .ci(n13777), .co(n13659), .s(
        n13780) );
  inv_1 U13303 ( .ip(n13780), .op(n13866) );
  fulladder U13304 ( .a(n13783), .b(n13782), .ci(n13781), .co(n13774), .s(
        n13865) );
  fulladder U13305 ( .a(n13786), .b(n13785), .ci(n13784), .co(n13777), .s(
        n13787) );
  inv_1 U13306 ( .ip(n13787), .op(n13869) );
  fulladder U13307 ( .a(n13790), .b(n13789), .ci(n13788), .co(n13783), .s(
        n13868) );
  fulladder U13308 ( .a(n13793), .b(n13792), .ci(n13791), .co(n13788), .s(
        n13929) );
  nor2_1 U13309 ( .ip1(n13795), .ip2(n13794), .op(n13797) );
  xor2_1 U13310 ( .ip1(n13797), .ip2(n13796), .op(n13945) );
  nor2_1 U13311 ( .ip1(n13799), .ip2(n13798), .op(n13808) );
  nor2_1 U13312 ( .ip1(n13801), .ip2(n13800), .op(n13802) );
  or2_1 U13313 ( .ip1(m1Inputs[93]), .ip2(n13802), .op(n13805) );
  or2_1 U13314 ( .ip1(n13803), .ip2(n13802), .op(n13804) );
  nand2_1 U13315 ( .ip1(n13805), .ip2(n13804), .op(n13806) );
  nor2_1 U13316 ( .ip1(n13808), .ip2(n13806), .op(n13952) );
  or2_1 U13317 ( .ip1(n13952), .ip2(n13808), .op(n13810) );
  nor2_1 U13318 ( .ip1(n13807), .ip2(n14340), .op(n13951) );
  or2_1 U13319 ( .ip1(n13951), .ip2(n13808), .op(n13809) );
  nand2_1 U13320 ( .ip1(n13810), .ip2(n13809), .op(n13944) );
  nor2_1 U13321 ( .ip1(n13812), .ip2(n13811), .op(n13814) );
  xor2_1 U13322 ( .ip1(n13814), .ip2(n13813), .op(n13943) );
  fulladder U13323 ( .a(n13817), .b(n13816), .ci(n13815), .co(n13878), .s(
        n13940) );
  fulladder U13324 ( .a(n13820), .b(n13819), .ci(n13818), .co(n13877), .s(
        n13939) );
  fulladder U13325 ( .a(n13823), .b(n13822), .ci(n13821), .co(n13791), .s(
        n13937) );
  nand2_1 U13326 ( .ip1(m1Inputs[86]), .ip2(n4627), .op(n13826) );
  nor3_1 U13327 ( .ip1(n13825), .ip2(n14368), .ip3(n13824), .op(n13831) );
  or2_1 U13328 ( .ip1(n13826), .ip2(n13831), .op(n13829) );
  or2_1 U13329 ( .ip1(n13827), .ip2(n13831), .op(n13828) );
  nand2_1 U13330 ( .ip1(n13829), .ip2(n13828), .op(n13956) );
  or2_1 U13331 ( .ip1(n13956), .ip2(n13831), .op(n13833) );
  nor2_1 U13332 ( .ip1(n13830), .ip2(n14824), .op(n13955) );
  or2_1 U13333 ( .ip1(n13955), .ip2(n13831), .op(n13832) );
  nand2_1 U13334 ( .ip1(n13833), .ip2(n13832), .op(n13910) );
  nand2_1 U13335 ( .ip1(m1Inputs[88]), .ip2(\STAGE_1/weightReg [5]), .op(
        n13837) );
  nor3_1 U13336 ( .ip1(n13836), .ip2(n13835), .ip3(n13834), .op(n13842) );
  or2_1 U13337 ( .ip1(n13837), .ip2(n13842), .op(n13840) );
  or2_1 U13338 ( .ip1(n13838), .ip2(n13842), .op(n13839) );
  nand2_1 U13339 ( .ip1(n13840), .ip2(n13839), .op(n13954) );
  or2_1 U13340 ( .ip1(n13954), .ip2(n13842), .op(n13844) );
  nor2_1 U13341 ( .ip1(n13841), .ip2(n14902), .op(n13953) );
  or2_1 U13342 ( .ip1(n13953), .ip2(n13842), .op(n13843) );
  nand2_1 U13343 ( .ip1(n13844), .ip2(n13843), .op(n13909) );
  xor2_1 U13344 ( .ip1(n13846), .ip2(n13845), .op(n13908) );
  nor3_1 U13345 ( .ip1(n13766), .ip2(n13847), .ip3(n13984), .op(n13921) );
  or2_1 U13346 ( .ip1(m1Inputs[85]), .ip2(n13848), .op(n13850) );
  or2_1 U13347 ( .ip1(n14838), .ip2(n13848), .op(n13849) );
  nand2_1 U13348 ( .ip1(n13850), .ip2(n13849), .op(n13920) );
  nand2_1 U13349 ( .ip1(m1Inputs[83]), .ip2(\STAGE_1/weightReg [10]), .op(
        n13922) );
  nor2_1 U13350 ( .ip1(n13920), .ip2(n13922), .op(n13851) );
  nor2_1 U13351 ( .ip1(n13921), .ip2(n13851), .op(n13907) );
  nand2_1 U13352 ( .ip1(\STAGE_1/weightReg [2]), .ip2(m1Inputs[91]), .op(
        n13855) );
  nor3_1 U13353 ( .ip1(n13854), .ip2(n13853), .ip3(n13852), .op(n13860) );
  or2_1 U13354 ( .ip1(n13855), .ip2(n13860), .op(n13858) );
  or2_1 U13355 ( .ip1(n13856), .ip2(n13860), .op(n13857) );
  nand2_1 U13356 ( .ip1(n13858), .ip2(n13857), .op(n13896) );
  or2_1 U13357 ( .ip1(n13896), .ip2(n13860), .op(n13863) );
  nand2_1 U13358 ( .ip1(column[85]), .ip2(n13859), .op(n13895) );
  inv_1 U13359 ( .ip(n13895), .op(n13861) );
  or2_1 U13360 ( .ip1(n13861), .ip2(n13860), .op(n13862) );
  nand2_1 U13361 ( .ip1(n13863), .ip2(n13862), .op(n13906) );
  nand2_1 U13362 ( .ip1(m1Inputs[83]), .ip2(\STAGE_1/weightReg [11]), .op(
        n13905) );
  fulladder U13363 ( .a(n13866), .b(n13865), .ci(n13864), .co(n14042), .s(
        n14047) );
  fulladder U13364 ( .a(n13869), .b(n13868), .ci(n13867), .co(n13864), .s(
        n13926) );
  fulladder U13365 ( .a(n13872), .b(n13871), .ci(n13870), .co(n13781), .s(
        n13925) );
  fulladder U13366 ( .a(n13875), .b(n13874), .ci(n13873), .co(n13740), .s(
        n13876) );
  inv_1 U13367 ( .ip(n13876), .op(n13933) );
  fulladder U13368 ( .a(n13879), .b(n13878), .ci(n13877), .co(n13870), .s(
        n13932) );
  fulladder U13369 ( .a(n13882), .b(n13881), .ci(n13880), .co(n13875), .s(
        n13883) );
  inv_1 U13370 ( .ip(n13883), .op(n13968) );
  or2_1 U13371 ( .ip1(n13884), .ip2(n13886), .op(n13889) );
  inv_1 U13372 ( .ip(n13885), .op(n13887) );
  or2_1 U13373 ( .ip1(n13887), .ip2(n13886), .op(n13888) );
  nand2_1 U13374 ( .ip1(n13889), .ip2(n13888), .op(n13978) );
  or2_1 U13375 ( .ip1(n13890), .ip2(n13891), .op(n13894) );
  or2_1 U13376 ( .ip1(n13892), .ip2(n13891), .op(n13893) );
  nand2_1 U13377 ( .ip1(n13894), .ip2(n13893), .op(n13977) );
  xor2_1 U13378 ( .ip1(n13896), .ip2(n13895), .op(n13976) );
  nor2_1 U13379 ( .ip1(n13898), .ip2(n13897), .op(n13900) );
  xor2_1 U13380 ( .ip1(n13900), .ip2(n13899), .op(n13948) );
  nor2_1 U13381 ( .ip1(n13902), .ip2(n13901), .op(n13904) );
  xor2_1 U13382 ( .ip1(n13904), .ip2(n13903), .op(n13947) );
  fulladder U13383 ( .a(n13907), .b(n13906), .ci(n13905), .co(n13935), .s(
        n13981) );
  fulladder U13384 ( .a(n13910), .b(n13909), .ci(n13908), .co(n13936), .s(
        n13980) );
  or2_1 U13385 ( .ip1(n13911), .ip2(n13912), .op(n13915) );
  or2_1 U13386 ( .ip1(n13913), .ip2(n13912), .op(n13914) );
  nand2_1 U13387 ( .ip1(n13915), .ip2(n13914), .op(n13971) );
  nor2_1 U13388 ( .ip1(n13917), .ip2(n13916), .op(n13918) );
  nor2_1 U13389 ( .ip1(n13919), .ip2(n13918), .op(n13970) );
  nor2_1 U13390 ( .ip1(n13921), .ip2(n13920), .op(n13923) );
  xor2_1 U13391 ( .ip1(n13923), .ip2(n13922), .op(n13969) );
  fulladder U13392 ( .a(n13926), .b(n13925), .ci(n13924), .co(n14046), .s(
        n14051) );
  fulladder U13393 ( .a(n13929), .b(n13928), .ci(n13927), .co(n13867), .s(
        n13930) );
  inv_1 U13394 ( .ip(n13930), .op(n13960) );
  fulladder U13395 ( .a(n13933), .b(n13932), .ci(n13931), .co(n13924), .s(
        n13934) );
  inv_1 U13396 ( .ip(n13934), .op(n13959) );
  fulladder U13397 ( .a(n13937), .b(n13936), .ci(n13935), .co(n13927), .s(
        n13938) );
  inv_1 U13398 ( .ip(n13938), .op(n13964) );
  fulladder U13399 ( .a(n13941), .b(n13940), .ci(n13939), .co(n13928), .s(
        n13942) );
  inv_1 U13400 ( .ip(n13942), .op(n13963) );
  fulladder U13401 ( .a(n13945), .b(n13944), .ci(n13943), .co(n13941), .s(
        n13946) );
  inv_1 U13402 ( .ip(n13946), .op(n13996) );
  fulladder U13403 ( .a(n13949), .b(n13948), .ci(n13947), .co(n13967), .s(
        n13950) );
  inv_1 U13404 ( .ip(n13950), .op(n13995) );
  xor2_1 U13405 ( .ip1(n13952), .ip2(n13951), .op(n13974) );
  xor2_1 U13406 ( .ip1(n13954), .ip2(n13953), .op(n13973) );
  xor2_1 U13407 ( .ip1(n13956), .ip2(n13955), .op(n13972) );
  inv_1 U13408 ( .ip(n13957), .op(n14050) );
  fulladder U13409 ( .a(n13960), .b(n13959), .ci(n13958), .co(n13957), .s(
        n13961) );
  inv_1 U13410 ( .ip(n13961), .op(n14055) );
  fulladder U13411 ( .a(n13964), .b(n13963), .ci(n13962), .co(n13958), .s(
        n13965) );
  inv_1 U13412 ( .ip(n13965), .op(n13993) );
  fulladder U13413 ( .a(n13968), .b(n13967), .ci(n13966), .co(n13931), .s(
        n13992) );
  fulladder U13414 ( .a(n13971), .b(n13970), .ci(n13969), .co(n13979), .s(
        n14015) );
  fulladder U13415 ( .a(n13974), .b(n13973), .ci(n13972), .co(n13994), .s(
        n13975) );
  inv_1 U13416 ( .ip(n13975), .op(n14014) );
  fulladder U13417 ( .a(n13978), .b(n13977), .ci(n13976), .co(n13949), .s(
        n14013) );
  fulladder U13418 ( .a(n13981), .b(n13980), .ci(n13979), .co(n13966), .s(
        n13999) );
  fulladder U13419 ( .a(n13984), .b(n13983), .ci(n13982), .co(n14003), .s(
        n14005) );
  fulladder U13420 ( .a(n13987), .b(n13986), .ci(n13985), .co(n14002), .s(
        n14009) );
  fulladder U13421 ( .a(n13990), .b(n13989), .ci(n13988), .co(n14001), .s(
        n14021) );
  fulladder U13422 ( .a(n13993), .b(n13992), .ci(n13991), .co(n14054), .s(
        n14059) );
  fulladder U13423 ( .a(n13996), .b(n13995), .ci(n13994), .co(n13962), .s(
        n13997) );
  inv_1 U13424 ( .ip(n13997), .op(n14012) );
  fulladder U13425 ( .a(n14000), .b(n13999), .ci(n13998), .co(n13991), .s(
        n14011) );
  fulladder U13426 ( .a(n14003), .b(n14002), .ci(n14001), .co(n13998), .s(
        n14018) );
  fulladder U13427 ( .a(n14006), .b(n14005), .ci(n14004), .co(n14017), .s(
        n14020) );
  fulladder U13428 ( .a(n14009), .b(n14008), .ci(n14007), .co(n14016), .s(
        n14031) );
  fulladder U13429 ( .a(n14012), .b(n14011), .ci(n14010), .co(n14058), .s(
        n14063) );
  fulladder U13430 ( .a(n14015), .b(n14014), .ci(n14013), .co(n14000), .s(
        n14024) );
  fulladder U13431 ( .a(n14018), .b(n14017), .ci(n14016), .co(n14010), .s(
        n14023) );
  fulladder U13432 ( .a(n14021), .b(n14020), .ci(n14019), .co(n14022), .s(
        n14030) );
  fulladder U13433 ( .a(n14024), .b(n14023), .ci(n14022), .co(n14062), .s(
        n14067) );
  fulladder U13434 ( .a(n14027), .b(n14026), .ci(n14025), .co(n14028), .s(
        \STAGE_1/M6/sum [4]) );
  inv_1 U13435 ( .ip(n14028), .op(n14066) );
  fulladder U13436 ( .a(n14031), .b(n14030), .ci(n14029), .co(n14065), .s(
        n13410) );
  inv_1 U13437 ( .ip(n14032), .op(\STAGE_1/M6/sum [14]) );
  fulladder U13438 ( .a(n14035), .b(n14034), .ci(n14033), .co(n14106), .s(
        n14036) );
  inv_1 U13439 ( .ip(n14036), .op(\STAGE_1/M6/sum [13]) );
  fulladder U13440 ( .a(n14039), .b(n14038), .ci(n14037), .co(n14033), .s(
        n14040) );
  inv_1 U13441 ( .ip(n14040), .op(\STAGE_1/M6/sum [12]) );
  fulladder U13442 ( .a(n14043), .b(n14042), .ci(n14041), .co(n14037), .s(
        n14044) );
  inv_1 U13443 ( .ip(n14044), .op(\STAGE_1/M6/sum [11]) );
  fulladder U13444 ( .a(n14047), .b(n14046), .ci(n14045), .co(n14041), .s(
        n14048) );
  inv_1 U13445 ( .ip(n14048), .op(\STAGE_1/M6/sum [10]) );
  fulladder U13446 ( .a(n14051), .b(n14050), .ci(n14049), .co(n14045), .s(
        n14052) );
  inv_1 U13447 ( .ip(n14052), .op(\STAGE_1/M6/sum [9]) );
  fulladder U13448 ( .a(n14055), .b(n14054), .ci(n14053), .co(n14049), .s(
        n14056) );
  inv_1 U13449 ( .ip(n14056), .op(\STAGE_1/M6/sum [8]) );
  fulladder U13450 ( .a(n14059), .b(n14058), .ci(n14057), .co(n14053), .s(
        n14060) );
  inv_1 U13451 ( .ip(n14060), .op(\STAGE_1/M6/sum [7]) );
  fulladder U13452 ( .a(n14063), .b(n14062), .ci(n14061), .co(n14057), .s(
        n14064) );
  inv_1 U13453 ( .ip(n14064), .op(\STAGE_1/M6/sum [6]) );
  fulladder U13454 ( .a(n14067), .b(n14066), .ci(n14065), .co(n14061), .s(
        n14068) );
  inv_1 U13455 ( .ip(n14068), .op(\STAGE_1/M6/sum [5]) );
  nand2_1 U13456 ( .ip1(m1Inputs[95]), .ip2(n14975), .op(n14070) );
  nand2_1 U13457 ( .ip1(m1Inputs[89]), .ip2(\STAGE_1/weightReg [14]), .op(
        n14069) );
  xor2_1 U13458 ( .ip1(n14070), .ip2(n14069), .op(n14075) );
  fulladder U13459 ( .a(n14073), .b(n14072), .ci(n14071), .co(n14074), .s(
        n14077) );
  xor2_1 U13460 ( .ip1(n14075), .ip2(n14074), .op(n14085) );
  fulladder U13461 ( .a(n14078), .b(n14077), .ci(n14076), .co(n14083), .s(
        n14108) );
  fulladder U13462 ( .a(n14081), .b(n14080), .ci(n14079), .co(n14082), .s(
        n13501) );
  xor2_1 U13463 ( .ip1(n14083), .ip2(n14082), .op(n14084) );
  xor2_1 U13464 ( .ip1(n14085), .ip2(n14084), .op(n14087) );
  nand2_1 U13465 ( .ip1(m1Inputs[91]), .ip2(\STAGE_1/weightReg [12]), .op(
        n14086) );
  xor2_1 U13466 ( .ip1(n14087), .ip2(n14086), .op(n14132) );
  fulladder U13467 ( .a(n14090), .b(n14089), .ci(n14088), .co(n14095), .s(
        n14073) );
  fulladder U13468 ( .a(n14093), .b(n14092), .ci(n14091), .co(n14094), .s(
        n13516) );
  xor2_1 U13469 ( .ip1(n14095), .ip2(n14094), .op(n14096) );
  xor2_1 U13470 ( .ip1(n14097), .ip2(n14096), .op(n14125) );
  fulladder U13471 ( .a(n14100), .b(n14099), .ci(n14098), .co(n14105), .s(
        n14072) );
  fulladder U13472 ( .a(n14103), .b(n14102), .ci(n14101), .co(n14104), .s(
        n14079) );
  xor2_1 U13473 ( .ip1(n14105), .ip2(n14104), .op(n14115) );
  fulladder U13474 ( .a(n14108), .b(n14107), .ci(n14106), .co(n14113), .s(
        n14032) );
  fulladder U13475 ( .a(n14111), .b(n14110), .ci(n14109), .co(n14112), .s(
        n13509) );
  xor2_1 U13476 ( .ip1(n14113), .ip2(n14112), .op(n14114) );
  xor2_1 U13477 ( .ip1(n14115), .ip2(n14114), .op(n14123) );
  nand2_1 U13478 ( .ip1(m1Inputs[90]), .ip2(\STAGE_1/weightReg [13]), .op(
        n14117) );
  nand2_1 U13479 ( .ip1(m1Inputs[88]), .ip2(\STAGE_1/weightReg [15]), .op(
        n14116) );
  xor2_1 U13480 ( .ip1(n14117), .ip2(n14116), .op(n14121) );
  nand2_1 U13481 ( .ip1(m1Inputs[94]), .ip2(n14994), .op(n14119) );
  nand2_1 U13482 ( .ip1(m1Inputs[93]), .ip2(\STAGE_1/weightReg [10]), .op(
        n14118) );
  xor2_1 U13483 ( .ip1(n14119), .ip2(n14118), .op(n14120) );
  xor2_1 U13484 ( .ip1(n14121), .ip2(n14120), .op(n14122) );
  xor2_1 U13485 ( .ip1(n14123), .ip2(n14122), .op(n14124) );
  xor2_1 U13486 ( .ip1(n14125), .ip2(n14124), .op(n14130) );
  nand3_1 U13487 ( .ip1(column[94]), .ip2(n15042), .ip3(n14126), .op(n14127)
         );
  nand2_1 U13488 ( .ip1(n14128), .ip2(n14127), .op(n14129) );
  xor2_1 U13489 ( .ip1(n14130), .ip2(n14129), .op(n14131) );
  xor2_1 U13490 ( .ip1(n14132), .ip2(n14131), .op(n14134) );
  nand2_1 U13491 ( .ip1(n15042), .ip2(column[95]), .op(n14133) );
  xor2_1 U13492 ( .ip1(n14134), .ip2(n14133), .op(\STAGE_1/M6/sum [15]) );
  fulladder U13493 ( .a(n14137), .b(n14136), .ci(n14135), .co(n7684), .s(
        n14138) );
  inv_1 U13494 ( .ip(n14138), .op(\STAGE_1/M7/sum [12]) );
  fulladder U13495 ( .a(n14141), .b(n14140), .ci(n14139), .co(n14135), .s(
        n14142) );
  inv_1 U13496 ( .ip(n14142), .op(\STAGE_1/M7/sum [11]) );
  fulladder U13497 ( .a(n14145), .b(n14144), .ci(n14143), .co(n14139), .s(
        n14146) );
  inv_1 U13498 ( .ip(n14146), .op(\STAGE_1/M7/sum [10]) );
  fulladder U13499 ( .a(n14149), .b(n14148), .ci(n14147), .co(n14143), .s(
        n14150) );
  inv_1 U13500 ( .ip(n14150), .op(\STAGE_1/M7/sum [9]) );
  fulladder U13501 ( .a(n14153), .b(n14152), .ci(n14151), .co(n14147), .s(
        n14154) );
  inv_1 U13502 ( .ip(n14154), .op(\STAGE_1/M7/sum [8]) );
  fulladder U13503 ( .a(n14157), .b(n14156), .ci(n14155), .co(n14151), .s(
        n14158) );
  inv_1 U13504 ( .ip(n14158), .op(\STAGE_1/M7/sum [7]) );
  fulladder U13505 ( .a(n14161), .b(n14160), .ci(n14159), .co(n14211), .s(
        n14198) );
  nand4_1 U13506 ( .ip1(\STAGE_1/weightReg [11]), .ip2(\STAGE_1/weightReg [10]), .ip3(m1Inputs[108]), .ip4(m1Inputs[107]), .op(n14266) );
  inv_1 U13507 ( .ip(n14266), .op(n14163) );
  or2_1 U13508 ( .ip1(n14162), .ip2(n14163), .op(n14166) );
  nand2_1 U13509 ( .ip1(n14629), .ip2(m1Inputs[108]), .op(n14164) );
  or2_1 U13510 ( .ip1(n14164), .ip2(n14163), .op(n14165) );
  nand2_1 U13511 ( .ip1(n14166), .ip2(n14165), .op(n14264) );
  inv_1 U13512 ( .ip(n14264), .op(n14168) );
  nand2_1 U13513 ( .ip1(column[110]), .ip2(n14768), .op(n14167) );
  mux2_1 U13514 ( .ip1(n14168), .ip2(n14264), .s(n14167), .op(n14219) );
  nor2_1 U13515 ( .ip1(n14842), .ip2(n14169), .op(n14216) );
  nor2_1 U13516 ( .ip1(n12083), .ip2(n14170), .op(n14215) );
  nand2_1 U13517 ( .ip1(m1Inputs[111]), .ip2(\STAGE_1/weightReg [7]), .op(
        n14214) );
  fulladder U13518 ( .a(n14173), .b(n14172), .ci(n14171), .co(n14217), .s(
        n14182) );
  inv_1 U13519 ( .ip(n14174), .op(n14177) );
  nand3_1 U13520 ( .ip1(column[109]), .ip2(n15042), .ip3(n14175), .op(n14176)
         );
  nand2_1 U13521 ( .ip1(n14177), .ip2(n14176), .op(n14235) );
  fulladder U13522 ( .a(n14180), .b(n14179), .ci(n14178), .co(n14234), .s(
        n14183) );
  fulladder U13523 ( .a(n14183), .b(n14182), .ci(n14181), .co(n14242), .s(
        n7035) );
  fulladder U13524 ( .a(n14186), .b(n14185), .ci(n14184), .co(n14228), .s(
        n14195) );
  nor2_1 U13525 ( .ip1(n14188), .ip2(n14187), .op(n14247) );
  nor2_1 U13526 ( .ip1(n6503), .ip2(n14189), .op(n14246) );
  nand2_1 U13527 ( .ip1(n14976), .ip2(m1Inputs[103]), .op(n14245) );
  fulladder U13528 ( .a(n14192), .b(n14191), .ci(n14190), .co(n14226), .s(
        n7049) );
  fulladder U13529 ( .a(n14195), .b(n14194), .ci(n14193), .co(n14237), .s(
        n7031) );
  inv_1 U13530 ( .ip(n14196), .op(n14210) );
  fulladder U13531 ( .a(n14199), .b(n14198), .ci(n14197), .co(n14209), .s(
        n7068) );
  inv_1 U13532 ( .ip(n14200), .op(n14231) );
  fulladder U13533 ( .a(n14203), .b(n14202), .ci(n14201), .co(n14230), .s(
        n14206) );
  fulladder U13534 ( .a(n14206), .b(n14205), .ci(n14204), .co(n14229), .s(
        \STAGE_1/M7/sum [13]) );
  nand2_1 U13535 ( .ip1(m1Inputs[110]), .ip2(n14994), .op(n14208) );
  nand2_1 U13536 ( .ip1(m1Inputs[104]), .ip2(\STAGE_1/weightReg [15]), .op(
        n14207) );
  xor2_1 U13537 ( .ip1(n14208), .ip2(n14207), .op(n14213) );
  fulladder U13538 ( .a(n14211), .b(n14210), .ci(n14209), .co(n14212), .s(
        n14200) );
  xor2_1 U13539 ( .ip1(n14213), .ip2(n14212), .op(n14223) );
  fulladder U13540 ( .a(n14216), .b(n14215), .ci(n14214), .co(n14221), .s(
        n14218) );
  fulladder U13541 ( .a(n14219), .b(n14218), .ci(n14217), .co(n14220), .s(
        n14244) );
  xor2_1 U13542 ( .ip1(n14221), .ip2(n14220), .op(n14222) );
  xor2_1 U13543 ( .ip1(n14223), .ip2(n14222), .op(n14225) );
  nand2_1 U13544 ( .ip1(m1Inputs[107]), .ip2(\STAGE_1/weightReg [12]), .op(
        n14224) );
  xor2_1 U13545 ( .ip1(n14225), .ip2(n14224), .op(n14270) );
  fulladder U13546 ( .a(n14228), .b(n14227), .ci(n14226), .co(n14255), .s(
        n14238) );
  fulladder U13547 ( .a(n14231), .b(n14230), .ci(n14229), .co(n14233), .s(
        \STAGE_1/M7/sum [14]) );
  nand2_1 U13548 ( .ip1(m1Inputs[105]), .ip2(\STAGE_1/weightReg [14]), .op(
        n14232) );
  xor2_1 U13549 ( .ip1(n14233), .ip2(n14232), .op(n14253) );
  fulladder U13550 ( .a(n14236), .b(n14235), .ci(n14234), .co(n14241), .s(
        n14243) );
  fulladder U13551 ( .a(n14239), .b(n14238), .ci(n14237), .co(n14240), .s(
        n14196) );
  xor2_1 U13552 ( .ip1(n14241), .ip2(n14240), .op(n14251) );
  fulladder U13553 ( .a(n14244), .b(n14243), .ci(n14242), .co(n14249), .s(
        n14239) );
  fulladder U13554 ( .a(n14247), .b(n14246), .ci(n14245), .co(n14248), .s(
        n14227) );
  xor2_1 U13555 ( .ip1(n14249), .ip2(n14248), .op(n14250) );
  xor2_1 U13556 ( .ip1(n14251), .ip2(n14250), .op(n14252) );
  xor2_1 U13557 ( .ip1(n14253), .ip2(n14252), .op(n14254) );
  xor2_1 U13558 ( .ip1(n14255), .ip2(n14254), .op(n14263) );
  nand2_1 U13559 ( .ip1(m1Inputs[111]), .ip2(n14975), .op(n14257) );
  nand2_1 U13560 ( .ip1(m1Inputs[106]), .ip2(\STAGE_1/weightReg [13]), .op(
        n14256) );
  xor2_1 U13561 ( .ip1(n14257), .ip2(n14256), .op(n14258) );
  xor2_1 U13562 ( .ip1(n14259), .ip2(n14258), .op(n14261) );
  nand2_1 U13563 ( .ip1(n14876), .ip2(m1Inputs[109]), .op(n14260) );
  xor2_1 U13564 ( .ip1(n14261), .ip2(n14260), .op(n14262) );
  xor2_1 U13565 ( .ip1(n14263), .ip2(n14262), .op(n14268) );
  nand3_1 U13566 ( .ip1(column[110]), .ip2(n15042), .ip3(n14264), .op(n14265)
         );
  nand2_1 U13567 ( .ip1(n14266), .ip2(n14265), .op(n14267) );
  xor2_1 U13568 ( .ip1(n14268), .ip2(n14267), .op(n14269) );
  xor2_1 U13569 ( .ip1(n14270), .ip2(n14269), .op(n14272) );
  nand2_1 U13570 ( .ip1(n15042), .ip2(column[111]), .op(n14271) );
  xor2_1 U13571 ( .ip1(n14272), .ip2(n14271), .op(\STAGE_1/M7/sum [15]) );
  nand2_1 U13572 ( .ip1(n14629), .ip2(m1Inputs[122]), .op(n14377) );
  nor2_1 U13573 ( .ip1(n14377), .ip2(n14276), .op(n14364) );
  nor2_1 U13574 ( .ip1(n13766), .ip2(n14433), .op(n14341) );
  or2_1 U13575 ( .ip1(m1Inputs[121]), .ip2(n14341), .op(n14274) );
  or2_1 U13576 ( .ip1(n14876), .ip2(n14341), .op(n14273) );
  nand2_1 U13577 ( .ip1(n14274), .ip2(n14273), .op(n14362) );
  or2_1 U13578 ( .ip1(n14364), .ip2(n14362), .op(n14275) );
  nand2_1 U13579 ( .ip1(column[123]), .ip2(n14768), .op(n14361) );
  xor2_1 U13580 ( .ip1(n14275), .ip2(n14361), .op(n14406) );
  fulladder U13581 ( .a(n14278), .b(n14277), .ci(n14276), .co(n14279), .s(
        n7748) );
  inv_1 U13582 ( .ip(n14279), .op(n14405) );
  fulladder U13583 ( .a(n14282), .b(n14281), .ci(n14280), .co(n14404), .s(
        n14326) );
  inv_1 U13584 ( .ip(n14283), .op(n14471) );
  nand2_1 U13585 ( .ip1(m1Inputs[119]), .ip2(\STAGE_1/weightReg [12]), .op(
        n14285) );
  nand2_1 U13586 ( .ip1(m1Inputs[120]), .ip2(\STAGE_1/weightReg [11]), .op(
        n14284) );
  xor2_1 U13587 ( .ip1(n14285), .ip2(n14284), .op(n14350) );
  nor2_1 U13588 ( .ip1(n14842), .ip2(n14286), .op(n14352) );
  xor2_1 U13589 ( .ip1(n14350), .ip2(n14352), .op(n14403) );
  nand2_1 U13590 ( .ip1(m1Inputs[124]), .ip2(\STAGE_1/weightReg [7]), .op(
        n14357) );
  nor2_1 U13591 ( .ip1(n14287), .ip2(n14783), .op(n14356) );
  nand2_1 U13592 ( .ip1(m1Inputs[126]), .ip2(n14369), .op(n14355) );
  inv_1 U13593 ( .ip(n14288), .op(n14402) );
  nor2_1 U13594 ( .ip1(n14419), .ip2(n14289), .op(n14367) );
  nor2_1 U13595 ( .ip1(n6503), .ip2(n14290), .op(n14366) );
  nand2_1 U13596 ( .ip1(n14976), .ip2(m1Inputs[116]), .op(n14365) );
  inv_1 U13597 ( .ip(n14291), .op(n14470) );
  fulladder U13598 ( .a(n14294), .b(n14293), .ci(n14292), .co(n14469), .s(
        n14300) );
  fulladder U13599 ( .a(n14297), .b(n14296), .ci(n14295), .co(n14298), .s(
        n7795) );
  inv_1 U13600 ( .ip(n14298), .op(n14483) );
  fulladder U13601 ( .a(n14301), .b(n14300), .ci(n14299), .co(n14482), .s(
        n14329) );
  and3_1 U13602 ( .ip1(\STAGE_1/weightReg [10]), .ip2(m1Inputs[122]), .ip3(
        n14302), .op(n14305) );
  or2_1 U13603 ( .ip1(n14303), .ip2(n14305), .op(n14308) );
  inv_1 U13604 ( .ip(n14304), .op(n14306) );
  or2_1 U13605 ( .ip1(n14306), .ip2(n14305), .op(n14307) );
  nand2_1 U13606 ( .ip1(n14308), .ip2(n14307), .op(n14396) );
  nand2_1 U13607 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[118]), .op(
        n14395) );
  nor2_1 U13608 ( .ip1(n14310), .ip2(n14309), .op(n14311) );
  nor2_1 U13609 ( .ip1(n14312), .ip2(n14311), .op(n14394) );
  inv_1 U13610 ( .ip(n14313), .op(n14459) );
  fulladder U13611 ( .a(n14316), .b(n14315), .ci(n14314), .co(n14317), .s(
        n14301) );
  inv_1 U13612 ( .ip(n14317), .op(n14458) );
  fulladder U13613 ( .a(n14320), .b(n14319), .ci(n14318), .co(n14457), .s(
        n14323) );
  fulladder U13614 ( .a(n14323), .b(n14322), .ci(n14321), .co(n14466), .s(
        n14296) );
  fulladder U13615 ( .a(n14326), .b(n14325), .ci(n14324), .co(n14465), .s(
        n14297) );
  inv_1 U13616 ( .ip(n14327), .op(n14493) );
  fulladder U13617 ( .a(n14330), .b(n14329), .ci(n14328), .co(n14492), .s(
        n14333) );
  inv_1 U13618 ( .ip(n14331), .op(n14490) );
  fulladder U13619 ( .a(n14334), .b(n14333), .ci(n14332), .co(n14335), .s(
        n7956) );
  inv_1 U13620 ( .ip(n14335), .op(n14489) );
  fulladder U13621 ( .a(n14338), .b(n14337), .ci(n14336), .co(n14488), .s(
        \STAGE_1/M8/sum [10]) );
  nor2_1 U13622 ( .ip1(n14842), .ip2(n14339), .op(n14432) );
  nor2_1 U13623 ( .ip1(n14340), .ip2(n14418), .op(n14431) );
  nand3_1 U13624 ( .ip1(n14629), .ip2(m1Inputs[123]), .ip3(n14341), .op(n14346) );
  nand2_1 U13625 ( .ip1(m1Inputs[123]), .ip2(n14994), .op(n14342) );
  nand2_1 U13626 ( .ip1(n14342), .ip2(n14377), .op(n14343) );
  nand2_1 U13627 ( .ip1(n14343), .ip2(n14346), .op(n14360) );
  inv_1 U13628 ( .ip(n14360), .op(n14344) );
  nand3_1 U13629 ( .ip1(column[124]), .ip2(n15042), .ip3(n14344), .op(n14345)
         );
  nand2_1 U13630 ( .ip1(n14346), .ip2(n14345), .op(n14430) );
  nand2_1 U13631 ( .ip1(m1Inputs[119]), .ip2(\STAGE_1/weightReg [13]), .op(
        n14348) );
  nand2_1 U13632 ( .ip1(m1Inputs[121]), .ip2(\STAGE_1/weightReg [11]), .op(
        n14347) );
  xor2_1 U13633 ( .ip1(n14348), .ip2(n14347), .op(n14371) );
  nand2_1 U13634 ( .ip1(n14816), .ip2(m1Inputs[118]), .op(n14349) );
  xor2_1 U13635 ( .ip1(n14371), .ip2(n14349), .op(n14455) );
  nor2_1 U13636 ( .ip1(n14902), .ip2(n14418), .op(n14387) );
  and2_1 U13637 ( .ip1(n14374), .ip2(n14387), .op(n14351) );
  or2_1 U13638 ( .ip1(n14350), .ip2(n14351), .op(n14354) );
  or2_1 U13639 ( .ip1(n14352), .ip2(n14351), .op(n14353) );
  nand2_1 U13640 ( .ip1(n14354), .ip2(n14353), .op(n14454) );
  fulladder U13641 ( .a(n14357), .b(n14356), .ci(n14355), .co(n14453), .s(
        n14288) );
  inv_1 U13642 ( .ip(n14358), .op(n14439) );
  nand2_1 U13643 ( .ip1(column[124]), .ip2(n14768), .op(n14359) );
  xor2_1 U13644 ( .ip1(n14360), .ip2(n14359), .op(n14400) );
  nor2_1 U13645 ( .ip1(n14362), .ip2(n14361), .op(n14363) );
  or2_1 U13646 ( .ip1(n14364), .ip2(n14363), .op(n14399) );
  fulladder U13647 ( .a(n14367), .b(n14366), .ci(n14365), .co(n14398), .s(
        n14401) );
  nor2_1 U13648 ( .ip1(n13766), .ip2(n14517), .op(n14426) );
  nor2_1 U13649 ( .ip1(n14434), .ip2(n14368), .op(n14425) );
  nand2_1 U13650 ( .ip1(n14976), .ip2(m1Inputs[118]), .op(n14424) );
  nor2_1 U13651 ( .ip1(n14902), .ip2(n14372), .op(n14410) );
  nor2_1 U13652 ( .ip1(n6503), .ip2(n14419), .op(n14409) );
  nand2_1 U13653 ( .ip1(m1Inputs[127]), .ip2(n12981), .op(n14408) );
  nor2_1 U13654 ( .ip1(n14434), .ip2(n14836), .op(n14392) );
  nor2_1 U13655 ( .ip1(n6503), .ip2(n14517), .op(n14391) );
  nand2_1 U13656 ( .ip1(m1Inputs[127]), .ip2(n14369), .op(n14390) );
  inv_1 U13657 ( .ip(n14370), .op(n14444) );
  nand3_1 U13658 ( .ip1(n14816), .ip2(n14371), .ip3(m1Inputs[118]), .op(n14376) );
  nor2_1 U13659 ( .ip1(n14373), .ip2(n14372), .op(n14562) );
  nand2_1 U13660 ( .ip1(n14374), .ip2(n14562), .op(n14375) );
  nand2_1 U13661 ( .ip1(n14376), .ip2(n14375), .op(n14437) );
  nand2_1 U13662 ( .ip1(n14629), .ip2(m1Inputs[123]), .op(n14378) );
  nand2_1 U13663 ( .ip1(n14847), .ip2(m1Inputs[123]), .op(n14411) );
  nor2_1 U13664 ( .ip1(n14411), .ip2(n14377), .op(n14420) );
  or2_1 U13665 ( .ip1(n14378), .ip2(n14420), .op(n14381) );
  nand2_1 U13666 ( .ip1(n14847), .ip2(m1Inputs[122]), .op(n14379) );
  or2_1 U13667 ( .ip1(n14379), .ip2(n14420), .op(n14380) );
  nand2_1 U13668 ( .ip1(n14381), .ip2(n14380), .op(n14421) );
  inv_1 U13669 ( .ip(n14421), .op(n14383) );
  nand2_1 U13670 ( .ip1(column[125]), .ip2(n14768), .op(n14382) );
  mux2_1 U13671 ( .ip1(n14383), .ip2(n14421), .s(n14382), .op(n14436) );
  nor2_1 U13672 ( .ip1(n14419), .ip2(n14384), .op(n14388) );
  nand2_1 U13673 ( .ip1(n14976), .ip2(m1Inputs[117]), .op(n14386) );
  inv_1 U13674 ( .ip(n14385), .op(n14443) );
  fulladder U13675 ( .a(n14388), .b(n14387), .ci(n14386), .co(n14435), .s(
        n14389) );
  inv_1 U13676 ( .ip(n14389), .op(n14451) );
  fulladder U13677 ( .a(n14392), .b(n14391), .ci(n14390), .co(n14427), .s(
        n14393) );
  inv_1 U13678 ( .ip(n14393), .op(n14450) );
  fulladder U13679 ( .a(n14396), .b(n14395), .ci(n14394), .co(n14449), .s(
        n14313) );
  inv_1 U13680 ( .ip(n14397), .op(n14446) );
  fulladder U13681 ( .a(n14400), .b(n14399), .ci(n14398), .co(n14438), .s(
        n14463) );
  fulladder U13682 ( .a(n14403), .b(n14402), .ci(n14401), .co(n14462), .s(
        n14291) );
  fulladder U13683 ( .a(n14406), .b(n14405), .ci(n14404), .co(n14461), .s(
        n14283) );
  inv_1 U13684 ( .ip(n14407), .op(n14554) );
  fulladder U13685 ( .a(n14410), .b(n14409), .ci(n14408), .co(n14531), .s(
        n14428) );
  nand4_1 U13686 ( .ip1(\STAGE_1/weightReg [11]), .ip2(\STAGE_1/weightReg [10]), .ip3(m1Inputs[124]), .ip4(m1Inputs[123]), .op(n14505) );
  inv_1 U13687 ( .ip(n14505), .op(n14412) );
  or2_1 U13688 ( .ip1(n14411), .ip2(n14412), .op(n14415) );
  nand2_1 U13689 ( .ip1(n14629), .ip2(m1Inputs[124]), .op(n14413) );
  or2_1 U13690 ( .ip1(n14413), .ip2(n14412), .op(n14414) );
  nand2_1 U13691 ( .ip1(n14415), .ip2(n14414), .op(n14504) );
  inv_1 U13692 ( .ip(n14504), .op(n14417) );
  nand2_1 U13693 ( .ip1(column[126]), .ip2(n14768), .op(n14416) );
  mux2_1 U13694 ( .ip1(n14417), .ip2(n14504), .s(n14416), .op(n14530) );
  nor2_1 U13695 ( .ip1(n14842), .ip2(n14418), .op(n14520) );
  nor2_1 U13696 ( .ip1(n12083), .ip2(n14419), .op(n14519) );
  nand2_1 U13697 ( .ip1(m1Inputs[127]), .ip2(n14835), .op(n14518) );
  inv_1 U13698 ( .ip(n14420), .op(n14423) );
  nand3_1 U13699 ( .ip1(column[125]), .ip2(n15042), .ip3(n14421), .op(n14422)
         );
  nand2_1 U13700 ( .ip1(n14423), .ip2(n14422), .op(n14561) );
  fulladder U13701 ( .a(n14426), .b(n14425), .ci(n14424), .co(n14560), .s(
        n14429) );
  fulladder U13702 ( .a(n14429), .b(n14428), .ci(n14427), .co(n14526), .s(
        n14370) );
  fulladder U13703 ( .a(n14432), .b(n14431), .ci(n14430), .co(n14514), .s(
        n14440) );
  nor2_1 U13704 ( .ip1(n14902), .ip2(n14433), .op(n14559) );
  nor2_1 U13705 ( .ip1(n6504), .ip2(n14434), .op(n14558) );
  nand2_1 U13706 ( .ip1(n14976), .ip2(m1Inputs[119]), .op(n14557) );
  fulladder U13707 ( .a(n14437), .b(n14436), .ci(n14435), .co(n14512), .s(
        n14385) );
  fulladder U13708 ( .a(n14440), .b(n14439), .ci(n14438), .co(n14509), .s(
        n14447) );
  inv_1 U13709 ( .ip(n14441), .op(n14553) );
  fulladder U13710 ( .a(n14444), .b(n14443), .ci(n14442), .co(n14552), .s(
        n14397) );
  fulladder U13711 ( .a(n14447), .b(n14446), .ci(n14445), .co(n14407), .s(
        n14448) );
  inv_1 U13712 ( .ip(n14448), .op(n14474) );
  fulladder U13713 ( .a(n14451), .b(n14450), .ci(n14449), .co(n14442), .s(
        n14452) );
  inv_1 U13714 ( .ip(n14452), .op(n14477) );
  fulladder U13715 ( .a(n14455), .b(n14454), .ci(n14453), .co(n14358), .s(
        n14456) );
  inv_1 U13716 ( .ip(n14456), .op(n14476) );
  fulladder U13717 ( .a(n14459), .b(n14458), .ci(n14457), .co(n14475), .s(
        n14467) );
  inv_1 U13718 ( .ip(n14460), .op(n14473) );
  fulladder U13719 ( .a(n14463), .b(n14462), .ci(n14461), .co(n14445), .s(
        n14464) );
  inv_1 U13720 ( .ip(n14464), .op(n14481) );
  fulladder U13721 ( .a(n14467), .b(n14466), .ci(n14465), .co(n14468), .s(
        n14327) );
  inv_1 U13722 ( .ip(n14468), .op(n14480) );
  fulladder U13723 ( .a(n14471), .b(n14470), .ci(n14469), .co(n14479), .s(
        n14484) );
  fulladder U13724 ( .a(n14474), .b(n14473), .ci(n14472), .co(n14522), .s(
        n14498) );
  fulladder U13725 ( .a(n14477), .b(n14476), .ci(n14475), .co(n14460), .s(
        n14478) );
  inv_1 U13726 ( .ip(n14478), .op(n14487) );
  fulladder U13727 ( .a(n14481), .b(n14480), .ci(n14479), .co(n14472), .s(
        n14486) );
  fulladder U13728 ( .a(n14484), .b(n14483), .ci(n14482), .co(n14485), .s(
        n14494) );
  fulladder U13729 ( .a(n14487), .b(n14486), .ci(n14485), .co(n14497), .s(
        n14502) );
  fulladder U13730 ( .a(n14490), .b(n14489), .ci(n14488), .co(n14491), .s(
        \STAGE_1/M8/sum [11]) );
  inv_1 U13731 ( .ip(n14491), .op(n14501) );
  fulladder U13732 ( .a(n14494), .b(n14493), .ci(n14492), .co(n14500), .s(
        n14331) );
  inv_1 U13733 ( .ip(n14495), .op(\STAGE_1/M8/sum [14]) );
  fulladder U13734 ( .a(n14498), .b(n14497), .ci(n14496), .co(n14521), .s(
        n14499) );
  inv_1 U13735 ( .ip(n14499), .op(\STAGE_1/M8/sum [13]) );
  fulladder U13736 ( .a(n14502), .b(n14501), .ci(n14500), .co(n14496), .s(
        n14503) );
  inv_1 U13737 ( .ip(n14503), .op(\STAGE_1/M8/sum [12]) );
  nand2_1 U13738 ( .ip1(column[127]), .ip2(n14768), .op(n14508) );
  nand3_1 U13739 ( .ip1(column[126]), .ip2(n15042), .ip3(n14504), .op(n14506)
         );
  nand2_1 U13740 ( .ip1(n14506), .ip2(n14505), .op(n14507) );
  xor2_1 U13741 ( .ip1(n14508), .ip2(n14507), .op(n14541) );
  fulladder U13742 ( .a(n14511), .b(n14510), .ci(n14509), .co(n14516), .s(
        n14441) );
  fulladder U13743 ( .a(n14514), .b(n14513), .ci(n14512), .co(n14515), .s(
        n14510) );
  xor2_1 U13744 ( .ip1(n14516), .ip2(n14515), .op(n14539) );
  nor2_1 U13745 ( .ip1(n14824), .ip2(n14517), .op(n14537) );
  fulladder U13746 ( .a(n14520), .b(n14519), .ci(n14518), .co(n14525), .s(
        n14529) );
  fulladder U13747 ( .a(n14523), .b(n14522), .ci(n14521), .co(n14524), .s(
        n14495) );
  xor2_1 U13748 ( .ip1(n14525), .ip2(n14524), .op(n14535) );
  fulladder U13749 ( .a(n14528), .b(n14527), .ci(n14526), .co(n14533), .s(
        n14511) );
  fulladder U13750 ( .a(n14531), .b(n14530), .ci(n14529), .co(n14532), .s(
        n14528) );
  xor2_1 U13751 ( .ip1(n14533), .ip2(n14532), .op(n14534) );
  xor2_1 U13752 ( .ip1(n14535), .ip2(n14534), .op(n14536) );
  xor2_1 U13753 ( .ip1(n14537), .ip2(n14536), .op(n14538) );
  xor2_1 U13754 ( .ip1(n14539), .ip2(n14538), .op(n14540) );
  xor2_1 U13755 ( .ip1(n14541), .ip2(n14540), .op(n14549) );
  nand2_1 U13756 ( .ip1(m1Inputs[122]), .ip2(n15028), .op(n14543) );
  nand2_1 U13757 ( .ip1(m1Inputs[125]), .ip2(\STAGE_1/weightReg [10]), .op(
        n14542) );
  xor2_1 U13758 ( .ip1(n14543), .ip2(n14542), .op(n14547) );
  nand2_1 U13759 ( .ip1(m1Inputs[127]), .ip2(n14975), .op(n14545) );
  nand2_1 U13760 ( .ip1(m1Inputs[120]), .ip2(\STAGE_1/weightReg [15]), .op(
        n14544) );
  xor2_1 U13761 ( .ip1(n14545), .ip2(n14544), .op(n14546) );
  xor2_1 U13762 ( .ip1(n14547), .ip2(n14546), .op(n14548) );
  xor2_1 U13763 ( .ip1(n14549), .ip2(n14548), .op(n14570) );
  nand2_1 U13764 ( .ip1(m1Inputs[121]), .ip2(\STAGE_1/weightReg [14]), .op(
        n14551) );
  nand2_1 U13765 ( .ip1(m1Inputs[123]), .ip2(\STAGE_1/weightReg [12]), .op(
        n14550) );
  xor2_1 U13766 ( .ip1(n14551), .ip2(n14550), .op(n14556) );
  fulladder U13767 ( .a(n14554), .b(n14553), .ci(n14552), .co(n14555), .s(
        n14523) );
  xor2_1 U13768 ( .ip1(n14556), .ip2(n14555), .op(n14566) );
  fulladder U13769 ( .a(n14559), .b(n14558), .ci(n14557), .co(n14564), .s(
        n14513) );
  fulladder U13770 ( .a(n14562), .b(n14561), .ci(n14560), .co(n14563), .s(
        n14527) );
  xor2_1 U13771 ( .ip1(n14564), .ip2(n14563), .op(n14565) );
  xor2_1 U13772 ( .ip1(n14566), .ip2(n14565), .op(n14568) );
  nand2_1 U13773 ( .ip1(m1Inputs[126]), .ip2(n14994), .op(n14567) );
  xor2_1 U13774 ( .ip1(n14568), .ip2(n14567), .op(n14569) );
  xor2_1 U13775 ( .ip1(n14570), .ip2(n14569), .op(\STAGE_1/M8/sum [15]) );
  nand2_1 U13776 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[136]), .op(
        n14649) );
  and3_1 U13777 ( .ip1(column[140]), .ip2(n13039), .ip3(n14571), .op(n14572)
         );
  nor2_1 U13778 ( .ip1(n14573), .ip2(n14572), .op(n14648) );
  nand2_1 U13779 ( .ip1(n14816), .ip2(m1Inputs[135]), .op(n14647) );
  fulladder U13780 ( .a(n14576), .b(n14575), .ci(n14574), .co(n14657), .s(
        n8997) );
  fulladder U13781 ( .a(n14579), .b(n14578), .ci(n14577), .co(n14656), .s(
        n9099) );
  inv_1 U13782 ( .ip(n14580), .op(n14623) );
  nand2_1 U13783 ( .ip1(m1Inputs[142]), .ip2(n14835), .op(n14643) );
  nor2_1 U13784 ( .ip1(n14853), .ip2(n14587), .op(n14642) );
  nand2_1 U13785 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[140]), .op(
        n14641) );
  nand2_1 U13786 ( .ip1(n14838), .ip2(m1Inputs[141]), .op(n14627) );
  nor2_1 U13787 ( .ip1(n14581), .ip2(n14836), .op(n14626) );
  nand2_1 U13788 ( .ip1(n15025), .ip2(m1Inputs[137]), .op(n14625) );
  fulladder U13789 ( .a(n14584), .b(n14583), .ci(n14582), .co(n14644), .s(
        n14600) );
  nand2_1 U13790 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[137]), .op(
        n14712) );
  nor2_1 U13791 ( .ip1(n14585), .ip2(n14712), .op(n14589) );
  nor3_1 U13792 ( .ip1(n14842), .ip2(n14587), .ip3(n14586), .op(n14588) );
  nor2_1 U13793 ( .ip1(n14589), .ip2(n14588), .op(n14655) );
  nand2_1 U13794 ( .ip1(n14847), .ip2(m1Inputs[139]), .op(n14628) );
  nor2_1 U13795 ( .ip1(n14628), .ip2(n14590), .op(n14640) );
  or2_1 U13796 ( .ip1(n14591), .ip2(n14640), .op(n14594) );
  nand2_1 U13797 ( .ip1(n14847), .ip2(m1Inputs[138]), .op(n14592) );
  or2_1 U13798 ( .ip1(n14592), .ip2(n14640), .op(n14593) );
  nand2_1 U13799 ( .ip1(n14594), .ip2(n14593), .op(n14638) );
  nand2_1 U13800 ( .ip1(column[141]), .ip2(n14768), .op(n14595) );
  xor2_1 U13801 ( .ip1(n14638), .ip2(n14595), .op(n14654) );
  fulladder U13802 ( .a(n14598), .b(n14597), .ci(n14596), .co(n14653), .s(
        n14601) );
  fulladder U13803 ( .a(n14601), .b(n14600), .ci(n14599), .co(n14659), .s(
        n9090) );
  inv_1 U13804 ( .ip(n14602), .op(n14622) );
  fulladder U13805 ( .a(n14605), .b(n14604), .ci(n14603), .co(n14621), .s(
        n9015) );
  inv_1 U13806 ( .ip(n14606), .op(n14668) );
  fulladder U13807 ( .a(n14609), .b(n14608), .ci(n14607), .co(n14610), .s(
        n14616) );
  inv_1 U13808 ( .ip(n14610), .op(n14667) );
  fulladder U13809 ( .a(n14613), .b(n14612), .ci(n14611), .co(n14666), .s(
        n9086) );
  inv_1 U13810 ( .ip(n14614), .op(n14664) );
  fulladder U13811 ( .a(n14617), .b(n14616), .ci(n14615), .co(n14663), .s(
        n14620) );
  fulladder U13812 ( .a(n14620), .b(n14619), .ci(n14618), .co(n14662), .s(
        \STAGE_1/M9/sum [12]) );
  fulladder U13813 ( .a(n14623), .b(n14622), .ci(n14621), .co(n14624), .s(
        n14606) );
  inv_1 U13814 ( .ip(n14624), .op(n14709) );
  fulladder U13815 ( .a(n14627), .b(n14626), .ci(n14625), .co(n14694), .s(
        n14645) );
  nand4_1 U13816 ( .ip1(\STAGE_1/weightReg [11]), .ip2(n14876), .ip3(
        m1Inputs[140]), .ip4(m1Inputs[139]), .op(n14733) );
  inv_1 U13817 ( .ip(n14733), .op(n14630) );
  or2_1 U13818 ( .ip1(n14628), .ip2(n14630), .op(n14633) );
  nand2_1 U13819 ( .ip1(n14629), .ip2(m1Inputs[140]), .op(n14631) );
  or2_1 U13820 ( .ip1(n14631), .ip2(n14630), .op(n14632) );
  nand2_1 U13821 ( .ip1(n14633), .ip2(n14632), .op(n14731) );
  nand2_1 U13822 ( .ip1(column[142]), .ip2(n14768), .op(n14634) );
  xor2_1 U13823 ( .ip1(n14731), .ip2(n14634), .op(n14693) );
  nor2_1 U13824 ( .ip1(n14842), .ip2(n14635), .op(n14701) );
  nor2_1 U13825 ( .ip1(n13766), .ip2(n14636), .op(n14700) );
  nand2_1 U13826 ( .ip1(m1Inputs[143]), .ip2(n14835), .op(n14699) );
  inv_1 U13827 ( .ip(n14637), .op(n14692) );
  and3_1 U13828 ( .ip1(column[141]), .ip2(n14768), .ip3(n14638), .op(n14639)
         );
  nor2_1 U13829 ( .ip1(n14640), .ip2(n14639), .op(n14711) );
  fulladder U13830 ( .a(n14643), .b(n14642), .ci(n14641), .co(n14710), .s(
        n14646) );
  fulladder U13831 ( .a(n14646), .b(n14645), .ci(n14644), .co(n14689), .s(
        n14661) );
  fulladder U13832 ( .a(n14649), .b(n14648), .ci(n14647), .co(n14674), .s(
        n14658) );
  nor2_1 U13833 ( .ip1(n14902), .ip2(n14650), .op(n14704) );
  nor2_1 U13834 ( .ip1(n6503), .ip2(n14651), .op(n14703) );
  nand2_1 U13835 ( .ip1(n14976), .ip2(m1Inputs[135]), .op(n14702) );
  inv_1 U13836 ( .ip(n14652), .op(n14673) );
  fulladder U13837 ( .a(n14655), .b(n14654), .ci(n14653), .co(n14672), .s(
        n14660) );
  fulladder U13838 ( .a(n14658), .b(n14657), .ci(n14656), .co(n14677), .s(
        n14580) );
  fulladder U13839 ( .a(n14661), .b(n14660), .ci(n14659), .co(n14707), .s(
        n14602) );
  fulladder U13840 ( .a(n14664), .b(n14663), .ci(n14662), .co(n14665), .s(
        \STAGE_1/M9/sum [13]) );
  inv_1 U13841 ( .ip(n14665), .op(n14681) );
  fulladder U13842 ( .a(n14668), .b(n14667), .ci(n14666), .co(n14680), .s(
        n14614) );
  inv_1 U13843 ( .ip(n14669), .op(\STAGE_1/M9/sum [14]) );
  nand2_1 U13844 ( .ip1(m1Inputs[137]), .ip2(\STAGE_1/weightReg [14]), .op(
        n14671) );
  nand2_1 U13845 ( .ip1(m1Inputs[139]), .ip2(\STAGE_1/weightReg [12]), .op(
        n14670) );
  xor2_1 U13846 ( .ip1(n14671), .ip2(n14670), .op(n14676) );
  fulladder U13847 ( .a(n14674), .b(n14673), .ci(n14672), .co(n14675), .s(
        n14678) );
  xor2_1 U13848 ( .ip1(n14676), .ip2(n14675), .op(n14686) );
  fulladder U13849 ( .a(n14679), .b(n14678), .ci(n14677), .co(n14684), .s(
        n14708) );
  fulladder U13850 ( .a(n14682), .b(n14681), .ci(n14680), .co(n14683), .s(
        n14669) );
  xor2_1 U13851 ( .ip1(n14684), .ip2(n14683), .op(n14685) );
  xor2_1 U13852 ( .ip1(n14686), .ip2(n14685), .op(n14688) );
  nand2_1 U13853 ( .ip1(m1Inputs[142]), .ip2(n14994), .op(n14687) );
  xor2_1 U13854 ( .ip1(n14688), .ip2(n14687), .op(n14730) );
  fulladder U13855 ( .a(n14691), .b(n14690), .ci(n14689), .co(n14696), .s(
        n14679) );
  fulladder U13856 ( .a(n14694), .b(n14693), .ci(n14692), .co(n14695), .s(
        n14691) );
  xor2_1 U13857 ( .ip1(n14696), .ip2(n14695), .op(n14697) );
  xor2_1 U13858 ( .ip1(n14698), .ip2(n14697), .op(n14726) );
  fulladder U13859 ( .a(n14701), .b(n14700), .ci(n14699), .co(n14706), .s(
        n14637) );
  fulladder U13860 ( .a(n14704), .b(n14703), .ci(n14702), .co(n14705), .s(
        n14652) );
  xor2_1 U13861 ( .ip1(n14706), .ip2(n14705), .op(n14716) );
  fulladder U13862 ( .a(n14709), .b(n14708), .ci(n14707), .co(n14714), .s(
        n14682) );
  fulladder U13863 ( .a(n14712), .b(n14711), .ci(n14710), .co(n14713), .s(
        n14690) );
  xor2_1 U13864 ( .ip1(n14714), .ip2(n14713), .op(n14715) );
  xor2_1 U13865 ( .ip1(n14716), .ip2(n14715), .op(n14724) );
  nand2_1 U13866 ( .ip1(m1Inputs[143]), .ip2(n14975), .op(n14718) );
  nand2_1 U13867 ( .ip1(m1Inputs[136]), .ip2(\STAGE_1/weightReg [15]), .op(
        n14717) );
  xor2_1 U13868 ( .ip1(n14718), .ip2(n14717), .op(n14722) );
  nand2_1 U13869 ( .ip1(m1Inputs[138]), .ip2(n15028), .op(n14720) );
  nand2_1 U13870 ( .ip1(m1Inputs[141]), .ip2(\STAGE_1/weightReg [10]), .op(
        n14719) );
  xor2_1 U13871 ( .ip1(n14720), .ip2(n14719), .op(n14721) );
  xor2_1 U13872 ( .ip1(n14722), .ip2(n14721), .op(n14723) );
  xor2_1 U13873 ( .ip1(n14724), .ip2(n14723), .op(n14725) );
  xor2_1 U13874 ( .ip1(n14726), .ip2(n14725), .op(n14728) );
  nand2_1 U13875 ( .ip1(n15042), .ip2(column[143]), .op(n14727) );
  xor2_1 U13876 ( .ip1(n14728), .ip2(n14727), .op(n14729) );
  xor2_1 U13877 ( .ip1(n14730), .ip2(n14729), .op(n14735) );
  nand3_1 U13878 ( .ip1(column[142]), .ip2(n15042), .ip3(n14731), .op(n14732)
         );
  nand2_1 U13879 ( .ip1(n14733), .ip2(n14732), .op(n14734) );
  xor2_1 U13880 ( .ip1(n14735), .ip2(n14734), .op(\STAGE_1/M9/sum [15]) );
  nand2_1 U13881 ( .ip1(n14876), .ip2(m1Inputs[154]), .op(n14845) );
  nor3_1 U13882 ( .ip1(n6503), .ip2(n14882), .ip3(n14845), .op(n14738) );
  and3_1 U13883 ( .ip1(column[154]), .ip2(n15042), .ip3(n14736), .op(n14737)
         );
  nor2_1 U13884 ( .ip1(n14738), .ip2(n14737), .op(n14862) );
  nand2_1 U13885 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[150]), .op(
        n14861) );
  or2_1 U13886 ( .ip1(n14739), .ip2(n14740), .op(n14743) );
  or2_1 U13887 ( .ip1(n14741), .ip2(n14740), .op(n14742) );
  nand2_1 U13888 ( .ip1(n14743), .ip2(n14742), .op(n14860) );
  inv_1 U13889 ( .ip(n14744), .op(n14928) );
  fulladder U13890 ( .a(n14747), .b(n14746), .ci(n14745), .co(n14748), .s(
        n14794) );
  inv_1 U13891 ( .ip(n14748), .op(n14927) );
  fulladder U13892 ( .a(n14751), .b(n14750), .ci(n14749), .co(n14926), .s(
        n14754) );
  fulladder U13893 ( .a(n14754), .b(n14753), .ci(n14752), .co(n14935), .s(
        n14797) );
  fulladder U13894 ( .a(n14757), .b(n14756), .ci(n14755), .co(n14934), .s(
        n14798) );
  inv_1 U13895 ( .ip(n14758), .op(n14965) );
  fulladder U13896 ( .a(n14761), .b(n14760), .ci(n14759), .co(n14873), .s(
        n14756) );
  nand2_1 U13897 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[154]), .op(
        n14762) );
  nor3_1 U13898 ( .ip1(n12083), .ip2(n14825), .ip3(n14845), .op(n14818) );
  or2_1 U13899 ( .ip1(n14762), .ip2(n14818), .op(n14765) );
  nand2_1 U13900 ( .ip1(n14876), .ip2(m1Inputs[153]), .op(n14763) );
  or2_1 U13901 ( .ip1(n14763), .ip2(n14818), .op(n14764) );
  nand2_1 U13902 ( .ip1(n14765), .ip2(n14764), .op(n14766) );
  inv_1 U13903 ( .ip(n14766), .op(n14767) );
  and3_1 U13904 ( .ip1(column[155]), .ip2(n15042), .ip3(n14766), .op(n14817)
         );
  or2_1 U13905 ( .ip1(n14767), .ip2(n14817), .op(n14771) );
  nand2_1 U13906 ( .ip1(column[155]), .ip2(n14768), .op(n14769) );
  or2_1 U13907 ( .ip1(n14769), .ip2(n14817), .op(n14770) );
  nand2_1 U13908 ( .ip1(n14771), .ip2(n14770), .op(n14872) );
  fulladder U13909 ( .a(n14774), .b(n14773), .ci(n14772), .co(n14871), .s(
        n14757) );
  inv_1 U13910 ( .ip(n14775), .op(n14940) );
  nand2_1 U13911 ( .ip1(m1Inputs[152]), .ip2(\STAGE_1/weightReg [11]), .op(
        n14778) );
  nor2_1 U13912 ( .ip1(n14902), .ip2(n14776), .op(n14777) );
  xor2_1 U13913 ( .ip1(n14778), .ip2(n14777), .op(n14779) );
  nor3_1 U13914 ( .ip1(n14842), .ip2(n14852), .ip3(n14779), .op(n14829) );
  or2_1 U13915 ( .ip1(n14779), .ip2(n14829), .op(n14782) );
  nand2_1 U13916 ( .ip1(n14816), .ip2(m1Inputs[149]), .op(n14780) );
  or2_1 U13917 ( .ip1(n14780), .ip2(n14829), .op(n14781) );
  nand2_1 U13918 ( .ip1(n14782), .ip2(n14781), .op(n14870) );
  nor2_1 U13919 ( .ip1(n14837), .ip2(n14783), .op(n14833) );
  nand2_1 U13920 ( .ip1(m1Inputs[156]), .ip2(n14835), .op(n14832) );
  nand2_1 U13921 ( .ip1(m1Inputs[158]), .ip2(\STAGE_1/weightReg [5]), .op(
        n14831) );
  inv_1 U13922 ( .ip(n14784), .op(n14869) );
  nand2_1 U13923 ( .ip1(m1Inputs[157]), .ip2(n12981), .op(n14821) );
  nor2_1 U13924 ( .ip1(n14853), .ip2(n14785), .op(n14820) );
  nand2_1 U13925 ( .ip1(n14838), .ip2(m1Inputs[155]), .op(n14819) );
  inv_1 U13926 ( .ip(n14786), .op(n14868) );
  inv_1 U13927 ( .ip(n14787), .op(n14939) );
  fulladder U13928 ( .a(n14790), .b(n14789), .ci(n14788), .co(n14938), .s(
        n14793) );
  inv_1 U13929 ( .ip(n14791), .op(n14953) );
  fulladder U13930 ( .a(n14794), .b(n14793), .ci(n14792), .co(n14795), .s(
        n14802) );
  inv_1 U13931 ( .ip(n14795), .op(n14952) );
  fulladder U13932 ( .a(n14798), .b(n14797), .ci(n14796), .co(n14951), .s(
        n8413) );
  inv_1 U13933 ( .ip(n14799), .op(n14964) );
  fulladder U13934 ( .a(n14802), .b(n14801), .ci(n14800), .co(n14963), .s(
        n14805) );
  inv_1 U13935 ( .ip(n14803), .op(n14961) );
  fulladder U13936 ( .a(n14806), .b(n14805), .ci(n14804), .co(n14807), .s(
        n8577) );
  inv_1 U13937 ( .ip(n14807), .op(n14960) );
  fulladder U13938 ( .a(n14810), .b(n14809), .ci(n14808), .co(n14959), .s(
        \STAGE_1/M10/sum [10]) );
  nand2_1 U13939 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[152]), .op(
        n14900) );
  nand2_1 U13940 ( .ip1(\STAGE_1/weightReg [10]), .ip2(m1Inputs[155]), .op(
        n14846) );
  nor3_1 U13941 ( .ip1(n12083), .ip2(n14846), .ip3(n14901), .op(n14815) );
  or2_1 U13942 ( .ip1(n14845), .ip2(n14815), .op(n14813) );
  nand2_1 U13943 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[155]), .op(
        n14811) );
  or2_1 U13944 ( .ip1(n14811), .ip2(n14815), .op(n14812) );
  nand2_1 U13945 ( .ip1(n14813), .ip2(n14812), .op(n14823) );
  and3_1 U13946 ( .ip1(column[156]), .ip2(n13859), .ip3(n14823), .op(n14814)
         );
  nor2_1 U13947 ( .ip1(n14815), .ip2(n14814), .op(n14899) );
  nand2_1 U13948 ( .ip1(n14816), .ip2(m1Inputs[151]), .op(n14898) );
  nor2_1 U13949 ( .ip1(n14818), .ip2(n14817), .op(n14866) );
  fulladder U13950 ( .a(n14821), .b(n14820), .ci(n14819), .co(n14865), .s(
        n14786) );
  nand2_1 U13951 ( .ip1(column[156]), .ip2(n13498), .op(n14822) );
  xor2_1 U13952 ( .ip1(n14823), .ip2(n14822), .op(n14864) );
  nor2_1 U13953 ( .ip1(n14842), .ip2(n14841), .op(n14828) );
  nor2_1 U13954 ( .ip1(n14825), .ip2(n14824), .op(n14827) );
  nand2_1 U13955 ( .ip1(m1Inputs[151]), .ip2(n15028), .op(n14826) );
  xor2_1 U13956 ( .ip1(n14827), .ip2(n14826), .op(n14840) );
  xor2_1 U13957 ( .ip1(n14828), .ip2(n14840), .op(n14924) );
  nand2_1 U13958 ( .ip1(n15025), .ip2(m1Inputs[152]), .op(n14855) );
  nor2_1 U13959 ( .ip1(n14839), .ip2(n14855), .op(n14830) );
  nor2_1 U13960 ( .ip1(n14830), .ip2(n14829), .op(n14923) );
  fulladder U13961 ( .a(n14833), .b(n14832), .ci(n14831), .co(n14922), .s(
        n14784) );
  inv_1 U13962 ( .ip(n14834), .op(n14916) );
  nand2_1 U13963 ( .ip1(m1Inputs[158]), .ip2(n14835), .op(n14894) );
  nor2_1 U13964 ( .ip1(n14853), .ip2(n14841), .op(n14893) );
  nand2_1 U13965 ( .ip1(\STAGE_1/weightReg [9]), .ip2(m1Inputs[156]), .op(
        n14892) );
  nand2_1 U13966 ( .ip1(n14838), .ip2(m1Inputs[157]), .op(n14888) );
  nor2_1 U13967 ( .ip1(n14837), .ip2(n14836), .op(n14887) );
  nand2_1 U13968 ( .ip1(n15025), .ip2(m1Inputs[153]), .op(n14886) );
  nor2_1 U13969 ( .ip1(n14837), .ip2(n13835), .op(n14859) );
  nand2_1 U13970 ( .ip1(m1Inputs[158]), .ip2(n12981), .op(n14858) );
  nand2_1 U13971 ( .ip1(n14838), .ip2(m1Inputs[156]), .op(n14857) );
  nand2_1 U13972 ( .ip1(\STAGE_1/weightReg [13]), .ip2(m1Inputs[153]), .op(
        n15002) );
  nor2_1 U13973 ( .ip1(n14839), .ip2(n15002), .op(n14844) );
  nor3_1 U13974 ( .ip1(n14842), .ip2(n14841), .ip3(n14840), .op(n14843) );
  nor2_1 U13975 ( .ip1(n14844), .ip2(n14843), .op(n14907) );
  nand2_1 U13976 ( .ip1(n14847), .ip2(m1Inputs[155]), .op(n14875) );
  nor2_1 U13977 ( .ip1(n14875), .ip2(n14845), .op(n14891) );
  or2_1 U13978 ( .ip1(n14846), .ip2(n14891), .op(n14850) );
  nand2_1 U13979 ( .ip1(n14847), .ip2(m1Inputs[154]), .op(n14848) );
  or2_1 U13980 ( .ip1(n14848), .ip2(n14891), .op(n14849) );
  nand2_1 U13981 ( .ip1(n14850), .ip2(n14849), .op(n14889) );
  nand2_1 U13982 ( .ip1(column[157]), .ip2(n15042), .op(n14851) );
  xor2_1 U13983 ( .ip1(n14889), .ip2(n14851), .op(n14906) );
  nor2_1 U13984 ( .ip1(n14853), .ip2(n14852), .op(n14856) );
  nand2_1 U13985 ( .ip1(m1Inputs[157]), .ip2(\STAGE_1/weightReg [7]), .op(
        n14854) );
  fulladder U13986 ( .a(n14856), .b(n14855), .ci(n14854), .co(n14905), .s(
        n14920) );
  fulladder U13987 ( .a(n14859), .b(n14858), .ci(n14857), .co(n14895), .s(
        n14919) );
  fulladder U13988 ( .a(n14862), .b(n14861), .ci(n14860), .co(n14918), .s(
        n14744) );
  inv_1 U13989 ( .ip(n14863), .op(n14915) );
  fulladder U13990 ( .a(n14866), .b(n14865), .ci(n14864), .co(n14909), .s(
        n14867) );
  inv_1 U13991 ( .ip(n14867), .op(n14932) );
  fulladder U13992 ( .a(n14870), .b(n14869), .ci(n14868), .co(n14931), .s(
        n14787) );
  fulladder U13993 ( .a(n14873), .b(n14872), .ci(n14871), .co(n14930), .s(
        n14775) );
  inv_1 U13994 ( .ip(n14874), .op(n14989) );
  nand4_1 U13995 ( .ip1(\STAGE_1/weightReg [11]), .ip2(\STAGE_1/weightReg [10]), .ip3(m1Inputs[156]), .ip4(m1Inputs[155]), .op(n15044) );
  inv_1 U13996 ( .ip(n15044), .op(n14877) );
  or2_1 U13997 ( .ip1(n14875), .ip2(n14877), .op(n14880) );
  nand2_1 U13998 ( .ip1(n14876), .ip2(m1Inputs[156]), .op(n14878) );
  or2_1 U13999 ( .ip1(n14878), .ip2(n14877), .op(n14879) );
  nand2_1 U14000 ( .ip1(n14880), .ip2(n14879), .op(n15041) );
  nand2_1 U14001 ( .ip1(column[158]), .ip2(n14768), .op(n14881) );
  xor2_1 U14002 ( .ip1(n15041), .ip2(n14881), .op(n15020) );
  nor2_1 U14003 ( .ip1(n14883), .ip2(n14882), .op(n14999) );
  nor2_1 U14004 ( .ip1(n12083), .ip2(n14884), .op(n14998) );
  nand2_1 U14005 ( .ip1(m1Inputs[159]), .ip2(\STAGE_1/weightReg [7]), .op(
        n14997) );
  inv_1 U14006 ( .ip(n14885), .op(n15019) );
  fulladder U14007 ( .a(n14888), .b(n14887), .ci(n14886), .co(n15018), .s(
        n14896) );
  and3_1 U14008 ( .ip1(column[157]), .ip2(n14768), .ip3(n14889), .op(n14890)
         );
  nor2_1 U14009 ( .ip1(n14891), .ip2(n14890), .op(n15001) );
  fulladder U14010 ( .a(n14894), .b(n14893), .ci(n14892), .co(n15000), .s(
        n14897) );
  fulladder U14011 ( .a(n14897), .b(n14896), .ci(n14895), .co(n15007), .s(
        n14913) );
  fulladder U14012 ( .a(n14900), .b(n14899), .ci(n14898), .co(n15012), .s(
        n14910) );
  nor2_1 U14013 ( .ip1(n14902), .ip2(n14901), .op(n15017) );
  nor2_1 U14014 ( .ip1(n6503), .ip2(n14903), .op(n15016) );
  nand2_1 U14015 ( .ip1(n14976), .ip2(m1Inputs[151]), .op(n15015) );
  inv_1 U14016 ( .ip(n14904), .op(n15011) );
  fulladder U14017 ( .a(n14907), .b(n14906), .ci(n14905), .co(n15010), .s(
        n14912) );
  fulladder U14018 ( .a(n14910), .b(n14909), .ci(n14908), .co(n14979), .s(
        n14834) );
  fulladder U14019 ( .a(n14913), .b(n14912), .ci(n14911), .co(n14987), .s(
        n14863) );
  fulladder U14020 ( .a(n14916), .b(n14915), .ci(n14914), .co(n14874), .s(
        n14917) );
  inv_1 U14021 ( .ip(n14917), .op(n14943) );
  fulladder U14022 ( .a(n14920), .b(n14919), .ci(n14918), .co(n14911), .s(
        n14921) );
  inv_1 U14023 ( .ip(n14921), .op(n14946) );
  fulladder U14024 ( .a(n14924), .b(n14923), .ci(n14922), .co(n14908), .s(
        n14925) );
  inv_1 U14025 ( .ip(n14925), .op(n14945) );
  fulladder U14026 ( .a(n14928), .b(n14927), .ci(n14926), .co(n14944), .s(
        n14936) );
  inv_1 U14027 ( .ip(n14929), .op(n14942) );
  fulladder U14028 ( .a(n14932), .b(n14931), .ci(n14930), .co(n14914), .s(
        n14933) );
  inv_1 U14029 ( .ip(n14933), .op(n14949) );
  fulladder U14030 ( .a(n14936), .b(n14935), .ci(n14934), .co(n14937), .s(
        n14758) );
  inv_1 U14031 ( .ip(n14937), .op(n14948) );
  fulladder U14032 ( .a(n14940), .b(n14939), .ci(n14938), .co(n14947), .s(
        n14791) );
  fulladder U14033 ( .a(n14943), .b(n14942), .ci(n14941), .co(n14985), .s(
        n14969) );
  fulladder U14034 ( .a(n14946), .b(n14945), .ci(n14944), .co(n14929), .s(
        n14957) );
  fulladder U14035 ( .a(n14949), .b(n14948), .ci(n14947), .co(n14941), .s(
        n14950) );
  inv_1 U14036 ( .ip(n14950), .op(n14956) );
  fulladder U14037 ( .a(n14953), .b(n14952), .ci(n14951), .co(n14955), .s(
        n14799) );
  inv_1 U14038 ( .ip(n14954), .op(n14968) );
  fulladder U14039 ( .a(n14957), .b(n14956), .ci(n14955), .co(n14954), .s(
        n14958) );
  inv_1 U14040 ( .ip(n14958), .op(n14973) );
  fulladder U14041 ( .a(n14961), .b(n14960), .ci(n14959), .co(n14962), .s(
        \STAGE_1/M10/sum [11]) );
  inv_1 U14042 ( .ip(n14962), .op(n14972) );
  fulladder U14043 ( .a(n14965), .b(n14964), .ci(n14963), .co(n14971), .s(
        n14803) );
  inv_1 U14044 ( .ip(n14966), .op(\STAGE_1/M10/sum [14]) );
  fulladder U14045 ( .a(n14969), .b(n14968), .ci(n14967), .co(n14984), .s(
        n14970) );
  inv_1 U14046 ( .ip(n14970), .op(\STAGE_1/M10/sum [13]) );
  fulladder U14047 ( .a(n14973), .b(n14972), .ci(n14971), .co(n14967), .s(
        n14974) );
  inv_1 U14048 ( .ip(n14974), .op(\STAGE_1/M10/sum [12]) );
  nand2_1 U14049 ( .ip1(m1Inputs[159]), .ip2(n14975), .op(n14978) );
  nand2_1 U14050 ( .ip1(m1Inputs[152]), .ip2(n14976), .op(n14977) );
  xor2_1 U14051 ( .ip1(n14978), .ip2(n14977), .op(n14983) );
  fulladder U14052 ( .a(n14981), .b(n14980), .ci(n14979), .co(n14982), .s(
        n14988) );
  xor2_1 U14053 ( .ip1(n14983), .ip2(n14982), .op(n14993) );
  fulladder U14054 ( .a(n14986), .b(n14985), .ci(n14984), .co(n14991), .s(
        n14966) );
  fulladder U14055 ( .a(n14989), .b(n14988), .ci(n14987), .co(n14990), .s(
        n14986) );
  xor2_1 U14056 ( .ip1(n14991), .ip2(n14990), .op(n14992) );
  xor2_1 U14057 ( .ip1(n14993), .ip2(n14992), .op(n14996) );
  nand2_1 U14058 ( .ip1(m1Inputs[158]), .ip2(n14994), .op(n14995) );
  xor2_1 U14059 ( .ip1(n14996), .ip2(n14995), .op(n15040) );
  fulladder U14060 ( .a(n14999), .b(n14998), .ci(n14997), .co(n15004), .s(
        n14885) );
  fulladder U14061 ( .a(n15002), .b(n15001), .ci(n15000), .co(n15003), .s(
        n15008) );
  xor2_1 U14062 ( .ip1(n15004), .ip2(n15003), .op(n15005) );
  xor2_1 U14063 ( .ip1(n15006), .ip2(n15005), .op(n15036) );
  fulladder U14064 ( .a(n15009), .b(n15008), .ci(n15007), .co(n15014), .s(
        n14981) );
  fulladder U14065 ( .a(n15012), .b(n15011), .ci(n15010), .co(n15013), .s(
        n14980) );
  xor2_1 U14066 ( .ip1(n15014), .ip2(n15013), .op(n15024) );
  fulladder U14067 ( .a(n15017), .b(n15016), .ci(n15015), .co(n15022), .s(
        n14904) );
  fulladder U14068 ( .a(n15020), .b(n15019), .ci(n15018), .co(n15021), .s(
        n15009) );
  xor2_1 U14069 ( .ip1(n15022), .ip2(n15021), .op(n15023) );
  xor2_1 U14070 ( .ip1(n15024), .ip2(n15023), .op(n15034) );
  nand2_1 U14071 ( .ip1(m1Inputs[153]), .ip2(\STAGE_1/weightReg [14]), .op(
        n15027) );
  nand2_1 U14072 ( .ip1(m1Inputs[155]), .ip2(n15025), .op(n15026) );
  xor2_1 U14073 ( .ip1(n15027), .ip2(n15026), .op(n15032) );
  nand2_1 U14074 ( .ip1(m1Inputs[154]), .ip2(n15028), .op(n15030) );
  nand2_1 U14075 ( .ip1(m1Inputs[157]), .ip2(\STAGE_1/weightReg [10]), .op(
        n15029) );
  xor2_1 U14076 ( .ip1(n15030), .ip2(n15029), .op(n15031) );
  xor2_1 U14077 ( .ip1(n15032), .ip2(n15031), .op(n15033) );
  xor2_1 U14078 ( .ip1(n15034), .ip2(n15033), .op(n15035) );
  xor2_1 U14079 ( .ip1(n15036), .ip2(n15035), .op(n15038) );
  nand2_1 U14080 ( .ip1(n15042), .ip2(column[159]), .op(n15037) );
  xor2_1 U14081 ( .ip1(n15038), .ip2(n15037), .op(n15039) );
  xor2_1 U14082 ( .ip1(n15040), .ip2(n15039), .op(n15046) );
  nand3_1 U14083 ( .ip1(column[158]), .ip2(n15042), .ip3(n15041), .op(n15043)
         );
  nand2_1 U14084 ( .ip1(n15044), .ip2(n15043), .op(n15045) );
  xor2_1 U14085 ( .ip1(n15046), .ip2(n15045), .op(\STAGE_1/M10/sum [15]) );
  nand3_1 U14086 ( .ip1(\CNTRL/count_layer1_784Q [0]), .ip2(
        \CNTRL/count_layer1_784Q [1]), .ip3(\CNTRL/count_layer1_784Q [2]), 
        .op(n15066) );
  inv_1 U14087 ( .ip(\CNTRL/count_layer1_784Q [3]), .op(n15065) );
  nor2_1 U14088 ( .ip1(n15066), .ip2(n15065), .op(n15070) );
  nand4_1 U14089 ( .ip1(n15070), .ip2(\CNTRL/count_layer1_784Q [8]), .ip3(
        \CNTRL/count_layer1_784Q [9]), .ip4(n15047), .op(n15150) );
  inv_1 U14090 ( .ip(n15150), .op(n15057) );
  inv_1 U14091 ( .ip(\CNTRL/count_layer1_200Q [2]), .op(n15151) );
  and4_1 U14092 ( .ip1(\CNTRL/count_layer1_200Q [3]), .ip2(
        \CNTRL/count_layer1_200Q [6]), .ip3(\CNTRL/count_layer1_200Q [7]), 
        .ip4(n15151), .op(n15049) );
  nor4_1 U14093 ( .ip1(\CNTRL/count_layer1_200Q [0]), .ip2(
        \CNTRL/count_layer1_200Q [1]), .ip3(\CNTRL/count_layer1_200Q [4]), 
        .ip4(\CNTRL/count_layer1_200Q [5]), .op(n15048) );
  nand2_1 U14094 ( .ip1(n15049), .ip2(n15048), .op(n15060) );
  inv_1 U14095 ( .ip(n15113), .op(n15050) );
  nor3_1 U14096 ( .ip1(n15060), .ip2(n15051), .ip3(n15050), .op(n15056) );
  inv_1 U14097 ( .ip(\CNTRL/count_10_2Q [2]), .op(n15122) );
  inv_1 U14098 ( .ip(\CNTRL/count_10_2Q [1]), .op(n15121) );
  and4_1 U14099 ( .ip1(n15122), .ip2(n15121), .ip3(\CNTRL/count_10_2Q [0]), 
        .ip4(\CNTRL/count_10_2Q [3]), .op(n15119) );
  or2_1 U14100 ( .ip1(n15119), .ip2(n15052), .op(n15054) );
  or2_1 U14101 ( .ip1(n15113), .ip2(n15052), .op(n15053) );
  nand2_1 U14102 ( .ip1(n15054), .ip2(n15053), .op(n15055) );
  or2_1 U14103 ( .ip1(n15056), .ip2(n15055), .op(n15095) );
  not_ab_or_c_or_d U14104 ( .ip1(\CNTRL/currentState [1]), .ip2(n15058), .ip3(
        n15057), .ip4(n15095), .op(n15059) );
  nor2_1 U14105 ( .ip1(reset), .ip2(n15059), .op(n4107) );
  nand3_1 U14106 ( .ip1(n15159), .ip2(n15150), .ip3(n15060), .op(n15080) );
  nor2_1 U14107 ( .ip1(\CNTRL/count_layer1_784Q [0]), .ip2(n15080), .op(
        \CNTRL/N233 ) );
  and2_1 U14108 ( .ip1(\CNTRL/count_layer1_784Q [0]), .ip2(
        \CNTRL/count_layer1_784Q [1]), .op(n15062) );
  nor3_1 U14109 ( .ip1(n15062), .ip2(n15061), .ip3(n15080), .op(\CNTRL/N234 )
         );
  nor2_1 U14110 ( .ip1(n15062), .ip2(\CNTRL/count_layer1_784Q [2]), .op(n15064) );
  inv_1 U14111 ( .ip(n15066), .op(n15063) );
  nor3_1 U14112 ( .ip1(n15064), .ip2(n15063), .ip3(n15080), .op(\CNTRL/N235 )
         );
  not_ab_or_c_or_d U14113 ( .ip1(n15066), .ip2(n15065), .ip3(n15070), .ip4(
        n15080), .op(\CNTRL/N236 ) );
  inv_1 U14114 ( .ip(n15070), .op(n15068) );
  inv_1 U14115 ( .ip(\CNTRL/count_layer1_784Q [4]), .op(n15067) );
  nor2_1 U14116 ( .ip1(n15068), .ip2(n15067), .op(n15069) );
  not_ab_or_c_or_d U14117 ( .ip1(n15068), .ip2(n15067), .ip3(n15069), .ip4(
        n15080), .op(\CNTRL/N237 ) );
  nor2_1 U14118 ( .ip1(\CNTRL/count_layer1_784Q [5]), .ip2(n15069), .op(n15072) );
  nand3_1 U14119 ( .ip1(n15070), .ip2(\CNTRL/count_layer1_784Q [4]), .ip3(
        \CNTRL/count_layer1_784Q [5]), .op(n15073) );
  inv_1 U14120 ( .ip(n15073), .op(n15071) );
  nor3_1 U14121 ( .ip1(n15072), .ip2(n15071), .ip3(n15080), .op(\CNTRL/N238 )
         );
  nor2_1 U14122 ( .ip1(n15074), .ip2(n15073), .op(n15075) );
  not_ab_or_c_or_d U14123 ( .ip1(n15074), .ip2(n15073), .ip3(n15075), .ip4(
        n15080), .op(\CNTRL/N239 ) );
  nor2_1 U14124 ( .ip1(\CNTRL/count_layer1_784Q [7]), .ip2(n15075), .op(n15077) );
  nand2_1 U14125 ( .ip1(\CNTRL/count_layer1_784Q [7]), .ip2(n15075), .op(
        n15078) );
  inv_1 U14126 ( .ip(n15078), .op(n15076) );
  nor3_1 U14127 ( .ip1(n15077), .ip2(n15076), .ip3(n15080), .op(\CNTRL/N240 )
         );
  nor2_1 U14128 ( .ip1(n15079), .ip2(n15078), .op(n15082) );
  not_ab_or_c_or_d U14129 ( .ip1(n15079), .ip2(n15078), .ip3(n15082), .ip4(
        n15080), .op(\CNTRL/N241 ) );
  nor2_1 U14130 ( .ip1(\CNTRL/count_layer1_784Q [9]), .ip2(n15082), .op(n15081) );
  not_ab_or_c_or_d U14131 ( .ip1(\CNTRL/count_layer1_784Q [9]), .ip2(n15082), 
        .ip3(n15081), .ip4(n15080), .op(\CNTRL/N242 ) );
  nand4_1 U14132 ( .ip1(\CNTRL/currentState [1]), .ip2(\CNTRL/currentState [0]), .ip3(\CNTRL/count_20Q [0]), .ip4(n15083), .op(n15084) );
  inv_1 U14133 ( .ip(n15084), .op(n17241) );
  or2_1 U14134 ( .ip1(n17241), .ip2(n17229), .op(n16860) );
  or2_1 U14135 ( .ip1(n15086), .ip2(n15085), .op(n15088) );
  nand2_1 U14136 ( .ip1(n15088), .ip2(n15087), .op(n15188) );
  nand2_1 U14137 ( .ip1(\CNTRL/count_20Q [1]), .ip2(n15188), .op(n15165) );
  nor2_1 U14138 ( .ip1(n15165), .ip2(n15167), .op(n15379) );
  and2_1 U14139 ( .ip1(n16860), .ip2(n15379), .op(weight2_loadNextRow) );
  nor4_1 U14140 ( .ip1(n15110), .ip2(n15174), .ip3(n15100), .ip4(n15098), .op(
        n15090) );
  mux2_1 U14141 ( .ip1(n15090), .ip2(n15089), .s(\CNTRL/count_20Q [4]), .op(
        n4111) );
  nand3_1 U14142 ( .ip1(n15092), .ip2(n15113), .ip3(n15091), .op(n15093) );
  and3_1 U14143 ( .ip1(\CNTRL/currentState [2]), .ip2(n15094), .ip3(n15093), 
        .op(n15096) );
  nor3_1 U14144 ( .ip1(n15096), .ip2(n15095), .ip3(weight2_loadNextRow), .op(
        n15097) );
  nor2_1 U14145 ( .ip1(reset), .ip2(n15097), .op(n4109) );
  inv_1 U14146 ( .ip(n15098), .op(n15103) );
  mux2_1 U14147 ( .ip1(n15103), .ip2(n15099), .s(\CNTRL/count_20Q [0]), .op(
        n4106) );
  nand2_1 U14148 ( .ip1(n15103), .ip2(n15100), .op(n15101) );
  nand2_1 U14149 ( .ip1(n15102), .ip2(n15101), .op(n15112) );
  inv_1 U14150 ( .ip(n15112), .op(n15107) );
  or2_1 U14151 ( .ip1(\CNTRL/count_20Q [0]), .ip2(\CNTRL/count_20Q [1]), .op(
        n15105) );
  or2_1 U14152 ( .ip1(n15103), .ip2(\CNTRL/count_20Q [1]), .op(n15104) );
  nand2_1 U14153 ( .ip1(n15105), .ip2(n15104), .op(n15106) );
  nor2_1 U14154 ( .ip1(n15107), .ip2(n15106), .op(n4105) );
  and2_1 U14155 ( .ip1(n15109), .ip2(n15108), .op(n15111) );
  mux2_1 U14156 ( .ip1(n15112), .ip2(n15111), .s(n15110), .op(n4104) );
  inv_1 U14157 ( .ip(\CNTRL/count_10_2Q [0]), .op(n15115) );
  nand2_1 U14158 ( .ip1(n16714), .ip2(n15113), .op(n15116) );
  nor2_1 U14159 ( .ip1(n15115), .ip2(n15116), .op(n15114) );
  not_ab_or_c_or_d U14160 ( .ip1(n15115), .ip2(n15116), .ip3(reset), .ip4(
        n15114), .op(n4102) );
  nand2_1 U14161 ( .ip1(n15115), .ip2(n15159), .op(n15118) );
  nand2_1 U14162 ( .ip1(n15159), .ip2(n15116), .op(n15117) );
  nand2_1 U14163 ( .ip1(n15118), .ip2(n15117), .op(n15120) );
  nor2_1 U14164 ( .ip1(n15121), .ip2(n15120), .op(n15124) );
  nor2_1 U14165 ( .ip1(reset), .ip2(n15119), .op(n15126) );
  nor2_1 U14166 ( .ip1(n15126), .ip2(n15120), .op(n15129) );
  not_ab_or_c_or_d U14167 ( .ip1(n15121), .ip2(n15120), .ip3(n15124), .ip4(
        n15129), .op(n4101) );
  inv_1 U14168 ( .ip(n15124), .op(n15123) );
  nor2_1 U14169 ( .ip1(n15123), .ip2(n15122), .op(n15130) );
  or2_1 U14170 ( .ip1(n15124), .ip2(\CNTRL/count_10_2Q [2]), .op(n15125) );
  nand2_1 U14171 ( .ip1(n15126), .ip2(n15125), .op(n15127) );
  nor2_1 U14172 ( .ip1(n15130), .ip2(n15127), .op(n4100) );
  nor2_1 U14173 ( .ip1(\CNTRL/count_10_2Q [3]), .ip2(n15130), .op(n15128) );
  not_ab_or_c_or_d U14174 ( .ip1(\CNTRL/count_10_2Q [3]), .ip2(n15130), .ip3(
        n15129), .ip4(n15128), .op(n4099) );
  inv_1 U14175 ( .ip(n15131), .op(n15141) );
  nor2_1 U14176 ( .ip1(n15132), .ip2(n15141), .op(n15134) );
  mux2_1 U14177 ( .ip1(n15134), .ip2(n15133), .s(\CNTRL/count_10Q [1]), .op(
        n4097) );
  nor2_1 U14178 ( .ip1(n15140), .ip2(n15136), .op(n15138) );
  nand2_1 U14179 ( .ip1(\CNTRL/count_10Q [0]), .ip2(\CNTRL/count_10Q [1]), 
        .op(n15135) );
  and3_1 U14180 ( .ip1(\CNTRL/count_10Q [0]), .ip2(\CNTRL/count_10Q [1]), 
        .ip3(\CNTRL/count_10Q [2]), .op(n15143) );
  not_ab_or_c_or_d U14181 ( .ip1(n15136), .ip2(n15135), .ip3(n15143), .ip4(
        n15141), .op(n15137) );
  or2_1 U14182 ( .ip1(n15138), .ip2(n15137), .op(n4096) );
  nor2_1 U14183 ( .ip1(n15140), .ip2(n15139), .op(n15145) );
  nor2_1 U14184 ( .ip1(\CNTRL/count_10Q [3]), .ip2(n15143), .op(n15142) );
  not_ab_or_c_or_d U14185 ( .ip1(\CNTRL/count_10Q [3]), .ip2(n15143), .ip3(
        n15142), .ip4(n15141), .op(n15144) );
  or2_1 U14186 ( .ip1(n15145), .ip2(n15144), .op(n4095) );
  inv_1 U14187 ( .ip(\CNTRL/count_layer1_200Q [0]), .op(n15149) );
  nor2_1 U14188 ( .ip1(n15150), .ip2(n15149), .op(n15148) );
  nor2_1 U14189 ( .ip1(n15148), .ip2(\CNTRL/count_layer1_200Q [1]), .op(n15147) );
  nand2_1 U14190 ( .ip1(n15148), .ip2(\CNTRL/count_layer1_200Q [1]), .op(
        n15152) );
  inv_1 U14191 ( .ip(n15152), .op(n15146) );
  nor3_1 U14192 ( .ip1(n15147), .ip2(reset), .ip3(n15146), .op(n4094) );
  not_ab_or_c_or_d U14193 ( .ip1(n15150), .ip2(n15149), .ip3(reset), .ip4(
        n15148), .op(n4093) );
  nor2_1 U14194 ( .ip1(n15152), .ip2(n15151), .op(n15153) );
  not_ab_or_c_or_d U14195 ( .ip1(n15152), .ip2(n15151), .ip3(reset), .ip4(
        n15153), .op(n4092) );
  nor2_1 U14196 ( .ip1(n15153), .ip2(\CNTRL/count_layer1_200Q [3]), .op(n15155) );
  nand2_1 U14197 ( .ip1(n15153), .ip2(\CNTRL/count_layer1_200Q [3]), .op(
        n15157) );
  inv_1 U14198 ( .ip(n15157), .op(n15154) );
  nor3_1 U14199 ( .ip1(n15155), .ip2(reset), .ip3(n15154), .op(n4091) );
  inv_1 U14200 ( .ip(\CNTRL/count_layer1_200Q [4]), .op(n15156) );
  nor2_1 U14201 ( .ip1(n15157), .ip2(n15156), .op(n15160) );
  not_ab_or_c_or_d U14202 ( .ip1(n15157), .ip2(n15156), .ip3(reset), .ip4(
        n15160), .op(n4090) );
  nor2_1 U14203 ( .ip1(n15160), .ip2(\CNTRL/count_layer1_200Q [5]), .op(n15158) );
  not_ab_or_c_or_d U14204 ( .ip1(n15160), .ip2(\CNTRL/count_layer1_200Q [5]), 
        .ip3(reset), .ip4(n15158), .op(n4089) );
  nand3_1 U14205 ( .ip1(n15160), .ip2(\CNTRL/count_layer1_200Q [5]), .ip3(
        n15159), .op(n15162) );
  inv_1 U14206 ( .ip(\CNTRL/count_layer1_200Q [6]), .op(n15161) );
  nor2_1 U14207 ( .ip1(n15162), .ip2(n15161), .op(n15164) );
  not_ab_or_c_or_d U14208 ( .ip1(n15162), .ip2(n15161), .ip3(reset), .ip4(
        n15164), .op(n4088) );
  nor2_1 U14209 ( .ip1(n15164), .ip2(reset), .op(n15163) );
  mux2_1 U14210 ( .ip1(n15164), .ip2(n15163), .s(\CNTRL/count_layer1_200Q [7]), 
        .op(n4087) );
  inv_1 U14211 ( .ip(n15165), .op(n15172) );
  nand2_1 U14212 ( .ip1(n15172), .ip2(n15184), .op(n15177) );
  nand3_1 U14213 ( .ip1(\CNTRL/count_20Q [2]), .ip2(\CNTRL/count_20Q [3]), 
        .ip3(n15188), .op(n15173) );
  nor2_1 U14214 ( .ip1(n15177), .ip2(n15173), .op(n16855) );
  nand2_1 U14215 ( .ip1(n16855), .ip2(\ROUTEDATA/regData [112]), .op(n15191)
         );
  nor4_1 U14216 ( .ip1(\CNTRL/count_20Q [2]), .ip2(\CNTRL/count_20Q [4]), 
        .ip3(n15174), .ip4(n15165), .op(n16847) );
  nand2_1 U14217 ( .ip1(n15188), .ip2(n15186), .op(n15166) );
  nor4_1 U14218 ( .ip1(\CNTRL/count_20Q [2]), .ip2(\CNTRL/count_20Q [4]), 
        .ip3(n15174), .ip4(n15166), .op(n16843) );
  nand2_1 U14219 ( .ip1(n16843), .ip2(\ROUTEDATA/regData [64]), .op(n15170) );
  inv_1 U14220 ( .ip(n15188), .op(n15171) );
  nor3_1 U14221 ( .ip1(\CNTRL/count_20Q [1]), .ip2(n15171), .ip3(n15167), .op(
        n16859) );
  nand2_1 U14222 ( .ip1(n16859), .ip2(\ROUTEDATA/regData [128]), .op(n15169)
         );
  nand2_1 U14223 ( .ip1(n15379), .ip2(\ROUTEDATA/regData [144]), .op(n15168)
         );
  nand3_1 U14224 ( .ip1(n15170), .ip2(n15169), .ip3(n15168), .op(n15183) );
  nor2_1 U14225 ( .ip1(n15184), .ip2(n15171), .op(n15192) );
  or2_1 U14226 ( .ip1(n15192), .ip2(n15172), .op(n15176) );
  nor2_1 U14227 ( .ip1(n15173), .ip2(n15176), .op(n16851) );
  nand2_1 U14228 ( .ip1(n16851), .ip2(\ROUTEDATA/regData [96]), .op(n15181) );
  nand3_1 U14229 ( .ip1(\CNTRL/count_20Q [2]), .ip2(n15188), .ip3(n15174), 
        .op(n15175) );
  nor2_1 U14230 ( .ip1(n15177), .ip2(n15175), .op(n16839) );
  nand2_1 U14231 ( .ip1(n16839), .ip2(\ROUTEDATA/regData [48]), .op(n15180) );
  nor2_1 U14232 ( .ip1(n15176), .ip2(n15175), .op(n16835) );
  nand2_1 U14233 ( .ip1(n16835), .ip2(\ROUTEDATA/regData [32]), .op(n15179) );
  inv_1 U14234 ( .ip(n15185), .op(n15193) );
  nor2_1 U14235 ( .ip1(n15193), .ip2(n15177), .op(n16831) );
  nand2_1 U14236 ( .ip1(n16831), .ip2(\ROUTEDATA/regData [16]), .op(n15178) );
  nand4_1 U14237 ( .ip1(n15181), .ip2(n15180), .ip3(n15179), .ip4(n15178), 
        .op(n15182) );
  not_ab_or_c_or_d U14238 ( .ip1(n16847), .ip2(\ROUTEDATA/regData [80]), .ip3(
        n15183), .ip4(n15182), .op(n15190) );
  nand3_1 U14239 ( .ip1(n15186), .ip2(n15185), .ip3(n15184), .op(n15187) );
  nand2_1 U14240 ( .ip1(n15188), .ip2(n15187), .op(n17243) );
  nand2_1 U14241 ( .ip1(n17243), .ip2(\ROUTEDATA/regData [0]), .op(n15189) );
  nand3_1 U14242 ( .ip1(n15191), .ip2(n15190), .ip3(n15189), .op(n15196) );
  or2_1 U14243 ( .ip1(n15192), .ip2(n16860), .op(n15195) );
  or2_1 U14244 ( .ip1(n15193), .ip2(n16860), .op(n15194) );
  nand2_1 U14245 ( .ip1(n15195), .ip2(n15194), .op(n15392) );
  mux2_1 U14246 ( .ip1(m2DataIn[0]), .ip2(n15196), .s(n15392), .op(n4086) );
  nand2_1 U14247 ( .ip1(\ROUTEDATA/regData [97]), .ip2(n16851), .op(n15208) );
  nand2_1 U14248 ( .ip1(\ROUTEDATA/regData [65]), .ip2(n16843), .op(n15199) );
  nand2_1 U14249 ( .ip1(n15379), .ip2(\ROUTEDATA/regData [145]), .op(n15198)
         );
  nand2_1 U14250 ( .ip1(n16859), .ip2(\ROUTEDATA/regData [129]), .op(n15197)
         );
  nand3_1 U14251 ( .ip1(n15199), .ip2(n15198), .ip3(n15197), .op(n15205) );
  nand2_1 U14252 ( .ip1(n16839), .ip2(\ROUTEDATA/regData [49]), .op(n15203) );
  nand2_1 U14253 ( .ip1(n17243), .ip2(\ROUTEDATA/regData [1]), .op(n15202) );
  nand2_1 U14254 ( .ip1(n16835), .ip2(\ROUTEDATA/regData [33]), .op(n15201) );
  nand2_1 U14255 ( .ip1(n16855), .ip2(\ROUTEDATA/regData [113]), .op(n15200)
         );
  nand4_1 U14256 ( .ip1(n15203), .ip2(n15202), .ip3(n15201), .ip4(n15200), 
        .op(n15204) );
  not_ab_or_c_or_d U14257 ( .ip1(n16847), .ip2(\ROUTEDATA/regData [81]), .ip3(
        n15205), .ip4(n15204), .op(n15207) );
  nand2_1 U14258 ( .ip1(n16831), .ip2(\ROUTEDATA/regData [17]), .op(n15206) );
  nand3_1 U14259 ( .ip1(n15208), .ip2(n15207), .ip3(n15206), .op(n15209) );
  mux2_1 U14260 ( .ip1(m2DataIn[1]), .ip2(n15209), .s(n15392), .op(n4085) );
  nand2_1 U14261 ( .ip1(n16839), .ip2(\ROUTEDATA/regData [50]), .op(n15221) );
  nand2_1 U14262 ( .ip1(n16843), .ip2(\ROUTEDATA/regData [66]), .op(n15212) );
  nand2_1 U14263 ( .ip1(n15379), .ip2(\ROUTEDATA/regData [146]), .op(n15211)
         );
  nand2_1 U14264 ( .ip1(n16859), .ip2(\ROUTEDATA/regData [130]), .op(n15210)
         );
  nand3_1 U14265 ( .ip1(n15212), .ip2(n15211), .ip3(n15210), .op(n15218) );
  nand2_1 U14266 ( .ip1(n16831), .ip2(\ROUTEDATA/regData [18]), .op(n15216) );
  nand2_1 U14267 ( .ip1(n16851), .ip2(\ROUTEDATA/regData [98]), .op(n15215) );
  nand2_1 U14268 ( .ip1(n17243), .ip2(\ROUTEDATA/regData [2]), .op(n15214) );
  nand2_1 U14269 ( .ip1(n16855), .ip2(\ROUTEDATA/regData [114]), .op(n15213)
         );
  nand4_1 U14270 ( .ip1(n15216), .ip2(n15215), .ip3(n15214), .ip4(n15213), 
        .op(n15217) );
  not_ab_or_c_or_d U14271 ( .ip1(n16847), .ip2(\ROUTEDATA/regData [82]), .ip3(
        n15218), .ip4(n15217), .op(n15220) );
  nand2_1 U14272 ( .ip1(n16835), .ip2(\ROUTEDATA/regData [34]), .op(n15219) );
  nand3_1 U14273 ( .ip1(n15221), .ip2(n15220), .ip3(n15219), .op(n15222) );
  mux2_1 U14274 ( .ip1(m2DataIn[2]), .ip2(n15222), .s(n15392), .op(n4084) );
  nand2_1 U14275 ( .ip1(n16855), .ip2(\ROUTEDATA/regData [115]), .op(n15234)
         );
  nand2_1 U14276 ( .ip1(n16843), .ip2(\ROUTEDATA/regData [67]), .op(n15225) );
  nand2_1 U14277 ( .ip1(n16859), .ip2(\ROUTEDATA/regData [131]), .op(n15224)
         );
  nand2_1 U14278 ( .ip1(n15379), .ip2(\ROUTEDATA/regData [147]), .op(n15223)
         );
  nand3_1 U14279 ( .ip1(n15225), .ip2(n15224), .ip3(n15223), .op(n15231) );
  nand2_1 U14280 ( .ip1(n16839), .ip2(\ROUTEDATA/regData [51]), .op(n15229) );
  nand2_1 U14281 ( .ip1(n16831), .ip2(\ROUTEDATA/regData [19]), .op(n15228) );
  nand2_1 U14282 ( .ip1(n16851), .ip2(\ROUTEDATA/regData [99]), .op(n15227) );
  nand2_1 U14283 ( .ip1(n17243), .ip2(\ROUTEDATA/regData [3]), .op(n15226) );
  nand4_1 U14284 ( .ip1(n15229), .ip2(n15228), .ip3(n15227), .ip4(n15226), 
        .op(n15230) );
  not_ab_or_c_or_d U14285 ( .ip1(n16847), .ip2(\ROUTEDATA/regData [83]), .ip3(
        n15231), .ip4(n15230), .op(n15233) );
  nand2_1 U14286 ( .ip1(n16835), .ip2(\ROUTEDATA/regData [35]), .op(n15232) );
  nand3_1 U14287 ( .ip1(n15234), .ip2(n15233), .ip3(n15232), .op(n15235) );
  mux2_1 U14288 ( .ip1(m2DataIn[3]), .ip2(n15235), .s(n15392), .op(n4083) );
  nand2_1 U14289 ( .ip1(n16855), .ip2(\ROUTEDATA/regData [116]), .op(n15247)
         );
  nand2_1 U14290 ( .ip1(\ROUTEDATA/regData [68]), .ip2(n16843), .op(n15238) );
  nand2_1 U14291 ( .ip1(n15379), .ip2(\ROUTEDATA/regData [148]), .op(n15237)
         );
  nand2_1 U14292 ( .ip1(n16859), .ip2(\ROUTEDATA/regData [132]), .op(n15236)
         );
  nand3_1 U14293 ( .ip1(n15238), .ip2(n15237), .ip3(n15236), .op(n15244) );
  nand2_1 U14294 ( .ip1(n17243), .ip2(\ROUTEDATA/regData [4]), .op(n15242) );
  nand2_1 U14295 ( .ip1(n16839), .ip2(\ROUTEDATA/regData [52]), .op(n15241) );
  nand2_1 U14296 ( .ip1(n16831), .ip2(\ROUTEDATA/regData [20]), .op(n15240) );
  nand2_1 U14297 ( .ip1(n16835), .ip2(\ROUTEDATA/regData [36]), .op(n15239) );
  nand4_1 U14298 ( .ip1(n15242), .ip2(n15241), .ip3(n15240), .ip4(n15239), 
        .op(n15243) );
  not_ab_or_c_or_d U14299 ( .ip1(n16847), .ip2(\ROUTEDATA/regData [84]), .ip3(
        n15244), .ip4(n15243), .op(n15246) );
  nand2_1 U14300 ( .ip1(n16851), .ip2(\ROUTEDATA/regData [100]), .op(n15245)
         );
  nand3_1 U14301 ( .ip1(n15247), .ip2(n15246), .ip3(n15245), .op(n15248) );
  mux2_1 U14302 ( .ip1(m2DataIn[4]), .ip2(n15248), .s(n15392), .op(n4082) );
  nand2_1 U14303 ( .ip1(n16855), .ip2(\ROUTEDATA/regData [117]), .op(n15260)
         );
  nand2_1 U14304 ( .ip1(n16843), .ip2(\ROUTEDATA/regData [69]), .op(n15251) );
  nand2_1 U14305 ( .ip1(n16859), .ip2(\ROUTEDATA/regData [133]), .op(n15250)
         );
  nand2_1 U14306 ( .ip1(n15379), .ip2(\ROUTEDATA/regData [149]), .op(n15249)
         );
  nand3_1 U14307 ( .ip1(n15251), .ip2(n15250), .ip3(n15249), .op(n15257) );
  nand2_1 U14308 ( .ip1(n16835), .ip2(\ROUTEDATA/regData [37]), .op(n15255) );
  nand2_1 U14309 ( .ip1(n16831), .ip2(\ROUTEDATA/regData [21]), .op(n15254) );
  nand2_1 U14310 ( .ip1(n16839), .ip2(\ROUTEDATA/regData [53]), .op(n15253) );
  nand2_1 U14311 ( .ip1(n16851), .ip2(\ROUTEDATA/regData [101]), .op(n15252)
         );
  nand4_1 U14312 ( .ip1(n15255), .ip2(n15254), .ip3(n15253), .ip4(n15252), 
        .op(n15256) );
  not_ab_or_c_or_d U14313 ( .ip1(n16847), .ip2(\ROUTEDATA/regData [85]), .ip3(
        n15257), .ip4(n15256), .op(n15259) );
  nand2_1 U14314 ( .ip1(n17243), .ip2(\ROUTEDATA/regData [5]), .op(n15258) );
  nand3_1 U14315 ( .ip1(n15260), .ip2(n15259), .ip3(n15258), .op(n15261) );
  mux2_1 U14316 ( .ip1(m2DataIn[5]), .ip2(n15261), .s(n15392), .op(n4081) );
  nand2_1 U14317 ( .ip1(\ROUTEDATA/regData [6]), .ip2(n17243), .op(n15273) );
  nand2_1 U14318 ( .ip1(\ROUTEDATA/regData [70]), .ip2(n16843), .op(n15264) );
  nand2_1 U14319 ( .ip1(n16859), .ip2(\ROUTEDATA/regData [134]), .op(n15263)
         );
  nand2_1 U14320 ( .ip1(n15379), .ip2(\ROUTEDATA/regData [150]), .op(n15262)
         );
  nand3_1 U14321 ( .ip1(n15264), .ip2(n15263), .ip3(n15262), .op(n15270) );
  nand2_1 U14322 ( .ip1(n16851), .ip2(\ROUTEDATA/regData [102]), .op(n15268)
         );
  nand2_1 U14323 ( .ip1(n16855), .ip2(\ROUTEDATA/regData [118]), .op(n15267)
         );
  nand2_1 U14324 ( .ip1(n16831), .ip2(\ROUTEDATA/regData [22]), .op(n15266) );
  nand2_1 U14325 ( .ip1(n16835), .ip2(\ROUTEDATA/regData [38]), .op(n15265) );
  nand4_1 U14326 ( .ip1(n15268), .ip2(n15267), .ip3(n15266), .ip4(n15265), 
        .op(n15269) );
  not_ab_or_c_or_d U14327 ( .ip1(n16847), .ip2(\ROUTEDATA/regData [86]), .ip3(
        n15270), .ip4(n15269), .op(n15272) );
  nand2_1 U14328 ( .ip1(n16839), .ip2(\ROUTEDATA/regData [54]), .op(n15271) );
  nand3_1 U14329 ( .ip1(n15273), .ip2(n15272), .ip3(n15271), .op(n15274) );
  mux2_1 U14330 ( .ip1(m2DataIn[6]), .ip2(n15274), .s(n15392), .op(n4080) );
  nand2_1 U14331 ( .ip1(\ROUTEDATA/regData [55]), .ip2(n16839), .op(n15286) );
  nand2_1 U14332 ( .ip1(n16843), .ip2(\ROUTEDATA/regData [71]), .op(n15277) );
  nand2_1 U14333 ( .ip1(n16859), .ip2(\ROUTEDATA/regData [135]), .op(n15276)
         );
  nand2_1 U14334 ( .ip1(n15379), .ip2(\ROUTEDATA/regData [151]), .op(n15275)
         );
  nand3_1 U14335 ( .ip1(n15277), .ip2(n15276), .ip3(n15275), .op(n15283) );
  nand2_1 U14336 ( .ip1(n16851), .ip2(\ROUTEDATA/regData [103]), .op(n15281)
         );
  nand2_1 U14337 ( .ip1(n17243), .ip2(\ROUTEDATA/regData [7]), .op(n15280) );
  nand2_1 U14338 ( .ip1(n16855), .ip2(\ROUTEDATA/regData [119]), .op(n15279)
         );
  nand2_1 U14339 ( .ip1(n16835), .ip2(\ROUTEDATA/regData [39]), .op(n15278) );
  nand4_1 U14340 ( .ip1(n15281), .ip2(n15280), .ip3(n15279), .ip4(n15278), 
        .op(n15282) );
  not_ab_or_c_or_d U14341 ( .ip1(n16847), .ip2(\ROUTEDATA/regData [87]), .ip3(
        n15283), .ip4(n15282), .op(n15285) );
  nand2_1 U14342 ( .ip1(n16831), .ip2(\ROUTEDATA/regData [23]), .op(n15284) );
  nand3_1 U14343 ( .ip1(n15286), .ip2(n15285), .ip3(n15284), .op(n15287) );
  mux2_1 U14344 ( .ip1(m2DataIn[7]), .ip2(n15287), .s(n15392), .op(n4079) );
  nand2_1 U14345 ( .ip1(n16855), .ip2(\ROUTEDATA/regData [120]), .op(n15299)
         );
  nand2_1 U14346 ( .ip1(n16843), .ip2(\ROUTEDATA/regData [72]), .op(n15290) );
  nand2_1 U14347 ( .ip1(n15379), .ip2(\ROUTEDATA/regData [152]), .op(n15289)
         );
  nand2_1 U14348 ( .ip1(n16859), .ip2(\ROUTEDATA/regData [136]), .op(n15288)
         );
  nand3_1 U14349 ( .ip1(n15290), .ip2(n15289), .ip3(n15288), .op(n15296) );
  nand2_1 U14350 ( .ip1(n16839), .ip2(\ROUTEDATA/regData [56]), .op(n15294) );
  nand2_1 U14351 ( .ip1(n16835), .ip2(\ROUTEDATA/regData [40]), .op(n15293) );
  nand2_1 U14352 ( .ip1(n16831), .ip2(\ROUTEDATA/regData [24]), .op(n15292) );
  nand2_1 U14353 ( .ip1(n17243), .ip2(\ROUTEDATA/regData [8]), .op(n15291) );
  nand4_1 U14354 ( .ip1(n15294), .ip2(n15293), .ip3(n15292), .ip4(n15291), 
        .op(n15295) );
  not_ab_or_c_or_d U14355 ( .ip1(n16847), .ip2(\ROUTEDATA/regData [88]), .ip3(
        n15296), .ip4(n15295), .op(n15298) );
  nand2_1 U14356 ( .ip1(n16851), .ip2(\ROUTEDATA/regData [104]), .op(n15297)
         );
  nand3_1 U14357 ( .ip1(n15299), .ip2(n15298), .ip3(n15297), .op(n15300) );
  mux2_1 U14358 ( .ip1(m2DataIn[8]), .ip2(n15300), .s(n15392), .op(n4078) );
  nand2_1 U14359 ( .ip1(n16855), .ip2(\ROUTEDATA/regData [121]), .op(n15312)
         );
  nand2_1 U14360 ( .ip1(\ROUTEDATA/regData [73]), .ip2(n16843), .op(n15303) );
  nand2_1 U14361 ( .ip1(n16859), .ip2(\ROUTEDATA/regData [137]), .op(n15302)
         );
  nand2_1 U14362 ( .ip1(n15379), .ip2(\ROUTEDATA/regData [153]), .op(n15301)
         );
  nand3_1 U14363 ( .ip1(n15303), .ip2(n15302), .ip3(n15301), .op(n15309) );
  nand2_1 U14364 ( .ip1(n16831), .ip2(\ROUTEDATA/regData [25]), .op(n15307) );
  nand2_1 U14365 ( .ip1(n16851), .ip2(\ROUTEDATA/regData [105]), .op(n15306)
         );
  nand2_1 U14366 ( .ip1(n16835), .ip2(\ROUTEDATA/regData [41]), .op(n15305) );
  nand2_1 U14367 ( .ip1(n16839), .ip2(\ROUTEDATA/regData [57]), .op(n15304) );
  nand4_1 U14368 ( .ip1(n15307), .ip2(n15306), .ip3(n15305), .ip4(n15304), 
        .op(n15308) );
  not_ab_or_c_or_d U14369 ( .ip1(n16847), .ip2(\ROUTEDATA/regData [89]), .ip3(
        n15309), .ip4(n15308), .op(n15311) );
  nand2_1 U14370 ( .ip1(n17243), .ip2(\ROUTEDATA/regData [9]), .op(n15310) );
  nand3_1 U14371 ( .ip1(n15312), .ip2(n15311), .ip3(n15310), .op(n15313) );
  mux2_1 U14372 ( .ip1(m2DataIn[9]), .ip2(n15313), .s(n15392), .op(n4077) );
  nand2_1 U14373 ( .ip1(n16855), .ip2(\ROUTEDATA/regData [122]), .op(n15325)
         );
  nand2_1 U14374 ( .ip1(\ROUTEDATA/regData [74]), .ip2(n16843), .op(n15316) );
  nand2_1 U14375 ( .ip1(n15379), .ip2(\ROUTEDATA/regData [154]), .op(n15315)
         );
  nand2_1 U14376 ( .ip1(n16859), .ip2(\ROUTEDATA/regData [138]), .op(n15314)
         );
  nand3_1 U14377 ( .ip1(n15316), .ip2(n15315), .ip3(n15314), .op(n15322) );
  nand2_1 U14378 ( .ip1(n16831), .ip2(\ROUTEDATA/regData [26]), .op(n15320) );
  nand2_1 U14379 ( .ip1(n16835), .ip2(\ROUTEDATA/regData [42]), .op(n15319) );
  nand2_1 U14380 ( .ip1(n17243), .ip2(\ROUTEDATA/regData [10]), .op(n15318) );
  nand2_1 U14381 ( .ip1(n16851), .ip2(\ROUTEDATA/regData [106]), .op(n15317)
         );
  nand4_1 U14382 ( .ip1(n15320), .ip2(n15319), .ip3(n15318), .ip4(n15317), 
        .op(n15321) );
  not_ab_or_c_or_d U14383 ( .ip1(n16847), .ip2(\ROUTEDATA/regData [90]), .ip3(
        n15322), .ip4(n15321), .op(n15324) );
  nand2_1 U14384 ( .ip1(n16839), .ip2(\ROUTEDATA/regData [58]), .op(n15323) );
  nand3_1 U14385 ( .ip1(n15325), .ip2(n15324), .ip3(n15323), .op(n15326) );
  mux2_1 U14386 ( .ip1(m2DataIn[10]), .ip2(n15326), .s(n15392), .op(n4076) );
  nand2_1 U14387 ( .ip1(n16839), .ip2(\ROUTEDATA/regData [59]), .op(n15338) );
  nand2_1 U14388 ( .ip1(\ROUTEDATA/regData [75]), .ip2(n16843), .op(n15329) );
  nand2_1 U14389 ( .ip1(n15379), .ip2(\ROUTEDATA/regData [155]), .op(n15328)
         );
  nand2_1 U14390 ( .ip1(n16859), .ip2(\ROUTEDATA/regData [139]), .op(n15327)
         );
  nand3_1 U14391 ( .ip1(n15329), .ip2(n15328), .ip3(n15327), .op(n15335) );
  nand2_1 U14392 ( .ip1(n17243), .ip2(\ROUTEDATA/regData [11]), .op(n15333) );
  nand2_1 U14393 ( .ip1(n16831), .ip2(\ROUTEDATA/regData [27]), .op(n15332) );
  nand2_1 U14394 ( .ip1(n16855), .ip2(\ROUTEDATA/regData [123]), .op(n15331)
         );
  nand2_1 U14395 ( .ip1(n16851), .ip2(\ROUTEDATA/regData [107]), .op(n15330)
         );
  nand4_1 U14396 ( .ip1(n15333), .ip2(n15332), .ip3(n15331), .ip4(n15330), 
        .op(n15334) );
  not_ab_or_c_or_d U14397 ( .ip1(n16847), .ip2(\ROUTEDATA/regData [91]), .ip3(
        n15335), .ip4(n15334), .op(n15337) );
  nand2_1 U14398 ( .ip1(n16835), .ip2(\ROUTEDATA/regData [43]), .op(n15336) );
  nand3_1 U14399 ( .ip1(n15338), .ip2(n15337), .ip3(n15336), .op(n15339) );
  mux2_1 U14400 ( .ip1(m2DataIn[11]), .ip2(n15339), .s(n15392), .op(n4075) );
  nand2_1 U14401 ( .ip1(\ROUTEDATA/regData [12]), .ip2(n17243), .op(n15351) );
  nand2_1 U14402 ( .ip1(\ROUTEDATA/regData [76]), .ip2(n16843), .op(n15342) );
  nand2_1 U14403 ( .ip1(n16859), .ip2(\ROUTEDATA/regData [140]), .op(n15341)
         );
  nand2_1 U14404 ( .ip1(n15379), .ip2(\ROUTEDATA/regData [156]), .op(n15340)
         );
  nand3_1 U14405 ( .ip1(n15342), .ip2(n15341), .ip3(n15340), .op(n15348) );
  nand2_1 U14406 ( .ip1(n16855), .ip2(\ROUTEDATA/regData [124]), .op(n15346)
         );
  nand2_1 U14407 ( .ip1(n16839), .ip2(\ROUTEDATA/regData [60]), .op(n15345) );
  nand2_1 U14408 ( .ip1(n16831), .ip2(\ROUTEDATA/regData [28]), .op(n15344) );
  nand2_1 U14409 ( .ip1(n16835), .ip2(\ROUTEDATA/regData [44]), .op(n15343) );
  nand4_1 U14410 ( .ip1(n15346), .ip2(n15345), .ip3(n15344), .ip4(n15343), 
        .op(n15347) );
  not_ab_or_c_or_d U14411 ( .ip1(n16847), .ip2(\ROUTEDATA/regData [92]), .ip3(
        n15348), .ip4(n15347), .op(n15350) );
  nand2_1 U14412 ( .ip1(n16851), .ip2(\ROUTEDATA/regData [108]), .op(n15349)
         );
  nand3_1 U14413 ( .ip1(n15351), .ip2(n15350), .ip3(n15349), .op(n15352) );
  mux2_1 U14414 ( .ip1(m2DataIn[12]), .ip2(n15352), .s(n15392), .op(n4074) );
  nand2_1 U14415 ( .ip1(n17243), .ip2(\ROUTEDATA/regData [13]), .op(n15364) );
  nand2_1 U14416 ( .ip1(n16843), .ip2(\ROUTEDATA/regData [77]), .op(n15355) );
  nand2_1 U14417 ( .ip1(n15379), .ip2(\ROUTEDATA/regData [157]), .op(n15354)
         );
  nand2_1 U14418 ( .ip1(n16859), .ip2(\ROUTEDATA/regData [141]), .op(n15353)
         );
  nand3_1 U14419 ( .ip1(n15355), .ip2(n15354), .ip3(n15353), .op(n15361) );
  nand2_1 U14420 ( .ip1(n16831), .ip2(\ROUTEDATA/regData [29]), .op(n15359) );
  nand2_1 U14421 ( .ip1(n16851), .ip2(\ROUTEDATA/regData [109]), .op(n15358)
         );
  nand2_1 U14422 ( .ip1(n16835), .ip2(\ROUTEDATA/regData [45]), .op(n15357) );
  nand2_1 U14423 ( .ip1(n16855), .ip2(\ROUTEDATA/regData [125]), .op(n15356)
         );
  nand4_1 U14424 ( .ip1(n15359), .ip2(n15358), .ip3(n15357), .ip4(n15356), 
        .op(n15360) );
  not_ab_or_c_or_d U14425 ( .ip1(n16847), .ip2(\ROUTEDATA/regData [93]), .ip3(
        n15361), .ip4(n15360), .op(n15363) );
  nand2_1 U14426 ( .ip1(n16839), .ip2(\ROUTEDATA/regData [61]), .op(n15362) );
  nand3_1 U14427 ( .ip1(n15364), .ip2(n15363), .ip3(n15362), .op(n15365) );
  mux2_1 U14428 ( .ip1(m2DataIn[13]), .ip2(n15365), .s(n15392), .op(n4073) );
  nand2_1 U14429 ( .ip1(n16851), .ip2(\ROUTEDATA/regData [110]), .op(n15377)
         );
  nand2_1 U14430 ( .ip1(\ROUTEDATA/regData [78]), .ip2(n16843), .op(n15368) );
  nand2_1 U14431 ( .ip1(n15379), .ip2(\ROUTEDATA/regData [158]), .op(n15367)
         );
  nand2_1 U14432 ( .ip1(n16859), .ip2(\ROUTEDATA/regData [142]), .op(n15366)
         );
  nand3_1 U14433 ( .ip1(n15368), .ip2(n15367), .ip3(n15366), .op(n15374) );
  nand2_1 U14434 ( .ip1(n16831), .ip2(\ROUTEDATA/regData [30]), .op(n15372) );
  nand2_1 U14435 ( .ip1(n16855), .ip2(\ROUTEDATA/regData [126]), .op(n15371)
         );
  nand2_1 U14436 ( .ip1(n16839), .ip2(\ROUTEDATA/regData [62]), .op(n15370) );
  nand2_1 U14437 ( .ip1(n17243), .ip2(\ROUTEDATA/regData [14]), .op(n15369) );
  nand4_1 U14438 ( .ip1(n15372), .ip2(n15371), .ip3(n15370), .ip4(n15369), 
        .op(n15373) );
  not_ab_or_c_or_d U14439 ( .ip1(n16847), .ip2(\ROUTEDATA/regData [94]), .ip3(
        n15374), .ip4(n15373), .op(n15376) );
  nand2_1 U14440 ( .ip1(n16835), .ip2(\ROUTEDATA/regData [46]), .op(n15375) );
  nand3_1 U14441 ( .ip1(n15377), .ip2(n15376), .ip3(n15375), .op(n15378) );
  mux2_1 U14442 ( .ip1(m2DataIn[14]), .ip2(n15378), .s(n15392), .op(n4072) );
  nand2_1 U14443 ( .ip1(n16855), .ip2(\ROUTEDATA/regData [127]), .op(n15391)
         );
  nand2_1 U14444 ( .ip1(\ROUTEDATA/regData [79]), .ip2(n16843), .op(n15382) );
  nand2_1 U14445 ( .ip1(n15379), .ip2(\ROUTEDATA/regData [159]), .op(n15381)
         );
  nand2_1 U14446 ( .ip1(n16859), .ip2(\ROUTEDATA/regData [143]), .op(n15380)
         );
  nand3_1 U14447 ( .ip1(n15382), .ip2(n15381), .ip3(n15380), .op(n15388) );
  nand2_1 U14448 ( .ip1(n16831), .ip2(\ROUTEDATA/regData [31]), .op(n15386) );
  nand2_1 U14449 ( .ip1(n16835), .ip2(\ROUTEDATA/regData [47]), .op(n15385) );
  nand2_1 U14450 ( .ip1(n16851), .ip2(\ROUTEDATA/regData [111]), .op(n15384)
         );
  nand2_1 U14451 ( .ip1(n17243), .ip2(\ROUTEDATA/regData [15]), .op(n15383) );
  nand4_1 U14452 ( .ip1(n15386), .ip2(n15385), .ip3(n15384), .ip4(n15383), 
        .op(n15387) );
  not_ab_or_c_or_d U14453 ( .ip1(n16847), .ip2(\ROUTEDATA/regData [95]), .ip3(
        n15388), .ip4(n15387), .op(n15390) );
  nand2_1 U14454 ( .ip1(n16839), .ip2(\ROUTEDATA/regData [63]), .op(n15389) );
  nand3_1 U14455 ( .ip1(n15391), .ip2(n15390), .ip3(n15389), .op(n15393) );
  mux2_1 U14456 ( .ip1(m2DataIn[15]), .ip2(n15393), .s(n15392), .op(n4071) );
  nor2_1 U14457 ( .ip1(weight2AddrOffChip[3]), .ip2(n4113), .op(n15406) );
  nand2_1 U14458 ( .ip1(n15409), .ip2(n15406), .op(n15394) );
  mux2_1 U14459 ( .ip1(weight2[0]), .ip2(\WEIGHT_2/mem_w2[0][0] ), .s(n15394), 
        .op(n4070) );
  mux2_1 U14460 ( .ip1(weight2[1]), .ip2(\WEIGHT_2/mem_w2[0][1] ), .s(n15394), 
        .op(n4069) );
  mux2_1 U14461 ( .ip1(weight2[2]), .ip2(\WEIGHT_2/mem_w2[0][2] ), .s(n15394), 
        .op(n4068) );
  mux2_1 U14462 ( .ip1(weight2[3]), .ip2(\WEIGHT_2/mem_w2[0][3] ), .s(n15394), 
        .op(n4067) );
  mux2_1 U14463 ( .ip1(weight2[4]), .ip2(\WEIGHT_2/mem_w2[0][4] ), .s(n15394), 
        .op(n4066) );
  mux2_1 U14464 ( .ip1(weight2[5]), .ip2(\WEIGHT_2/mem_w2[0][5] ), .s(n15394), 
        .op(n4065) );
  mux2_1 U14465 ( .ip1(weight2[6]), .ip2(\WEIGHT_2/mem_w2[0][6] ), .s(n15394), 
        .op(n4064) );
  mux2_1 U14466 ( .ip1(weight2[7]), .ip2(\WEIGHT_2/mem_w2[0][7] ), .s(n15394), 
        .op(n4063) );
  mux2_1 U14467 ( .ip1(weight2[8]), .ip2(\WEIGHT_2/mem_w2[0][8] ), .s(n15394), 
        .op(n4062) );
  mux2_1 U14468 ( .ip1(weight2[9]), .ip2(\WEIGHT_2/mem_w2[0][9] ), .s(n15394), 
        .op(n4061) );
  mux2_1 U14469 ( .ip1(weight2[10]), .ip2(\WEIGHT_2/mem_w2[0][10] ), .s(n15394), .op(n4060) );
  mux2_1 U14470 ( .ip1(weight2[11]), .ip2(\WEIGHT_2/mem_w2[0][11] ), .s(n15394), .op(n4059) );
  mux2_1 U14471 ( .ip1(weight2[12]), .ip2(\WEIGHT_2/mem_w2[0][12] ), .s(n15394), .op(n4058) );
  mux2_1 U14472 ( .ip1(weight2[13]), .ip2(\WEIGHT_2/mem_w2[0][13] ), .s(n15394), .op(n4057) );
  mux2_1 U14473 ( .ip1(weight2[14]), .ip2(\WEIGHT_2/mem_w2[0][14] ), .s(n15394), .op(n4056) );
  mux2_1 U14474 ( .ip1(weight2[15]), .ip2(\WEIGHT_2/mem_w2[0][15] ), .s(n15394), .op(n4055) );
  nand2_1 U14475 ( .ip1(n15411), .ip2(n15406), .op(n15395) );
  mux2_1 U14476 ( .ip1(weight2[0]), .ip2(\WEIGHT_2/mem_w2[1][0] ), .s(n15395), 
        .op(n4054) );
  mux2_1 U14477 ( .ip1(weight2[1]), .ip2(\WEIGHT_2/mem_w2[1][1] ), .s(n15395), 
        .op(n4053) );
  mux2_1 U14478 ( .ip1(weight2[2]), .ip2(\WEIGHT_2/mem_w2[1][2] ), .s(n15395), 
        .op(n4052) );
  mux2_1 U14479 ( .ip1(weight2[3]), .ip2(\WEIGHT_2/mem_w2[1][3] ), .s(n15395), 
        .op(n4051) );
  mux2_1 U14480 ( .ip1(weight2[4]), .ip2(\WEIGHT_2/mem_w2[1][4] ), .s(n15395), 
        .op(n4050) );
  mux2_1 U14481 ( .ip1(weight2[5]), .ip2(\WEIGHT_2/mem_w2[1][5] ), .s(n15395), 
        .op(n4049) );
  mux2_1 U14482 ( .ip1(weight2[6]), .ip2(\WEIGHT_2/mem_w2[1][6] ), .s(n15395), 
        .op(n4048) );
  mux2_1 U14483 ( .ip1(weight2[7]), .ip2(\WEIGHT_2/mem_w2[1][7] ), .s(n15395), 
        .op(n4047) );
  mux2_1 U14484 ( .ip1(weight2[8]), .ip2(\WEIGHT_2/mem_w2[1][8] ), .s(n15395), 
        .op(n4046) );
  mux2_1 U14485 ( .ip1(weight2[9]), .ip2(\WEIGHT_2/mem_w2[1][9] ), .s(n15395), 
        .op(n4045) );
  mux2_1 U14486 ( .ip1(weight2[10]), .ip2(\WEIGHT_2/mem_w2[1][10] ), .s(n15395), .op(n4044) );
  mux2_1 U14487 ( .ip1(weight2[11]), .ip2(\WEIGHT_2/mem_w2[1][11] ), .s(n15395), .op(n4043) );
  mux2_1 U14488 ( .ip1(weight2[12]), .ip2(\WEIGHT_2/mem_w2[1][12] ), .s(n15395), .op(n4042) );
  mux2_1 U14489 ( .ip1(weight2[13]), .ip2(\WEIGHT_2/mem_w2[1][13] ), .s(n15395), .op(n4041) );
  mux2_1 U14490 ( .ip1(weight2[14]), .ip2(\WEIGHT_2/mem_w2[1][14] ), .s(n15395), .op(n4040) );
  mux2_1 U14491 ( .ip1(weight2[15]), .ip2(\WEIGHT_2/mem_w2[1][15] ), .s(n15395), .op(n4039) );
  nand2_1 U14492 ( .ip1(n15396), .ip2(n15406), .op(n15397) );
  mux2_1 U14493 ( .ip1(weight2[0]), .ip2(\WEIGHT_2/mem_w2[2][0] ), .s(n15397), 
        .op(n4038) );
  mux2_1 U14494 ( .ip1(weight2[1]), .ip2(\WEIGHT_2/mem_w2[2][1] ), .s(n15397), 
        .op(n4037) );
  mux2_1 U14495 ( .ip1(weight2[2]), .ip2(\WEIGHT_2/mem_w2[2][2] ), .s(n15397), 
        .op(n4036) );
  mux2_1 U14496 ( .ip1(weight2[3]), .ip2(\WEIGHT_2/mem_w2[2][3] ), .s(n15397), 
        .op(n4035) );
  mux2_1 U14497 ( .ip1(weight2[4]), .ip2(\WEIGHT_2/mem_w2[2][4] ), .s(n15397), 
        .op(n4034) );
  mux2_1 U14498 ( .ip1(weight2[5]), .ip2(\WEIGHT_2/mem_w2[2][5] ), .s(n15397), 
        .op(n4033) );
  mux2_1 U14499 ( .ip1(weight2[6]), .ip2(\WEIGHT_2/mem_w2[2][6] ), .s(n15397), 
        .op(n4032) );
  mux2_1 U14500 ( .ip1(weight2[7]), .ip2(\WEIGHT_2/mem_w2[2][7] ), .s(n15397), 
        .op(n4031) );
  mux2_1 U14501 ( .ip1(weight2[8]), .ip2(\WEIGHT_2/mem_w2[2][8] ), .s(n15397), 
        .op(n4030) );
  mux2_1 U14502 ( .ip1(weight2[9]), .ip2(\WEIGHT_2/mem_w2[2][9] ), .s(n15397), 
        .op(n4029) );
  mux2_1 U14503 ( .ip1(weight2[10]), .ip2(\WEIGHT_2/mem_w2[2][10] ), .s(n15397), .op(n4028) );
  mux2_1 U14504 ( .ip1(weight2[11]), .ip2(\WEIGHT_2/mem_w2[2][11] ), .s(n15397), .op(n4027) );
  mux2_1 U14505 ( .ip1(weight2[12]), .ip2(\WEIGHT_2/mem_w2[2][12] ), .s(n15397), .op(n4026) );
  mux2_1 U14506 ( .ip1(weight2[13]), .ip2(\WEIGHT_2/mem_w2[2][13] ), .s(n15397), .op(n4025) );
  mux2_1 U14507 ( .ip1(weight2[14]), .ip2(\WEIGHT_2/mem_w2[2][14] ), .s(n15397), .op(n4024) );
  mux2_1 U14508 ( .ip1(weight2[15]), .ip2(\WEIGHT_2/mem_w2[2][15] ), .s(n15397), .op(n4023) );
  nand2_1 U14509 ( .ip1(n15398), .ip2(n15406), .op(n15399) );
  mux2_1 U14510 ( .ip1(weight2[0]), .ip2(\WEIGHT_2/mem_w2[3][0] ), .s(n15399), 
        .op(n4022) );
  mux2_1 U14511 ( .ip1(weight2[1]), .ip2(\WEIGHT_2/mem_w2[3][1] ), .s(n15399), 
        .op(n4021) );
  mux2_1 U14512 ( .ip1(weight2[2]), .ip2(\WEIGHT_2/mem_w2[3][2] ), .s(n15399), 
        .op(n4020) );
  mux2_1 U14513 ( .ip1(weight2[3]), .ip2(\WEIGHT_2/mem_w2[3][3] ), .s(n15399), 
        .op(n4019) );
  mux2_1 U14514 ( .ip1(weight2[4]), .ip2(\WEIGHT_2/mem_w2[3][4] ), .s(n15399), 
        .op(n4018) );
  mux2_1 U14515 ( .ip1(weight2[5]), .ip2(\WEIGHT_2/mem_w2[3][5] ), .s(n15399), 
        .op(n4017) );
  mux2_1 U14516 ( .ip1(weight2[6]), .ip2(\WEIGHT_2/mem_w2[3][6] ), .s(n15399), 
        .op(n4016) );
  mux2_1 U14517 ( .ip1(weight2[7]), .ip2(\WEIGHT_2/mem_w2[3][7] ), .s(n15399), 
        .op(n4015) );
  mux2_1 U14518 ( .ip1(weight2[8]), .ip2(\WEIGHT_2/mem_w2[3][8] ), .s(n15399), 
        .op(n4014) );
  mux2_1 U14519 ( .ip1(weight2[9]), .ip2(\WEIGHT_2/mem_w2[3][9] ), .s(n15399), 
        .op(n4013) );
  mux2_1 U14520 ( .ip1(weight2[10]), .ip2(\WEIGHT_2/mem_w2[3][10] ), .s(n15399), .op(n4012) );
  mux2_1 U14521 ( .ip1(weight2[11]), .ip2(\WEIGHT_2/mem_w2[3][11] ), .s(n15399), .op(n4011) );
  mux2_1 U14522 ( .ip1(weight2[12]), .ip2(\WEIGHT_2/mem_w2[3][12] ), .s(n15399), .op(n4010) );
  mux2_1 U14523 ( .ip1(weight2[13]), .ip2(\WEIGHT_2/mem_w2[3][13] ), .s(n15399), .op(n4009) );
  mux2_1 U14524 ( .ip1(weight2[14]), .ip2(\WEIGHT_2/mem_w2[3][14] ), .s(n15399), .op(n4008) );
  mux2_1 U14525 ( .ip1(weight2[15]), .ip2(\WEIGHT_2/mem_w2[3][15] ), .s(n15399), .op(n4007) );
  nand2_1 U14526 ( .ip1(n15400), .ip2(n15406), .op(n15401) );
  mux2_1 U14527 ( .ip1(weight2[0]), .ip2(\WEIGHT_2/mem_w2[4][0] ), .s(n15401), 
        .op(n4006) );
  mux2_1 U14528 ( .ip1(weight2[1]), .ip2(\WEIGHT_2/mem_w2[4][1] ), .s(n15401), 
        .op(n4005) );
  mux2_1 U14529 ( .ip1(weight2[2]), .ip2(\WEIGHT_2/mem_w2[4][2] ), .s(n15401), 
        .op(n4004) );
  mux2_1 U14530 ( .ip1(weight2[3]), .ip2(\WEIGHT_2/mem_w2[4][3] ), .s(n15401), 
        .op(n4003) );
  mux2_1 U14531 ( .ip1(weight2[4]), .ip2(\WEIGHT_2/mem_w2[4][4] ), .s(n15401), 
        .op(n4002) );
  mux2_1 U14532 ( .ip1(weight2[5]), .ip2(\WEIGHT_2/mem_w2[4][5] ), .s(n15401), 
        .op(n4001) );
  mux2_1 U14533 ( .ip1(weight2[6]), .ip2(\WEIGHT_2/mem_w2[4][6] ), .s(n15401), 
        .op(n4000) );
  mux2_1 U14534 ( .ip1(weight2[7]), .ip2(\WEIGHT_2/mem_w2[4][7] ), .s(n15401), 
        .op(n3999) );
  mux2_1 U14535 ( .ip1(weight2[8]), .ip2(\WEIGHT_2/mem_w2[4][8] ), .s(n15401), 
        .op(n3998) );
  mux2_1 U14536 ( .ip1(weight2[9]), .ip2(\WEIGHT_2/mem_w2[4][9] ), .s(n15401), 
        .op(n3997) );
  mux2_1 U14537 ( .ip1(weight2[10]), .ip2(\WEIGHT_2/mem_w2[4][10] ), .s(n15401), .op(n3996) );
  mux2_1 U14538 ( .ip1(weight2[11]), .ip2(\WEIGHT_2/mem_w2[4][11] ), .s(n15401), .op(n3995) );
  mux2_1 U14539 ( .ip1(weight2[12]), .ip2(\WEIGHT_2/mem_w2[4][12] ), .s(n15401), .op(n3994) );
  mux2_1 U14540 ( .ip1(weight2[13]), .ip2(\WEIGHT_2/mem_w2[4][13] ), .s(n15401), .op(n3993) );
  mux2_1 U14541 ( .ip1(weight2[14]), .ip2(\WEIGHT_2/mem_w2[4][14] ), .s(n15401), .op(n3992) );
  mux2_1 U14542 ( .ip1(weight2[15]), .ip2(\WEIGHT_2/mem_w2[4][15] ), .s(n15401), .op(n3991) );
  nand2_1 U14543 ( .ip1(n15402), .ip2(n15406), .op(n15403) );
  mux2_1 U14544 ( .ip1(weight2[0]), .ip2(\WEIGHT_2/mem_w2[5][0] ), .s(n15403), 
        .op(n3990) );
  mux2_1 U14545 ( .ip1(weight2[1]), .ip2(\WEIGHT_2/mem_w2[5][1] ), .s(n15403), 
        .op(n3989) );
  mux2_1 U14546 ( .ip1(weight2[2]), .ip2(\WEIGHT_2/mem_w2[5][2] ), .s(n15403), 
        .op(n3988) );
  mux2_1 U14547 ( .ip1(weight2[3]), .ip2(\WEIGHT_2/mem_w2[5][3] ), .s(n15403), 
        .op(n3987) );
  mux2_1 U14548 ( .ip1(weight2[4]), .ip2(\WEIGHT_2/mem_w2[5][4] ), .s(n15403), 
        .op(n3986) );
  mux2_1 U14549 ( .ip1(weight2[5]), .ip2(\WEIGHT_2/mem_w2[5][5] ), .s(n15403), 
        .op(n3985) );
  mux2_1 U14550 ( .ip1(weight2[6]), .ip2(\WEIGHT_2/mem_w2[5][6] ), .s(n15403), 
        .op(n3984) );
  mux2_1 U14551 ( .ip1(weight2[7]), .ip2(\WEIGHT_2/mem_w2[5][7] ), .s(n15403), 
        .op(n3983) );
  mux2_1 U14552 ( .ip1(weight2[8]), .ip2(\WEIGHT_2/mem_w2[5][8] ), .s(n15403), 
        .op(n3982) );
  mux2_1 U14553 ( .ip1(weight2[9]), .ip2(\WEIGHT_2/mem_w2[5][9] ), .s(n15403), 
        .op(n3981) );
  mux2_1 U14554 ( .ip1(weight2[10]), .ip2(\WEIGHT_2/mem_w2[5][10] ), .s(n15403), .op(n3980) );
  mux2_1 U14555 ( .ip1(weight2[11]), .ip2(\WEIGHT_2/mem_w2[5][11] ), .s(n15403), .op(n3979) );
  mux2_1 U14556 ( .ip1(weight2[12]), .ip2(\WEIGHT_2/mem_w2[5][12] ), .s(n15403), .op(n3978) );
  mux2_1 U14557 ( .ip1(weight2[13]), .ip2(\WEIGHT_2/mem_w2[5][13] ), .s(n15403), .op(n3977) );
  mux2_1 U14558 ( .ip1(weight2[14]), .ip2(\WEIGHT_2/mem_w2[5][14] ), .s(n15403), .op(n3976) );
  mux2_1 U14559 ( .ip1(weight2[15]), .ip2(\WEIGHT_2/mem_w2[5][15] ), .s(n15403), .op(n3975) );
  nand2_1 U14560 ( .ip1(n15404), .ip2(n15406), .op(n15405) );
  mux2_1 U14561 ( .ip1(weight2[0]), .ip2(\WEIGHT_2/mem_w2[6][0] ), .s(n15405), 
        .op(n3974) );
  mux2_1 U14562 ( .ip1(weight2[1]), .ip2(\WEIGHT_2/mem_w2[6][1] ), .s(n15405), 
        .op(n3973) );
  mux2_1 U14563 ( .ip1(weight2[2]), .ip2(\WEIGHT_2/mem_w2[6][2] ), .s(n15405), 
        .op(n3972) );
  mux2_1 U14564 ( .ip1(weight2[3]), .ip2(\WEIGHT_2/mem_w2[6][3] ), .s(n15405), 
        .op(n3971) );
  mux2_1 U14565 ( .ip1(weight2[4]), .ip2(\WEIGHT_2/mem_w2[6][4] ), .s(n15405), 
        .op(n3970) );
  mux2_1 U14566 ( .ip1(weight2[5]), .ip2(\WEIGHT_2/mem_w2[6][5] ), .s(n15405), 
        .op(n3969) );
  mux2_1 U14567 ( .ip1(weight2[6]), .ip2(\WEIGHT_2/mem_w2[6][6] ), .s(n15405), 
        .op(n3968) );
  mux2_1 U14568 ( .ip1(weight2[7]), .ip2(\WEIGHT_2/mem_w2[6][7] ), .s(n15405), 
        .op(n3967) );
  mux2_1 U14569 ( .ip1(weight2[8]), .ip2(\WEIGHT_2/mem_w2[6][8] ), .s(n15405), 
        .op(n3966) );
  mux2_1 U14570 ( .ip1(weight2[9]), .ip2(\WEIGHT_2/mem_w2[6][9] ), .s(n15405), 
        .op(n3965) );
  mux2_1 U14571 ( .ip1(weight2[10]), .ip2(\WEIGHT_2/mem_w2[6][10] ), .s(n15405), .op(n3964) );
  mux2_1 U14572 ( .ip1(weight2[11]), .ip2(\WEIGHT_2/mem_w2[6][11] ), .s(n15405), .op(n3963) );
  mux2_1 U14573 ( .ip1(weight2[12]), .ip2(\WEIGHT_2/mem_w2[6][12] ), .s(n15405), .op(n3962) );
  mux2_1 U14574 ( .ip1(weight2[13]), .ip2(\WEIGHT_2/mem_w2[6][13] ), .s(n15405), .op(n3961) );
  mux2_1 U14575 ( .ip1(weight2[14]), .ip2(\WEIGHT_2/mem_w2[6][14] ), .s(n15405), .op(n3960) );
  mux2_1 U14576 ( .ip1(weight2[15]), .ip2(\WEIGHT_2/mem_w2[6][15] ), .s(n15405), .op(n3959) );
  nand2_1 U14577 ( .ip1(n15407), .ip2(n15406), .op(n15408) );
  mux2_1 U14578 ( .ip1(weight2[0]), .ip2(\WEIGHT_2/mem_w2[7][0] ), .s(n15408), 
        .op(n3958) );
  mux2_1 U14579 ( .ip1(weight2[1]), .ip2(\WEIGHT_2/mem_w2[7][1] ), .s(n15408), 
        .op(n3957) );
  mux2_1 U14580 ( .ip1(weight2[2]), .ip2(\WEIGHT_2/mem_w2[7][2] ), .s(n15408), 
        .op(n3956) );
  mux2_1 U14581 ( .ip1(weight2[3]), .ip2(\WEIGHT_2/mem_w2[7][3] ), .s(n15408), 
        .op(n3955) );
  mux2_1 U14582 ( .ip1(weight2[4]), .ip2(\WEIGHT_2/mem_w2[7][4] ), .s(n15408), 
        .op(n3954) );
  mux2_1 U14583 ( .ip1(weight2[5]), .ip2(\WEIGHT_2/mem_w2[7][5] ), .s(n15408), 
        .op(n3953) );
  mux2_1 U14584 ( .ip1(weight2[6]), .ip2(\WEIGHT_2/mem_w2[7][6] ), .s(n15408), 
        .op(n3952) );
  mux2_1 U14585 ( .ip1(weight2[7]), .ip2(\WEIGHT_2/mem_w2[7][7] ), .s(n15408), 
        .op(n3951) );
  mux2_1 U14586 ( .ip1(weight2[8]), .ip2(\WEIGHT_2/mem_w2[7][8] ), .s(n15408), 
        .op(n3950) );
  mux2_1 U14587 ( .ip1(weight2[9]), .ip2(\WEIGHT_2/mem_w2[7][9] ), .s(n15408), 
        .op(n3949) );
  mux2_1 U14588 ( .ip1(weight2[10]), .ip2(\WEIGHT_2/mem_w2[7][10] ), .s(n15408), .op(n3948) );
  mux2_1 U14589 ( .ip1(weight2[11]), .ip2(\WEIGHT_2/mem_w2[7][11] ), .s(n15408), .op(n3947) );
  mux2_1 U14590 ( .ip1(weight2[12]), .ip2(\WEIGHT_2/mem_w2[7][12] ), .s(n15408), .op(n3946) );
  mux2_1 U14591 ( .ip1(weight2[13]), .ip2(\WEIGHT_2/mem_w2[7][13] ), .s(n15408), .op(n3945) );
  mux2_1 U14592 ( .ip1(weight2[14]), .ip2(\WEIGHT_2/mem_w2[7][14] ), .s(n15408), .op(n3944) );
  mux2_1 U14593 ( .ip1(weight2[15]), .ip2(\WEIGHT_2/mem_w2[7][15] ), .s(n15408), .op(n3943) );
  nand3_1 U14594 ( .ip1(w2SramWeOffChip), .ip2(n15409), .ip3(
        weight2AddrOffChip[3]), .op(n15410) );
  mux2_1 U14595 ( .ip1(weight2[0]), .ip2(\WEIGHT_2/mem_w2[8][0] ), .s(n15410), 
        .op(n3942) );
  mux2_1 U14596 ( .ip1(weight2[1]), .ip2(\WEIGHT_2/mem_w2[8][1] ), .s(n15410), 
        .op(n3941) );
  mux2_1 U14597 ( .ip1(weight2[2]), .ip2(\WEIGHT_2/mem_w2[8][2] ), .s(n15410), 
        .op(n3940) );
  mux2_1 U14598 ( .ip1(weight2[3]), .ip2(\WEIGHT_2/mem_w2[8][3] ), .s(n15410), 
        .op(n3939) );
  mux2_1 U14599 ( .ip1(weight2[4]), .ip2(\WEIGHT_2/mem_w2[8][4] ), .s(n15410), 
        .op(n3938) );
  mux2_1 U14600 ( .ip1(weight2[5]), .ip2(\WEIGHT_2/mem_w2[8][5] ), .s(n15410), 
        .op(n3937) );
  mux2_1 U14601 ( .ip1(weight2[6]), .ip2(\WEIGHT_2/mem_w2[8][6] ), .s(n15410), 
        .op(n3936) );
  mux2_1 U14602 ( .ip1(weight2[7]), .ip2(\WEIGHT_2/mem_w2[8][7] ), .s(n15410), 
        .op(n3935) );
  mux2_1 U14603 ( .ip1(weight2[8]), .ip2(\WEIGHT_2/mem_w2[8][8] ), .s(n15410), 
        .op(n3934) );
  mux2_1 U14604 ( .ip1(weight2[9]), .ip2(\WEIGHT_2/mem_w2[8][9] ), .s(n15410), 
        .op(n3933) );
  mux2_1 U14605 ( .ip1(weight2[10]), .ip2(\WEIGHT_2/mem_w2[8][10] ), .s(n15410), .op(n3932) );
  mux2_1 U14606 ( .ip1(weight2[11]), .ip2(\WEIGHT_2/mem_w2[8][11] ), .s(n15410), .op(n3931) );
  mux2_1 U14607 ( .ip1(weight2[12]), .ip2(\WEIGHT_2/mem_w2[8][12] ), .s(n15410), .op(n3930) );
  mux2_1 U14608 ( .ip1(weight2[13]), .ip2(\WEIGHT_2/mem_w2[8][13] ), .s(n15410), .op(n3929) );
  mux2_1 U14609 ( .ip1(weight2[14]), .ip2(\WEIGHT_2/mem_w2[8][14] ), .s(n15410), .op(n3928) );
  mux2_1 U14610 ( .ip1(weight2[15]), .ip2(\WEIGHT_2/mem_w2[8][15] ), .s(n15410), .op(n3927) );
  nand3_1 U14611 ( .ip1(w2SramWeOffChip), .ip2(n15411), .ip3(
        weight2AddrOffChip[3]), .op(n15412) );
  mux2_1 U14612 ( .ip1(weight2[0]), .ip2(\WEIGHT_2/mem_w2[9][0] ), .s(n15412), 
        .op(n3926) );
  mux2_1 U14613 ( .ip1(weight2[1]), .ip2(\WEIGHT_2/mem_w2[9][1] ), .s(n15412), 
        .op(n3925) );
  mux2_1 U14614 ( .ip1(weight2[2]), .ip2(\WEIGHT_2/mem_w2[9][2] ), .s(n15412), 
        .op(n3924) );
  mux2_1 U14615 ( .ip1(weight2[3]), .ip2(\WEIGHT_2/mem_w2[9][3] ), .s(n15412), 
        .op(n3923) );
  mux2_1 U14616 ( .ip1(weight2[4]), .ip2(\WEIGHT_2/mem_w2[9][4] ), .s(n15412), 
        .op(n3922) );
  mux2_1 U14617 ( .ip1(weight2[5]), .ip2(\WEIGHT_2/mem_w2[9][5] ), .s(n15412), 
        .op(n3921) );
  mux2_1 U14618 ( .ip1(weight2[6]), .ip2(\WEIGHT_2/mem_w2[9][6] ), .s(n15412), 
        .op(n3920) );
  mux2_1 U14619 ( .ip1(weight2[7]), .ip2(\WEIGHT_2/mem_w2[9][7] ), .s(n15412), 
        .op(n3919) );
  mux2_1 U14620 ( .ip1(weight2[8]), .ip2(\WEIGHT_2/mem_w2[9][8] ), .s(n15412), 
        .op(n3918) );
  mux2_1 U14621 ( .ip1(weight2[9]), .ip2(\WEIGHT_2/mem_w2[9][9] ), .s(n15412), 
        .op(n3917) );
  mux2_1 U14622 ( .ip1(weight2[10]), .ip2(\WEIGHT_2/mem_w2[9][10] ), .s(n15412), .op(n3916) );
  mux2_1 U14623 ( .ip1(weight2[11]), .ip2(\WEIGHT_2/mem_w2[9][11] ), .s(n15412), .op(n3915) );
  mux2_1 U14624 ( .ip1(weight2[12]), .ip2(\WEIGHT_2/mem_w2[9][12] ), .s(n15412), .op(n3914) );
  mux2_1 U14625 ( .ip1(weight2[13]), .ip2(\WEIGHT_2/mem_w2[9][13] ), .s(n15412), .op(n3913) );
  mux2_1 U14626 ( .ip1(weight2[14]), .ip2(\WEIGHT_2/mem_w2[9][14] ), .s(n15412), .op(n3912) );
  mux2_1 U14627 ( .ip1(weight2[15]), .ip2(\WEIGHT_2/mem_w2[9][15] ), .s(n15412), .op(n3911) );
  inv_1 U14628 ( .ip(n15413), .op(n15414) );
  nand2_1 U14629 ( .ip1(n15415), .ip2(n15414), .op(n15450) );
  or2_1 U14630 ( .ip1(n15417), .ip2(n15416), .op(n15418) );
  nand2_1 U14631 ( .ip1(n15475), .ip2(n15418), .op(n15479) );
  nand2_1 U14632 ( .ip1(n15479), .ip2(n15419), .op(n15484) );
  nor2_1 U14633 ( .ip1(n15444), .ip2(n15420), .op(n15422) );
  nand4_1 U14634 ( .ip1(n15443), .ip2(n15447), .ip3(n15422), .ip4(n15421), 
        .op(n15452) );
  or2_1 U14635 ( .ip1(n15423), .ip2(n15422), .op(n15424) );
  nand2_1 U14636 ( .ip1(n15452), .ip2(n15424), .op(n15488) );
  nor4_1 U14637 ( .ip1(n15427), .ip2(n15426), .ip3(n15425), .ip4(n15488), .op(
        n15432) );
  inv_1 U14638 ( .ip(n15428), .op(n15430) );
  nand2_1 U14639 ( .ip1(n15430), .ip2(n15429), .op(n15457) );
  nand4_1 U14640 ( .ip1(n15433), .ip2(n15432), .ip3(n15457), .ip4(n15431), 
        .op(n15434) );
  not_ab_or_c_or_d U14641 ( .ip1(n15435), .ip2(n15470), .ip3(n15484), .ip4(
        n15434), .op(n15439) );
  inv_1 U14642 ( .ip(n15436), .op(n15483) );
  nand2_1 U14643 ( .ip1(n15483), .ip2(n15437), .op(n15438) );
  nand4_1 U14644 ( .ip1(n15486), .ip2(n15472), .ip3(n15439), .ip4(n15438), 
        .op(n15440) );
  nor4_1 U14645 ( .ip1(n15442), .ip2(n15441), .ip3(n15450), .ip4(n15440), .op(
        n15448) );
  nand3_1 U14646 ( .ip1(n15445), .ip2(n15444), .ip3(n15443), .op(n15446) );
  nand2_1 U14647 ( .ip1(n15447), .ip2(n15446), .op(n15489) );
  nor2_1 U14648 ( .ip1(n15448), .ip2(n15489), .op(n3910) );
  nand2_1 U14649 ( .ip1(n15449), .ip2(n15485), .op(n15461) );
  nor2_1 U14650 ( .ip1(n15451), .ip2(n15450), .op(n15478) );
  inv_1 U14651 ( .ip(n15452), .op(n15453) );
  not_ab_or_c_or_d U14652 ( .ip1(n15470), .ip2(n15455), .ip3(n15454), .ip4(
        n15453), .op(n15459) );
  not_ab_or_c_or_d U14653 ( .ip1(n15474), .ip2(n15464), .ip3(n15456), .ip4(
        n15484), .op(n15458) );
  nand4_1 U14654 ( .ip1(n15478), .ip2(n15459), .ip3(n15458), .ip4(n15457), 
        .op(n15460) );
  or4_1 U14655 ( .ip1(n15463), .ip2(n15462), .ip3(n15461), .ip4(n15460), .op(
        n3909) );
  and2_1 U14656 ( .ip1(n15465), .ip2(n15464), .op(n15482) );
  nor2_1 U14657 ( .ip1(n15467), .ip2(n15466), .op(n15481) );
  nand2_1 U14658 ( .ip1(n15469), .ip2(n15468), .op(n15471) );
  nand2_1 U14659 ( .ip1(n15471), .ip2(n15470), .op(n15473) );
  nand2_1 U14660 ( .ip1(n15473), .ip2(n15472), .op(n15487) );
  nand2_1 U14661 ( .ip1(n15475), .ip2(n15474), .op(n15477) );
  nand4_1 U14662 ( .ip1(n15479), .ip2(n15478), .ip3(n15477), .ip4(n15476), 
        .op(n15480) );
  or4_1 U14663 ( .ip1(n15482), .ip2(n15481), .ip3(n15487), .ip4(n15480), .op(
        n3907) );
  nor2_1 U14664 ( .ip1(n15484), .ip2(n15483), .op(n15492) );
  nand3_1 U14665 ( .ip1(n15486), .ip2(n15492), .ip3(n15485), .op(n3905) );
  nor3_1 U14666 ( .ip1(n15489), .ip2(n15488), .ip3(n15487), .op(n15490) );
  nand4_1 U14667 ( .ip1(n15493), .ip2(n15492), .ip3(n15491), .ip4(n15490), 
        .op(n15494) );
  nor2_1 U14668 ( .ip1(n3904), .ip2(n15494), .op(n3903) );
  inv_1 U14669 ( .ip(m2DataIn[3]), .op(n16369) );
  nand4_1 U14670 ( .ip1(m2DataIn[2]), .ip2(m2DataIn[1]), .ip3(q_w2[3]), .ip4(
        q_w2[4]), .op(n15516) );
  nor2_1 U14671 ( .ip1(n16369), .ip2(n15516), .op(n15497) );
  nand2_1 U14672 ( .ip1(m2DataIn[4]), .ip2(q_w2[2]), .op(n15526) );
  nand2_1 U14673 ( .ip1(n15516), .ip2(q_w2[3]), .op(n15495) );
  mux2_1 U14674 ( .ip1(n15516), .ip2(n15495), .s(m2DataIn[3]), .op(n15525) );
  nor2_1 U14675 ( .ip1(n15526), .ip2(n15525), .op(n15496) );
  nor2_1 U14676 ( .ip1(n15497), .ip2(n15496), .op(n15604) );
  inv_1 U14677 ( .ip(m2DataIn[0]), .op(n16145) );
  inv_1 U14678 ( .ip(q_w2[4]), .op(n16447) );
  nand2_1 U14679 ( .ip1(m2DataIn[3]), .ip2(q_w2[7]), .op(n15762) );
  nor3_1 U14680 ( .ip1(n16145), .ip2(n16447), .ip3(n15762), .op(n15597) );
  inv_1 U14681 ( .ip(q_w2[7]), .op(n16561) );
  nor2_1 U14682 ( .ip1(n16145), .ip2(n16561), .op(n15498) );
  or2_1 U14683 ( .ip1(q_w2[4]), .ip2(n15498), .op(n15500) );
  or2_1 U14684 ( .ip1(m2DataIn[3]), .ip2(n15498), .op(n15499) );
  nand2_1 U14685 ( .ip1(n15500), .ip2(n15499), .op(n15595) );
  nor2_1 U14686 ( .ip1(n15597), .ip2(n15595), .op(n15501) );
  nand2_1 U14687 ( .ip1(m2DataIn[2]), .ip2(q_w2[5]), .op(n15594) );
  xor2_1 U14688 ( .ip1(n15501), .ip2(n15594), .op(n15603) );
  inv_1 U14689 ( .ip(m2DataIn[5]), .op(n16496) );
  inv_1 U14690 ( .ip(q_w2[3]), .op(n16177) );
  nor3_1 U14691 ( .ip1(n16496), .ip2(n16177), .ip3(n15526), .op(n15601) );
  nor2_1 U14692 ( .ip1(n16445), .ip2(n16177), .op(n15502) );
  or2_1 U14693 ( .ip1(q_w2[2]), .ip2(n15502), .op(n15504) );
  or2_1 U14694 ( .ip1(m2DataIn[5]), .ip2(n15502), .op(n15503) );
  nand2_1 U14695 ( .ip1(n15504), .ip2(n15503), .op(n15599) );
  nor2_1 U14696 ( .ip1(n15601), .ip2(n15599), .op(n15505) );
  nand2_1 U14697 ( .ip1(m2DataIn[7]), .ip2(q_w2[0]), .op(n15598) );
  xor2_1 U14698 ( .ip1(n15505), .ip2(n15598), .op(n15602) );
  inv_1 U14699 ( .ip(n15506), .op(n15622) );
  inv_1 U14700 ( .ip(q_w2[5]), .op(n16497) );
  nor2_1 U14701 ( .ip1(n16145), .ip2(n16497), .op(n15531) );
  inv_1 U14702 ( .ip(q_w2[2]), .op(n16308) );
  nor2_1 U14703 ( .ip1(n16369), .ip2(n16308), .op(n15530) );
  inv_1 U14704 ( .ip(q_w2[0]), .op(n15973) );
  nor2_1 U14705 ( .ip1(n16496), .ip2(n15973), .op(n15529) );
  nand2_1 U14706 ( .ip1(m2DataIn[2]), .ip2(q_w2[4]), .op(n15507) );
  inv_1 U14707 ( .ip(m2DataIn[2]), .op(n16309) );
  inv_1 U14708 ( .ip(m2DataIn[1]), .op(n16222) );
  nor4_1 U14709 ( .ip1(n16309), .ip2(n16222), .ip3(n16447), .ip4(n16497), .op(
        n15592) );
  or2_1 U14710 ( .ip1(n15507), .ip2(n15592), .op(n15510) );
  nand2_1 U14711 ( .ip1(m2DataIn[1]), .ip2(q_w2[5]), .op(n15508) );
  or2_1 U14712 ( .ip1(n15508), .ip2(n15592), .op(n15509) );
  nand2_1 U14713 ( .ip1(n15510), .ip2(n15509), .op(n15523) );
  inv_1 U14714 ( .ip(q_w2[6]), .op(n16538) );
  nor2_1 U14715 ( .ip1(n16145), .ip2(n16538), .op(n15691) );
  inv_1 U14716 ( .ip(q_w2[1]), .op(n16144) );
  nor2_1 U14717 ( .ip1(n16496), .ip2(n16144), .op(n15515) );
  nor2_1 U14718 ( .ip1(n16273), .ip2(n15973), .op(n15514) );
  and3_1 U14719 ( .ip1(m2DataIn[1]), .ip2(q_w2[6]), .ip3(n15511), .op(n15661)
         );
  nor2_1 U14720 ( .ip1(n16222), .ip2(n16538), .op(n15512) );
  nor2_1 U14721 ( .ip1(n15512), .ip2(n15511), .op(n15513) );
  nor2_1 U14722 ( .ip1(n15661), .ip2(n15513), .op(n15621) );
  fulladder U14723 ( .a(n15691), .b(n15515), .ci(n15514), .co(n15591), .s(
        n15522) );
  nor2_1 U14724 ( .ip1(n16273), .ip2(n16144), .op(n15590) );
  nand2_1 U14725 ( .ip1(m2DataIn[1]), .ip2(q_w2[2]), .op(n15548) );
  nor3_1 U14726 ( .ip1(n16309), .ip2(n16177), .ip3(n15548), .op(n15539) );
  inv_1 U14727 ( .ip(n15516), .op(n15521) );
  nor2_1 U14728 ( .ip1(n16309), .ip2(n16177), .op(n15517) );
  or2_1 U14729 ( .ip1(q_w2[4]), .ip2(n15517), .op(n15519) );
  or2_1 U14730 ( .ip1(m2DataIn[1]), .ip2(n15517), .op(n15518) );
  nand2_1 U14731 ( .ip1(n15519), .ip2(n15518), .op(n15520) );
  nor2_1 U14732 ( .ip1(n15521), .ip2(n15520), .op(n15528) );
  nor2_1 U14733 ( .ip1(n16445), .ip2(n16144), .op(n15527) );
  fulladder U14734 ( .a(n15524), .b(n15523), .ci(n15522), .co(n15511), .s(
        n15541) );
  xor2_1 U14735 ( .ip1(n15526), .ip2(n15525), .op(n15540) );
  fulladder U14736 ( .a(n15539), .b(n15528), .ci(n15527), .co(n15542), .s(
        n15545) );
  nor2_1 U14737 ( .ip1(n16145), .ip2(n16447), .op(n15534) );
  nor2_1 U14738 ( .ip1(n16369), .ip2(n16144), .op(n15533) );
  nor2_1 U14739 ( .ip1(n16445), .ip2(n15973), .op(n15532) );
  fulladder U14740 ( .a(n15531), .b(n15530), .ci(n15529), .co(n15524), .s(
        n15543) );
  fulladder U14741 ( .a(n15534), .b(n15533), .ci(n15532), .co(n15544), .s(
        n15547) );
  nor4_1 U14742 ( .ip1(n16369), .ip2(n16222), .ip3(n15973), .ip4(n16308), .op(
        n15549) );
  nor2_1 U14743 ( .ip1(n16222), .ip2(n16177), .op(n15535) );
  or2_1 U14744 ( .ip1(q_w2[2]), .ip2(n15535), .op(n15537) );
  or2_1 U14745 ( .ip1(m2DataIn[2]), .ip2(n15535), .op(n15536) );
  nand2_1 U14746 ( .ip1(n15537), .ip2(n15536), .op(n15538) );
  nor2_1 U14747 ( .ip1(n15539), .ip2(n15538), .op(n15546) );
  fulladder U14748 ( .a(n15542), .b(n15541), .ci(n15540), .co(n15587), .s(
        n15583) );
  fulladder U14749 ( .a(n15545), .b(n15544), .ci(n15543), .co(n15582), .s(
        n15576) );
  or2_1 U14750 ( .ip1(n15583), .ip2(n15582), .op(n15579) );
  nand3_1 U14751 ( .ip1(n15576), .ip2(n15575), .ip3(n15579), .op(n15581) );
  fulladder U14752 ( .a(n15547), .b(n15549), .ci(n15546), .co(n15575), .s(
        n15569) );
  or2_1 U14753 ( .ip1(n15548), .ip2(n15549), .op(n15552) );
  nand2_1 U14754 ( .ip1(m2DataIn[3]), .ip2(q_w2[0]), .op(n15550) );
  or2_1 U14755 ( .ip1(n15550), .ip2(n15549), .op(n15551) );
  nand2_1 U14756 ( .ip1(n15552), .ip2(n15551), .op(n15559) );
  nand2_1 U14757 ( .ip1(m2DataIn[2]), .ip2(q_w2[1]), .op(n15567) );
  nor2_1 U14758 ( .ip1(n16145), .ip2(n16177), .op(n15565) );
  nor4_1 U14759 ( .ip1(n16309), .ip2(n16222), .ip3(n15973), .ip4(n16144), .op(
        n15566) );
  xnor2_1 U14760 ( .ip1(n15565), .ip2(n15566), .op(n15553) );
  xor2_1 U14761 ( .ip1(n15567), .ip2(n15553), .op(n15561) );
  nand2_1 U14762 ( .ip1(n15559), .ip2(n15561), .op(n15564) );
  nand2_1 U14763 ( .ip1(m2DataIn[2]), .ip2(q_w2[0]), .op(n15558) );
  nand2_1 U14764 ( .ip1(m2DataIn[1]), .ip2(q_w2[1]), .op(n15557) );
  or2_1 U14765 ( .ip1(q_w2[0]), .ip2(q_w2[2]), .op(n15555) );
  or2_1 U14766 ( .ip1(n16309), .ip2(q_w2[2]), .op(n15554) );
  nand2_1 U14767 ( .ip1(n15555), .ip2(n15554), .op(n15556) );
  not_ab_or_c_or_d U14768 ( .ip1(n15558), .ip2(n15557), .ip3(n15556), .ip4(
        n16145), .op(n15560) );
  nand2_1 U14769 ( .ip1(n15559), .ip2(n15560), .op(n15563) );
  nand2_1 U14770 ( .ip1(n15561), .ip2(n15560), .op(n15562) );
  nand3_1 U14771 ( .ip1(n15564), .ip2(n15563), .ip3(n15562), .op(n15571) );
  nand2_1 U14772 ( .ip1(n15569), .ip2(n15571), .op(n15574) );
  nor2_1 U14773 ( .ip1(n15566), .ip2(n15565), .op(n15568) );
  nor2_1 U14774 ( .ip1(n15568), .ip2(n15567), .op(n15570) );
  nand2_1 U14775 ( .ip1(n15569), .ip2(n15570), .op(n15573) );
  nand2_1 U14776 ( .ip1(n15571), .ip2(n15570), .op(n15572) );
  nand3_1 U14777 ( .ip1(n15574), .ip2(n15573), .ip3(n15572), .op(n15578) );
  or2_1 U14778 ( .ip1(n15576), .ip2(n15575), .op(n15577) );
  nand3_1 U14779 ( .ip1(n15579), .ip2(n15578), .ip3(n15577), .op(n15580) );
  nand2_1 U14780 ( .ip1(n15581), .ip2(n15580), .op(n15585) );
  and2_1 U14781 ( .ip1(n15583), .ip2(n15582), .op(n15584) );
  not_ab_or_c_or_d U14782 ( .ip1(n15586), .ip2(n15587), .ip3(n15585), .ip4(
        n15584), .op(n15589) );
  nor2_1 U14783 ( .ip1(n15587), .ip2(n15586), .op(n15588) );
  nor2_1 U14784 ( .ip1(n15589), .ip2(n15588), .op(n15712) );
  fulladder U14785 ( .a(n15592), .b(n15591), .ci(n15590), .co(n15593), .s(
        n15620) );
  inv_1 U14786 ( .ip(n15593), .op(n15708) );
  nor2_1 U14787 ( .ip1(n15595), .ip2(n15594), .op(n15596) );
  nor2_1 U14788 ( .ip1(n15597), .ip2(n15596), .op(n15705) );
  nand2_1 U14789 ( .ip1(m2DataIn[6]), .ip2(q_w2[2]), .op(n15704) );
  nor2_1 U14790 ( .ip1(n15599), .ip2(n15598), .op(n15600) );
  nor2_1 U14791 ( .ip1(n15601), .ip2(n15600), .op(n15703) );
  fulladder U14792 ( .a(n15604), .b(n15603), .ci(n15602), .co(n15706), .s(
        n15506) );
  inv_1 U14793 ( .ip(n15605), .op(n15662) );
  nand2_1 U14794 ( .ip1(m2DataIn[4]), .ip2(q_w2[4]), .op(n15606) );
  nand2_1 U14795 ( .ip1(m2DataIn[5]), .ip2(q_w2[4]), .op(n15698) );
  nor3_1 U14796 ( .ip1(n16445), .ip2(n16177), .ip3(n15698), .op(n15664) );
  or2_1 U14797 ( .ip1(n15606), .ip2(n15664), .op(n15609) );
  nand2_1 U14798 ( .ip1(m2DataIn[5]), .ip2(q_w2[3]), .op(n15607) );
  or2_1 U14799 ( .ip1(n15607), .ip2(n15664), .op(n15608) );
  nand2_1 U14800 ( .ip1(n15609), .ip2(n15608), .op(n15663) );
  inv_1 U14801 ( .ip(m2DataIn[7]), .op(n16550) );
  nor2_1 U14802 ( .ip1(n16550), .ip2(n16144), .op(n15665) );
  xor2_1 U14803 ( .ip1(n15663), .ip2(n15665), .op(n15689) );
  nand2_1 U14804 ( .ip1(m2DataIn[3]), .ip2(q_w2[8]), .op(n15790) );
  nor3_1 U14805 ( .ip1(n16145), .ip2(n16497), .ip3(n15790), .op(n15672) );
  inv_1 U14806 ( .ip(q_w2[8]), .op(n16596) );
  nor2_1 U14807 ( .ip1(n16145), .ip2(n16596), .op(n15610) );
  or2_1 U14808 ( .ip1(q_w2[5]), .ip2(n15610), .op(n15612) );
  or2_1 U14809 ( .ip1(m2DataIn[3]), .ip2(n15610), .op(n15611) );
  nand2_1 U14810 ( .ip1(n15612), .ip2(n15611), .op(n15613) );
  nor2_1 U14811 ( .ip1(n15672), .ip2(n15613), .op(n15671) );
  inv_1 U14812 ( .ip(m2DataIn[8]), .op(n16624) );
  nor2_1 U14813 ( .ip1(n16624), .ip2(n15973), .op(n15673) );
  xor2_1 U14814 ( .ip1(n15671), .ip2(n15673), .op(n15688) );
  inv_1 U14815 ( .ip(rdata[0]), .op(n15616) );
  nand2_1 U14816 ( .ip1(q_w2[6]), .ip2(m2DataIn[2]), .op(n15615) );
  nor2_1 U14817 ( .ip1(n16222), .ip2(n16561), .op(n15614) );
  xor2_1 U14818 ( .ip1(n15615), .ip2(n15614), .op(n15617) );
  nor2_1 U14819 ( .ip1(n15616), .ip2(n15617), .op(n15677) );
  or2_1 U14820 ( .ip1(n15616), .ip2(n15677), .op(n15619) );
  or2_1 U14821 ( .ip1(n15617), .ip2(n15677), .op(n15618) );
  nand2_1 U14822 ( .ip1(n15619), .ip2(n15618), .op(n15687) );
  fulladder U14823 ( .a(n15622), .b(n15621), .ci(n15620), .co(n15710), .s(
        n15586) );
  mux2_1 U14824 ( .ip1(n15623), .ip2(\SIGMOID/N64 ), .s(n16714), .op(n15644)
         );
  buf_1 U14825 ( .ip(n15644), .op(n15653) );
  and2_1 U14826 ( .ip1(n18800), .ip2(n18888), .op(n15647) );
  or2_1 U14827 ( .ip1(n15624), .ip2(n16714), .op(n15626) );
  or2_1 U14828 ( .ip1(\CNTRL/count_20Q [0]), .ip2(n16714), .op(n15625) );
  nand2_1 U14829 ( .ip1(n15626), .ip2(n15625), .op(n15641) );
  nor2_1 U14830 ( .ip1(n15641), .ip2(n18901), .op(n15627) );
  nand2_1 U14831 ( .ip1(n15627), .ip2(n17488), .op(n15646) );
  buf_1 U14832 ( .ip(n17506), .op(n17564) );
  inv_1 U14833 ( .ip(n18165), .op(n18092) );
  nor3_1 U14834 ( .ip1(n15646), .ip2(n17564), .ip3(n18092), .op(n15631) );
  nand2_1 U14835 ( .ip1(n15647), .ip2(n15631), .op(n16717) );
  mux2_1 U14836 ( .ip1(n15653), .ip2(\ANSWER/mem[0][0][0] ), .s(n16717), .op(
        n3902) );
  nand2_1 U14837 ( .ip1(n15631), .ip2(n15648), .op(n16718) );
  mux2_1 U14838 ( .ip1(n15653), .ip2(\ANSWER/mem[0][1][0] ), .s(n16718), .op(
        n3901) );
  and2_1 U14839 ( .ip1(n18888), .ip2(n18884), .op(n15649) );
  nand2_1 U14840 ( .ip1(n15631), .ip2(n15649), .op(n16719) );
  mux2_1 U14841 ( .ip1(n15653), .ip2(\ANSWER/mem[0][2][0] ), .s(n16719), .op(
        n3900) );
  and2_1 U14842 ( .ip1(n18888), .ip2(n18854), .op(n15650) );
  nand2_1 U14843 ( .ip1(n15631), .ip2(n15650), .op(n16720) );
  mux2_1 U14844 ( .ip1(n15653), .ip2(\ANSWER/mem[0][3][0] ), .s(n16720), .op(
        n3899) );
  and2_1 U14845 ( .ip1(n18888), .ip2(n18843), .op(n15651) );
  nand2_1 U14846 ( .ip1(n15631), .ip2(n15651), .op(n16721) );
  mux2_1 U14847 ( .ip1(n15653), .ip2(\ANSWER/mem[0][4][0] ), .s(n16721), .op(
        n3898) );
  and2_1 U14848 ( .ip1(n18888), .ip2(n18832), .op(n15652) );
  nand2_1 U14849 ( .ip1(n15631), .ip2(n15652), .op(n16722) );
  mux2_1 U14850 ( .ip1(n15653), .ip2(\ANSWER/mem[0][5][0] ), .s(n16722), .op(
        n3897) );
  and2_1 U14851 ( .ip1(n18888), .ip2(n18821), .op(n15654) );
  nand2_1 U14852 ( .ip1(n15631), .ip2(n15654), .op(n16723) );
  mux2_1 U14853 ( .ip1(n15653), .ip2(\ANSWER/mem[0][6][0] ), .s(n16723), .op(
        n3896) );
  and2_1 U14854 ( .ip1(n18888), .ip2(n18865), .op(n15655) );
  nand2_1 U14855 ( .ip1(n15631), .ip2(n15655), .op(n16724) );
  mux2_1 U14856 ( .ip1(n15653), .ip2(\ANSWER/mem[0][7][0] ), .s(n16724), .op(
        n3895) );
  inv_1 U14857 ( .ip(n18914), .op(n15628) );
  nor2_1 U14858 ( .ip1(n15630), .ip2(n15628), .op(n15656) );
  nand2_1 U14859 ( .ip1(n15631), .ip2(n15656), .op(n16725) );
  mux2_1 U14860 ( .ip1(n15653), .ip2(\ANSWER/mem[0][8][0] ), .s(n16725), .op(
        n3894) );
  inv_1 U14861 ( .ip(n18899), .op(n15629) );
  nor2_1 U14862 ( .ip1(n15630), .ip2(n15629), .op(n15658) );
  nand2_1 U14863 ( .ip1(n15631), .ip2(n15658), .op(n16726) );
  mux2_1 U14864 ( .ip1(n15653), .ip2(\ANSWER/mem[0][9][0] ), .s(n16726), .op(
        n3893) );
  nor3_1 U14865 ( .ip1(n4362), .ip2(n15646), .ip3(n18092), .op(n15632) );
  nand2_1 U14866 ( .ip1(n15647), .ip2(n15632), .op(n16727) );
  mux2_1 U14867 ( .ip1(n15653), .ip2(\ANSWER/mem[1][0][0] ), .s(n16727), .op(
        n3892) );
  nand2_1 U14868 ( .ip1(n15648), .ip2(n15632), .op(n16728) );
  mux2_1 U14869 ( .ip1(n15653), .ip2(\ANSWER/mem[1][1][0] ), .s(n16728), .op(
        n3891) );
  buf_1 U14870 ( .ip(n15644), .op(n15659) );
  nand2_1 U14871 ( .ip1(n15649), .ip2(n15632), .op(n16729) );
  mux2_1 U14872 ( .ip1(n15659), .ip2(\ANSWER/mem[1][2][0] ), .s(n16729), .op(
        n3890) );
  nand2_1 U14873 ( .ip1(n15650), .ip2(n15632), .op(n16730) );
  mux2_1 U14874 ( .ip1(n15659), .ip2(\ANSWER/mem[1][3][0] ), .s(n16730), .op(
        n3889) );
  nand2_1 U14875 ( .ip1(n15651), .ip2(n15632), .op(n16731) );
  mux2_1 U14876 ( .ip1(n15644), .ip2(\ANSWER/mem[1][4][0] ), .s(n16731), .op(
        n3888) );
  nand2_1 U14877 ( .ip1(n15652), .ip2(n15632), .op(n16732) );
  mux2_1 U14878 ( .ip1(n15644), .ip2(\ANSWER/mem[1][5][0] ), .s(n16732), .op(
        n3887) );
  nand2_1 U14879 ( .ip1(n15654), .ip2(n15632), .op(n16733) );
  mux2_1 U14880 ( .ip1(n15644), .ip2(\ANSWER/mem[1][6][0] ), .s(n16733), .op(
        n3886) );
  nand2_1 U14881 ( .ip1(n15655), .ip2(n15632), .op(n16734) );
  mux2_1 U14882 ( .ip1(n15644), .ip2(\ANSWER/mem[1][7][0] ), .s(n16734), .op(
        n3885) );
  nand2_1 U14883 ( .ip1(n15656), .ip2(n15632), .op(n16735) );
  mux2_1 U14884 ( .ip1(n15644), .ip2(\ANSWER/mem[1][8][0] ), .s(n16735), .op(
        n3884) );
  nand2_1 U14885 ( .ip1(n15658), .ip2(n15632), .op(n16736) );
  mux2_1 U14886 ( .ip1(n15644), .ip2(\ANSWER/mem[1][9][0] ), .s(n16736), .op(
        n3883) );
  buf_1 U14887 ( .ip(n18878), .op(n18815) );
  nand2_1 U14888 ( .ip1(n4362), .ip2(n18165), .op(n15638) );
  nor4_1 U14889 ( .ip1(n15641), .ip2(n4366), .ip3(n18815), .ip4(n15638), .op(
        n15633) );
  nand2_1 U14890 ( .ip1(n15647), .ip2(n15633), .op(n16737) );
  mux2_1 U14891 ( .ip1(n15644), .ip2(\ANSWER/mem[2][0][0] ), .s(n16737), .op(
        n3882) );
  nand2_1 U14892 ( .ip1(n15648), .ip2(n15633), .op(n16738) );
  mux2_1 U14893 ( .ip1(n15644), .ip2(\ANSWER/mem[2][1][0] ), .s(n16738), .op(
        n3881) );
  nand2_1 U14894 ( .ip1(n15649), .ip2(n15633), .op(n16739) );
  mux2_1 U14895 ( .ip1(n15644), .ip2(\ANSWER/mem[2][2][0] ), .s(n16739), .op(
        n3880) );
  nand2_1 U14896 ( .ip1(n15650), .ip2(n15633), .op(n16740) );
  mux2_1 U14897 ( .ip1(n15644), .ip2(\ANSWER/mem[2][3][0] ), .s(n16740), .op(
        n3879) );
  nand2_1 U14898 ( .ip1(n15651), .ip2(n15633), .op(n16741) );
  mux2_1 U14899 ( .ip1(n15659), .ip2(\ANSWER/mem[2][4][0] ), .s(n16741), .op(
        n3878) );
  nand2_1 U14900 ( .ip1(n15652), .ip2(n15633), .op(n16742) );
  mux2_1 U14901 ( .ip1(n15653), .ip2(\ANSWER/mem[2][5][0] ), .s(n16742), .op(
        n3877) );
  nand2_1 U14902 ( .ip1(n15654), .ip2(n15633), .op(n16743) );
  mux2_1 U14903 ( .ip1(n15653), .ip2(\ANSWER/mem[2][6][0] ), .s(n16743), .op(
        n3876) );
  nand2_1 U14904 ( .ip1(n15655), .ip2(n15633), .op(n16744) );
  mux2_1 U14905 ( .ip1(n15644), .ip2(\ANSWER/mem[2][7][0] ), .s(n16744), .op(
        n3875) );
  nand2_1 U14906 ( .ip1(n15656), .ip2(n15633), .op(n16745) );
  mux2_1 U14907 ( .ip1(n15659), .ip2(\ANSWER/mem[2][8][0] ), .s(n16745), .op(
        n3874) );
  nand2_1 U14908 ( .ip1(n15658), .ip2(n15633), .op(n16746) );
  mux2_1 U14909 ( .ip1(n15653), .ip2(\ANSWER/mem[2][9][0] ), .s(n16746), .op(
        n3873) );
  buf_1 U14910 ( .ip(n18878), .op(n18837) );
  nand2_1 U14911 ( .ip1(n18165), .ip2(n17610), .op(n15640) );
  nor4_1 U14912 ( .ip1(n15641), .ip2(n4366), .ip3(n18837), .ip4(n15640), .op(
        n15634) );
  nand2_1 U14913 ( .ip1(n15647), .ip2(n15634), .op(n16747) );
  mux2_1 U14914 ( .ip1(n15659), .ip2(\ANSWER/mem[3][0][0] ), .s(n16747), .op(
        n3872) );
  nand2_1 U14915 ( .ip1(n15648), .ip2(n15634), .op(n16748) );
  mux2_1 U14916 ( .ip1(n15644), .ip2(\ANSWER/mem[3][1][0] ), .s(n16748), .op(
        n3871) );
  nand2_1 U14917 ( .ip1(n15649), .ip2(n15634), .op(n16749) );
  mux2_1 U14918 ( .ip1(n15644), .ip2(\ANSWER/mem[3][2][0] ), .s(n16749), .op(
        n3870) );
  nand2_1 U14919 ( .ip1(n15650), .ip2(n15634), .op(n16750) );
  mux2_1 U14920 ( .ip1(n15644), .ip2(\ANSWER/mem[3][3][0] ), .s(n16750), .op(
        n3869) );
  nand2_1 U14921 ( .ip1(n15651), .ip2(n15634), .op(n16751) );
  mux2_1 U14922 ( .ip1(n15644), .ip2(\ANSWER/mem[3][4][0] ), .s(n16751), .op(
        n3868) );
  nand2_1 U14923 ( .ip1(n15652), .ip2(n15634), .op(n16752) );
  mux2_1 U14924 ( .ip1(n15644), .ip2(\ANSWER/mem[3][5][0] ), .s(n16752), .op(
        n3867) );
  nand2_1 U14925 ( .ip1(n15654), .ip2(n15634), .op(n16753) );
  mux2_1 U14926 ( .ip1(n15659), .ip2(\ANSWER/mem[3][6][0] ), .s(n16753), .op(
        n3866) );
  nand2_1 U14927 ( .ip1(n15655), .ip2(n15634), .op(n16754) );
  mux2_1 U14928 ( .ip1(n15659), .ip2(\ANSWER/mem[3][7][0] ), .s(n16754), .op(
        n3865) );
  nand2_1 U14929 ( .ip1(n15656), .ip2(n15634), .op(n16755) );
  mux2_1 U14930 ( .ip1(n15659), .ip2(\ANSWER/mem[3][8][0] ), .s(n16755), .op(
        n3864) );
  nand2_1 U14931 ( .ip1(n15658), .ip2(n15634), .op(n16756) );
  mux2_1 U14932 ( .ip1(n15659), .ip2(\ANSWER/mem[3][9][0] ), .s(n16756), .op(
        n3863) );
  nor4_1 U14933 ( .ip1(n15641), .ip2(n17488), .ip3(n15636), .ip4(n15638), .op(
        n15635) );
  nand2_1 U14934 ( .ip1(n15647), .ip2(n15635), .op(n16757) );
  mux2_1 U14935 ( .ip1(n15659), .ip2(\ANSWER/mem[4][0][0] ), .s(n16757), .op(
        n3862) );
  nand2_1 U14936 ( .ip1(n15648), .ip2(n15635), .op(n16758) );
  mux2_1 U14937 ( .ip1(n15659), .ip2(\ANSWER/mem[4][1][0] ), .s(n16758), .op(
        n3861) );
  nand2_1 U14938 ( .ip1(n15649), .ip2(n15635), .op(n16759) );
  mux2_1 U14939 ( .ip1(n15653), .ip2(\ANSWER/mem[4][2][0] ), .s(n16759), .op(
        n3860) );
  nand2_1 U14940 ( .ip1(n15650), .ip2(n15635), .op(n16760) );
  mux2_1 U14941 ( .ip1(n15644), .ip2(\ANSWER/mem[4][3][0] ), .s(n16760), .op(
        n3859) );
  nand2_1 U14942 ( .ip1(n15651), .ip2(n15635), .op(n16761) );
  mux2_1 U14943 ( .ip1(n15659), .ip2(\ANSWER/mem[4][4][0] ), .s(n16761), .op(
        n3858) );
  nand2_1 U14944 ( .ip1(n15652), .ip2(n15635), .op(n16762) );
  mux2_1 U14945 ( .ip1(n15659), .ip2(\ANSWER/mem[4][5][0] ), .s(n16762), .op(
        n3857) );
  nand2_1 U14946 ( .ip1(n15654), .ip2(n15635), .op(n16763) );
  mux2_1 U14947 ( .ip1(n15644), .ip2(\ANSWER/mem[4][6][0] ), .s(n16763), .op(
        n3856) );
  nand2_1 U14948 ( .ip1(n15655), .ip2(n15635), .op(n16764) );
  mux2_1 U14949 ( .ip1(n15659), .ip2(\ANSWER/mem[4][7][0] ), .s(n16764), .op(
        n3855) );
  nand2_1 U14950 ( .ip1(n15656), .ip2(n15635), .op(n16765) );
  mux2_1 U14951 ( .ip1(n15659), .ip2(\ANSWER/mem[4][8][0] ), .s(n16765), .op(
        n3854) );
  nand2_1 U14952 ( .ip1(n15658), .ip2(n15635), .op(n16766) );
  mux2_1 U14953 ( .ip1(n15644), .ip2(\ANSWER/mem[4][9][0] ), .s(n16766), .op(
        n3853) );
  nor4_1 U14954 ( .ip1(n15641), .ip2(n17488), .ip3(n15636), .ip4(n15640), .op(
        n15637) );
  nand2_1 U14955 ( .ip1(n15647), .ip2(n15637), .op(n16767) );
  mux2_1 U14956 ( .ip1(n15644), .ip2(\ANSWER/mem[5][0][0] ), .s(n16767), .op(
        n3852) );
  nand2_1 U14957 ( .ip1(n15648), .ip2(n15637), .op(n16768) );
  mux2_1 U14958 ( .ip1(n15659), .ip2(\ANSWER/mem[5][1][0] ), .s(n16768), .op(
        n3851) );
  nand2_1 U14959 ( .ip1(n15649), .ip2(n15637), .op(n16769) );
  mux2_1 U14960 ( .ip1(n15644), .ip2(\ANSWER/mem[5][2][0] ), .s(n16769), .op(
        n3850) );
  nand2_1 U14961 ( .ip1(n15650), .ip2(n15637), .op(n16770) );
  mux2_1 U14962 ( .ip1(n15644), .ip2(\ANSWER/mem[5][3][0] ), .s(n16770), .op(
        n3849) );
  nand2_1 U14963 ( .ip1(n15651), .ip2(n15637), .op(n16771) );
  mux2_1 U14964 ( .ip1(n15659), .ip2(\ANSWER/mem[5][4][0] ), .s(n16771), .op(
        n3848) );
  nand2_1 U14965 ( .ip1(n15652), .ip2(n15637), .op(n16772) );
  mux2_1 U14966 ( .ip1(n15644), .ip2(\ANSWER/mem[5][5][0] ), .s(n16772), .op(
        n3847) );
  nand2_1 U14967 ( .ip1(n15654), .ip2(n15637), .op(n16773) );
  mux2_1 U14968 ( .ip1(n15644), .ip2(\ANSWER/mem[5][6][0] ), .s(n16773), .op(
        n3846) );
  nand2_1 U14969 ( .ip1(n15655), .ip2(n15637), .op(n16774) );
  mux2_1 U14970 ( .ip1(n15659), .ip2(\ANSWER/mem[5][7][0] ), .s(n16774), .op(
        n3845) );
  nand2_1 U14971 ( .ip1(n15656), .ip2(n15637), .op(n16775) );
  mux2_1 U14972 ( .ip1(n15644), .ip2(\ANSWER/mem[5][8][0] ), .s(n16775), .op(
        n3844) );
  nand2_1 U14973 ( .ip1(n15658), .ip2(n15637), .op(n16776) );
  mux2_1 U14974 ( .ip1(n15644), .ip2(\ANSWER/mem[5][9][0] ), .s(n16776), .op(
        n3843) );
  nor4_1 U14975 ( .ip1(n15641), .ip2(n4366), .ip3(n17488), .ip4(n15638), .op(
        n15639) );
  nand2_1 U14976 ( .ip1(n15647), .ip2(n15639), .op(n16777) );
  mux2_1 U14977 ( .ip1(n15653), .ip2(\ANSWER/mem[6][0][0] ), .s(n16777), .op(
        n3842) );
  nand2_1 U14978 ( .ip1(n15648), .ip2(n15639), .op(n16778) );
  mux2_1 U14979 ( .ip1(n15653), .ip2(\ANSWER/mem[6][1][0] ), .s(n16778), .op(
        n3841) );
  nand2_1 U14980 ( .ip1(n15649), .ip2(n15639), .op(n16779) );
  mux2_1 U14981 ( .ip1(n15653), .ip2(\ANSWER/mem[6][2][0] ), .s(n16779), .op(
        n3840) );
  nand2_1 U14982 ( .ip1(n15650), .ip2(n15639), .op(n16780) );
  mux2_1 U14983 ( .ip1(n15644), .ip2(\ANSWER/mem[6][3][0] ), .s(n16780), .op(
        n3839) );
  nand2_1 U14984 ( .ip1(n15651), .ip2(n15639), .op(n16781) );
  mux2_1 U14985 ( .ip1(n15644), .ip2(\ANSWER/mem[6][4][0] ), .s(n16781), .op(
        n3838) );
  nand2_1 U14986 ( .ip1(n15652), .ip2(n15639), .op(n16782) );
  mux2_1 U14987 ( .ip1(n15659), .ip2(\ANSWER/mem[6][5][0] ), .s(n16782), .op(
        n3837) );
  nand2_1 U14988 ( .ip1(n15654), .ip2(n15639), .op(n16783) );
  mux2_1 U14989 ( .ip1(n15653), .ip2(\ANSWER/mem[6][6][0] ), .s(n16783), .op(
        n3836) );
  nand2_1 U14990 ( .ip1(n15655), .ip2(n15639), .op(n16784) );
  mux2_1 U14991 ( .ip1(n15653), .ip2(\ANSWER/mem[6][7][0] ), .s(n16784), .op(
        n3835) );
  nand2_1 U14992 ( .ip1(n15656), .ip2(n15639), .op(n16785) );
  mux2_1 U14993 ( .ip1(n15659), .ip2(\ANSWER/mem[6][8][0] ), .s(n16785), .op(
        n3834) );
  nand2_1 U14994 ( .ip1(n15658), .ip2(n15639), .op(n16786) );
  mux2_1 U14995 ( .ip1(n15653), .ip2(\ANSWER/mem[6][9][0] ), .s(n16786), .op(
        n3833) );
  nor4_1 U14996 ( .ip1(n15641), .ip2(n4366), .ip3(n17488), .ip4(n15640), .op(
        n15642) );
  nand2_1 U14997 ( .ip1(n15647), .ip2(n15642), .op(n16787) );
  mux2_1 U14998 ( .ip1(n15644), .ip2(\ANSWER/mem[7][0][0] ), .s(n16787), .op(
        n3832) );
  nand2_1 U14999 ( .ip1(n15648), .ip2(n15642), .op(n16788) );
  mux2_1 U15000 ( .ip1(n15644), .ip2(\ANSWER/mem[7][1][0] ), .s(n16788), .op(
        n3831) );
  nand2_1 U15001 ( .ip1(n15649), .ip2(n15642), .op(n16790) );
  mux2_1 U15002 ( .ip1(n15644), .ip2(\ANSWER/mem[7][2][0] ), .s(n16790), .op(
        n3830) );
  nand2_1 U15003 ( .ip1(n15650), .ip2(n15642), .op(n16791) );
  mux2_1 U15004 ( .ip1(n15644), .ip2(\ANSWER/mem[7][3][0] ), .s(n16791), .op(
        n3829) );
  nand2_1 U15005 ( .ip1(n15651), .ip2(n15642), .op(n16792) );
  mux2_1 U15006 ( .ip1(n15644), .ip2(\ANSWER/mem[7][4][0] ), .s(n16792), .op(
        n3828) );
  nand2_1 U15007 ( .ip1(n15652), .ip2(n15642), .op(n16793) );
  mux2_1 U15008 ( .ip1(n15644), .ip2(\ANSWER/mem[7][5][0] ), .s(n16793), .op(
        n3827) );
  nand2_1 U15009 ( .ip1(n15654), .ip2(n15642), .op(n16794) );
  mux2_1 U15010 ( .ip1(n15644), .ip2(\ANSWER/mem[7][6][0] ), .s(n16794), .op(
        n3826) );
  nand2_1 U15011 ( .ip1(n15655), .ip2(n15642), .op(n16795) );
  mux2_1 U15012 ( .ip1(n15644), .ip2(\ANSWER/mem[7][7][0] ), .s(n16795), .op(
        n3825) );
  nand2_1 U15013 ( .ip1(n15656), .ip2(n15642), .op(n16796) );
  mux2_1 U15014 ( .ip1(n15653), .ip2(\ANSWER/mem[7][8][0] ), .s(n16796), .op(
        n3824) );
  nand2_1 U15015 ( .ip1(n15658), .ip2(n15642), .op(n16797) );
  mux2_1 U15016 ( .ip1(n15659), .ip2(\ANSWER/mem[7][9][0] ), .s(n16797), .op(
        n3823) );
  nor3_1 U15017 ( .ip1(n18165), .ip2(n15643), .ip3(n15646), .op(n15645) );
  nand2_1 U15018 ( .ip1(n15647), .ip2(n15645), .op(n16798) );
  mux2_1 U15019 ( .ip1(n15653), .ip2(\ANSWER/mem[8][0][0] ), .s(n16798), .op(
        n3822) );
  nand2_1 U15020 ( .ip1(n15648), .ip2(n15645), .op(n16799) );
  mux2_1 U15021 ( .ip1(n15659), .ip2(\ANSWER/mem[8][1][0] ), .s(n16799), .op(
        n3821) );
  nand2_1 U15022 ( .ip1(n15649), .ip2(n15645), .op(n16800) );
  mux2_1 U15023 ( .ip1(n15659), .ip2(\ANSWER/mem[8][2][0] ), .s(n16800), .op(
        n3820) );
  nand2_1 U15024 ( .ip1(n15650), .ip2(n15645), .op(n16801) );
  mux2_1 U15025 ( .ip1(n15644), .ip2(\ANSWER/mem[8][3][0] ), .s(n16801), .op(
        n3819) );
  nand2_1 U15026 ( .ip1(n15651), .ip2(n15645), .op(n16803) );
  mux2_1 U15027 ( .ip1(n15659), .ip2(\ANSWER/mem[8][4][0] ), .s(n16803), .op(
        n3818) );
  nand2_1 U15028 ( .ip1(n15652), .ip2(n15645), .op(n16804) );
  mux2_1 U15029 ( .ip1(n15653), .ip2(\ANSWER/mem[8][5][0] ), .s(n16804), .op(
        n3817) );
  nand2_1 U15030 ( .ip1(n15654), .ip2(n15645), .op(n16805) );
  mux2_1 U15031 ( .ip1(n15644), .ip2(\ANSWER/mem[8][6][0] ), .s(n16805), .op(
        n3816) );
  nand2_1 U15032 ( .ip1(n15655), .ip2(n15645), .op(n16806) );
  mux2_1 U15033 ( .ip1(n15659), .ip2(\ANSWER/mem[8][7][0] ), .s(n16806), .op(
        n3815) );
  nand2_1 U15034 ( .ip1(n15656), .ip2(n15645), .op(n16807) );
  mux2_1 U15035 ( .ip1(n15653), .ip2(\ANSWER/mem[8][8][0] ), .s(n16807), .op(
        n3814) );
  nand2_1 U15036 ( .ip1(n15658), .ip2(n15645), .op(n16808) );
  mux2_1 U15037 ( .ip1(n15659), .ip2(\ANSWER/mem[8][9][0] ), .s(n16808), .op(
        n3813) );
  nor3_1 U15038 ( .ip1(n4362), .ip2(n18165), .ip3(n15646), .op(n15657) );
  nand2_1 U15039 ( .ip1(n15647), .ip2(n15657), .op(n16809) );
  mux2_1 U15040 ( .ip1(n15653), .ip2(\ANSWER/mem[9][0][0] ), .s(n16809), .op(
        n3812) );
  nand2_1 U15041 ( .ip1(n15648), .ip2(n15657), .op(n16810) );
  mux2_1 U15042 ( .ip1(n15653), .ip2(\ANSWER/mem[9][1][0] ), .s(n16810), .op(
        n3811) );
  nand2_1 U15043 ( .ip1(n15649), .ip2(n15657), .op(n16811) );
  mux2_1 U15044 ( .ip1(n15659), .ip2(\ANSWER/mem[9][2][0] ), .s(n16811), .op(
        n3810) );
  nand2_1 U15045 ( .ip1(n15650), .ip2(n15657), .op(n16812) );
  mux2_1 U15046 ( .ip1(n15653), .ip2(\ANSWER/mem[9][3][0] ), .s(n16812), .op(
        n3809) );
  nand2_1 U15047 ( .ip1(n15651), .ip2(n15657), .op(n16813) );
  mux2_1 U15048 ( .ip1(n15659), .ip2(\ANSWER/mem[9][4][0] ), .s(n16813), .op(
        n3808) );
  nand2_1 U15049 ( .ip1(n15652), .ip2(n15657), .op(n16814) );
  mux2_1 U15050 ( .ip1(n15653), .ip2(\ANSWER/mem[9][5][0] ), .s(n16814), .op(
        n3807) );
  nand2_1 U15051 ( .ip1(n15654), .ip2(n15657), .op(n16815) );
  mux2_1 U15052 ( .ip1(n15659), .ip2(\ANSWER/mem[9][6][0] ), .s(n16815), .op(
        n3806) );
  nand2_1 U15053 ( .ip1(n15655), .ip2(n15657), .op(n16816) );
  mux2_1 U15054 ( .ip1(n15659), .ip2(\ANSWER/mem[9][7][0] ), .s(n16816), .op(
        n3805) );
  nand2_1 U15055 ( .ip1(n15656), .ip2(n15657), .op(n16817) );
  mux2_1 U15056 ( .ip1(n15659), .ip2(\ANSWER/mem[9][8][0] ), .s(n16817), .op(
        n3804) );
  nand2_1 U15057 ( .ip1(n15658), .ip2(n15657), .op(n16818) );
  mux2_1 U15058 ( .ip1(n15659), .ip2(\ANSWER/mem[9][9][0] ), .s(n16818), .op(
        n3803) );
  fulladder U15059 ( .a(n15662), .b(n15661), .ci(n15660), .co(n15724), .s(
        n15711) );
  or2_1 U15060 ( .ip1(n15663), .ip2(n15664), .op(n15667) );
  or2_1 U15061 ( .ip1(n15665), .ip2(n15664), .op(n15666) );
  nand2_1 U15062 ( .ip1(n15667), .ip2(n15666), .op(n15768) );
  inv_1 U15063 ( .ip(rdata[1]), .op(n15746) );
  nand2_1 U15064 ( .ip1(m2DataIn[2]), .ip2(q_w2[8]), .op(n15749) );
  nor3_1 U15065 ( .ip1(n16222), .ip2(n16561), .ip3(n15749), .op(n15748) );
  inv_1 U15066 ( .ip(n15748), .op(n15670) );
  nand2_1 U15067 ( .ip1(m2DataIn[2]), .ip2(q_w2[7]), .op(n16191) );
  nand2_1 U15068 ( .ip1(m2DataIn[1]), .ip2(q_w2[8]), .op(n15668) );
  nand2_1 U15069 ( .ip1(n16191), .ip2(n15668), .op(n15669) );
  nand2_1 U15070 ( .ip1(n15670), .ip2(n15669), .op(n15745) );
  mux2_1 U15071 ( .ip1(rdata[1]), .ip2(n15746), .s(n15745), .op(n15767) );
  or2_1 U15072 ( .ip1(n15671), .ip2(n15672), .op(n15675) );
  or2_1 U15073 ( .ip1(n15673), .ip2(n15672), .op(n15674) );
  nand2_1 U15074 ( .ip1(n15675), .ip2(n15674), .op(n15766) );
  inv_1 U15075 ( .ip(n15676), .op(n15772) );
  nor4_1 U15076 ( .ip1(n16309), .ip2(n16222), .ip3(n16538), .ip4(n16561), .op(
        n15678) );
  nor2_1 U15077 ( .ip1(n15678), .ip2(n15677), .op(n15683) );
  nor3_1 U15078 ( .ip1(n16550), .ip2(n16177), .ip3(n15704), .op(n15761) );
  nor2_1 U15079 ( .ip1(n16273), .ip2(n16177), .op(n15679) );
  or2_1 U15080 ( .ip1(q_w2[2]), .ip2(n15679), .op(n15681) );
  or2_1 U15081 ( .ip1(m2DataIn[7]), .ip2(n15679), .op(n15680) );
  nand2_1 U15082 ( .ip1(n15681), .ip2(n15680), .op(n15682) );
  or2_1 U15083 ( .ip1(n15761), .ip2(n15682), .op(n15684) );
  nor2_1 U15084 ( .ip1(n15683), .ip2(n15684), .op(n15760) );
  or2_1 U15085 ( .ip1(n15683), .ip2(n15760), .op(n15686) );
  or2_1 U15086 ( .ip1(n15684), .ip2(n15760), .op(n15685) );
  nand2_1 U15087 ( .ip1(n15686), .ip2(n15685), .op(n15771) );
  fulladder U15088 ( .a(n15689), .b(n15688), .ci(n15687), .co(n15770), .s(
        n15660) );
  inv_1 U15089 ( .ip(n15690), .op(n15721) );
  inv_1 U15090 ( .ip(q_w2[9]), .op(n16552) );
  nor2_1 U15091 ( .ip1(n16369), .ip2(n16552), .op(n15879) );
  nand2_1 U15092 ( .ip1(n15879), .ip2(n15691), .op(n15743) );
  inv_1 U15093 ( .ip(n15743), .op(n15696) );
  nor2_1 U15094 ( .ip1(n16145), .ip2(n16552), .op(n15692) );
  or2_1 U15095 ( .ip1(q_w2[6]), .ip2(n15692), .op(n15694) );
  or2_1 U15096 ( .ip1(m2DataIn[3]), .ip2(n15692), .op(n15693) );
  nand2_1 U15097 ( .ip1(n15694), .ip2(n15693), .op(n15695) );
  nor2_1 U15098 ( .ip1(n15696), .ip2(n15695), .op(n15741) );
  nand2_1 U15099 ( .ip1(m2DataIn[9]), .ip2(q_w2[0]), .op(n15697) );
  xor2_1 U15100 ( .ip1(n15741), .ip2(n15697), .op(n15758) );
  nor2_1 U15101 ( .ip1(n16624), .ip2(n16144), .op(n15702) );
  nand2_1 U15102 ( .ip1(m2DataIn[5]), .ip2(q_w2[5]), .op(n15733) );
  nor3_1 U15103 ( .ip1(n16445), .ip2(n16447), .ip3(n15733), .op(n15755) );
  inv_1 U15104 ( .ip(n15755), .op(n15701) );
  nand2_1 U15105 ( .ip1(m2DataIn[4]), .ip2(q_w2[5]), .op(n15699) );
  nand2_1 U15106 ( .ip1(n15699), .ip2(n15698), .op(n15700) );
  nand2_1 U15107 ( .ip1(n15701), .ip2(n15700), .op(n15753) );
  xor2_1 U15108 ( .ip1(n15702), .ip2(n15753), .op(n15757) );
  fulladder U15109 ( .a(n15705), .b(n15704), .ci(n15703), .co(n15756), .s(
        n15707) );
  fulladder U15110 ( .a(n15708), .b(n15707), .ci(n15706), .co(n15719), .s(
        n15605) );
  inv_1 U15111 ( .ip(n15709), .op(n15723) );
  fulladder U15112 ( .a(n15712), .b(n15711), .ci(n15710), .co(n15722), .s(
        n15623) );
  inv_1 U15113 ( .ip(\SIGMOID/lut_out [1]), .op(n15714) );
  inv_1 U15114 ( .ip(\SIGMOID/sign_bit ), .op(n16164) );
  nand2_1 U15115 ( .ip1(\SIGMOID/N64 ), .ip2(n16164), .op(n15713) );
  mux2_1 U15116 ( .ip1(n15714), .ip2(\SIGMOID/lut_out [1]), .s(n15713), .op(
        n17039) );
  mux2_1 U15117 ( .ip1(n15715), .ip2(n17039), .s(n16714), .op(n15716) );
  mux2_1 U15118 ( .ip1(n15716), .ip2(\ANSWER/mem[0][0][1] ), .s(n16717), .op(
        n3802) );
  buf_1 U15119 ( .ip(n15716), .op(n15718) );
  mux2_1 U15120 ( .ip1(n15718), .ip2(\ANSWER/mem[0][1][1] ), .s(n16718), .op(
        n3801) );
  mux2_1 U15121 ( .ip1(n15718), .ip2(\ANSWER/mem[0][2][1] ), .s(n16719), .op(
        n3800) );
  buf_1 U15122 ( .ip(n15716), .op(n15717) );
  mux2_1 U15123 ( .ip1(n15717), .ip2(\ANSWER/mem[0][3][1] ), .s(n16720), .op(
        n3799) );
  mux2_1 U15124 ( .ip1(n15718), .ip2(\ANSWER/mem[0][4][1] ), .s(n16721), .op(
        n3798) );
  mux2_1 U15125 ( .ip1(n15717), .ip2(\ANSWER/mem[0][5][1] ), .s(n16722), .op(
        n3797) );
  mux2_1 U15126 ( .ip1(n15718), .ip2(\ANSWER/mem[0][6][1] ), .s(n16723), .op(
        n3796) );
  mux2_1 U15127 ( .ip1(n15717), .ip2(\ANSWER/mem[0][7][1] ), .s(n16724), .op(
        n3795) );
  mux2_1 U15128 ( .ip1(n15718), .ip2(\ANSWER/mem[0][8][1] ), .s(n16725), .op(
        n3794) );
  mux2_1 U15129 ( .ip1(n15717), .ip2(\ANSWER/mem[0][9][1] ), .s(n16726), .op(
        n3793) );
  mux2_1 U15130 ( .ip1(n15718), .ip2(\ANSWER/mem[1][0][1] ), .s(n16727), .op(
        n3792) );
  mux2_1 U15131 ( .ip1(n15717), .ip2(\ANSWER/mem[1][1][1] ), .s(n16728), .op(
        n3791) );
  mux2_1 U15132 ( .ip1(n15716), .ip2(\ANSWER/mem[1][2][1] ), .s(n16729), .op(
        n3790) );
  mux2_1 U15133 ( .ip1(n15716), .ip2(\ANSWER/mem[1][3][1] ), .s(n16730), .op(
        n3789) );
  mux2_1 U15134 ( .ip1(n15716), .ip2(\ANSWER/mem[1][4][1] ), .s(n16731), .op(
        n3788) );
  mux2_1 U15135 ( .ip1(n15716), .ip2(\ANSWER/mem[1][5][1] ), .s(n16732), .op(
        n3787) );
  mux2_1 U15136 ( .ip1(n15718), .ip2(\ANSWER/mem[1][6][1] ), .s(n16733), .op(
        n3786) );
  mux2_1 U15137 ( .ip1(n15718), .ip2(\ANSWER/mem[1][7][1] ), .s(n16734), .op(
        n3785) );
  mux2_1 U15138 ( .ip1(n15717), .ip2(\ANSWER/mem[1][8][1] ), .s(n16735), .op(
        n3784) );
  mux2_1 U15139 ( .ip1(n15717), .ip2(\ANSWER/mem[1][9][1] ), .s(n16736), .op(
        n3783) );
  mux2_1 U15140 ( .ip1(n15718), .ip2(\ANSWER/mem[2][0][1] ), .s(n16737), .op(
        n3782) );
  mux2_1 U15141 ( .ip1(n15716), .ip2(\ANSWER/mem[2][1][1] ), .s(n16738), .op(
        n3781) );
  mux2_1 U15142 ( .ip1(n15716), .ip2(\ANSWER/mem[2][2][1] ), .s(n16739), .op(
        n3780) );
  mux2_1 U15143 ( .ip1(n15716), .ip2(\ANSWER/mem[2][3][1] ), .s(n16740), .op(
        n3779) );
  mux2_1 U15144 ( .ip1(n15716), .ip2(\ANSWER/mem[2][4][1] ), .s(n16741), .op(
        n3778) );
  mux2_1 U15145 ( .ip1(n15716), .ip2(\ANSWER/mem[2][5][1] ), .s(n16742), .op(
        n3777) );
  mux2_1 U15146 ( .ip1(n15716), .ip2(\ANSWER/mem[2][6][1] ), .s(n16743), .op(
        n3776) );
  mux2_1 U15147 ( .ip1(n15716), .ip2(\ANSWER/mem[2][7][1] ), .s(n16744), .op(
        n3775) );
  mux2_1 U15148 ( .ip1(n15716), .ip2(\ANSWER/mem[2][8][1] ), .s(n16745), .op(
        n3774) );
  mux2_1 U15149 ( .ip1(n15716), .ip2(\ANSWER/mem[2][9][1] ), .s(n16746), .op(
        n3773) );
  mux2_1 U15150 ( .ip1(n15716), .ip2(\ANSWER/mem[3][0][1] ), .s(n16747), .op(
        n3772) );
  mux2_1 U15151 ( .ip1(n15716), .ip2(\ANSWER/mem[3][1][1] ), .s(n16748), .op(
        n3771) );
  mux2_1 U15152 ( .ip1(n15716), .ip2(\ANSWER/mem[3][2][1] ), .s(n16749), .op(
        n3770) );
  mux2_1 U15153 ( .ip1(n15716), .ip2(\ANSWER/mem[3][3][1] ), .s(n16750), .op(
        n3769) );
  mux2_1 U15154 ( .ip1(n15716), .ip2(\ANSWER/mem[3][4][1] ), .s(n16751), .op(
        n3768) );
  mux2_1 U15155 ( .ip1(n15716), .ip2(\ANSWER/mem[3][5][1] ), .s(n16752), .op(
        n3767) );
  mux2_1 U15156 ( .ip1(n15716), .ip2(\ANSWER/mem[3][6][1] ), .s(n16753), .op(
        n3766) );
  mux2_1 U15157 ( .ip1(n15716), .ip2(\ANSWER/mem[3][7][1] ), .s(n16754), .op(
        n3765) );
  mux2_1 U15158 ( .ip1(n15716), .ip2(\ANSWER/mem[3][8][1] ), .s(n16755), .op(
        n3764) );
  mux2_1 U15159 ( .ip1(n15716), .ip2(\ANSWER/mem[3][9][1] ), .s(n16756), .op(
        n3763) );
  mux2_1 U15160 ( .ip1(n15717), .ip2(\ANSWER/mem[4][0][1] ), .s(n16757), .op(
        n3762) );
  mux2_1 U15161 ( .ip1(n15718), .ip2(\ANSWER/mem[4][1][1] ), .s(n16758), .op(
        n3761) );
  mux2_1 U15162 ( .ip1(n15717), .ip2(\ANSWER/mem[4][2][1] ), .s(n16759), .op(
        n3760) );
  mux2_1 U15163 ( .ip1(n15717), .ip2(\ANSWER/mem[4][3][1] ), .s(n16760), .op(
        n3759) );
  mux2_1 U15164 ( .ip1(n15716), .ip2(\ANSWER/mem[4][4][1] ), .s(n16761), .op(
        n3758) );
  mux2_1 U15165 ( .ip1(n15716), .ip2(\ANSWER/mem[4][5][1] ), .s(n16762), .op(
        n3757) );
  mux2_1 U15166 ( .ip1(n15716), .ip2(\ANSWER/mem[4][6][1] ), .s(n16763), .op(
        n3756) );
  mux2_1 U15167 ( .ip1(n15716), .ip2(\ANSWER/mem[4][7][1] ), .s(n16764), .op(
        n3755) );
  mux2_1 U15168 ( .ip1(n15718), .ip2(\ANSWER/mem[4][8][1] ), .s(n16765), .op(
        n3754) );
  mux2_1 U15169 ( .ip1(n15718), .ip2(\ANSWER/mem[4][9][1] ), .s(n16766), .op(
        n3753) );
  mux2_1 U15170 ( .ip1(n15718), .ip2(\ANSWER/mem[5][0][1] ), .s(n16767), .op(
        n3752) );
  mux2_1 U15171 ( .ip1(n15718), .ip2(\ANSWER/mem[5][1][1] ), .s(n16768), .op(
        n3751) );
  mux2_1 U15172 ( .ip1(n15717), .ip2(\ANSWER/mem[5][2][1] ), .s(n16769), .op(
        n3750) );
  mux2_1 U15173 ( .ip1(n15716), .ip2(\ANSWER/mem[5][3][1] ), .s(n16770), .op(
        n3749) );
  mux2_1 U15174 ( .ip1(n15718), .ip2(\ANSWER/mem[5][4][1] ), .s(n16771), .op(
        n3748) );
  mux2_1 U15175 ( .ip1(n15717), .ip2(\ANSWER/mem[5][5][1] ), .s(n16772), .op(
        n3747) );
  mux2_1 U15176 ( .ip1(n15716), .ip2(\ANSWER/mem[5][6][1] ), .s(n16773), .op(
        n3746) );
  mux2_1 U15177 ( .ip1(n15718), .ip2(\ANSWER/mem[5][7][1] ), .s(n16774), .op(
        n3745) );
  mux2_1 U15178 ( .ip1(n15717), .ip2(\ANSWER/mem[5][8][1] ), .s(n16775), .op(
        n3744) );
  mux2_1 U15179 ( .ip1(n15716), .ip2(\ANSWER/mem[5][9][1] ), .s(n16776), .op(
        n3743) );
  mux2_1 U15180 ( .ip1(n15718), .ip2(\ANSWER/mem[6][0][1] ), .s(n16777), .op(
        n3742) );
  mux2_1 U15181 ( .ip1(n15717), .ip2(\ANSWER/mem[6][1][1] ), .s(n16778), .op(
        n3741) );
  mux2_1 U15182 ( .ip1(n15718), .ip2(\ANSWER/mem[6][2][1] ), .s(n16779), .op(
        n3740) );
  mux2_1 U15183 ( .ip1(n15718), .ip2(\ANSWER/mem[6][3][1] ), .s(n16780), .op(
        n3739) );
  mux2_1 U15184 ( .ip1(n15718), .ip2(\ANSWER/mem[6][4][1] ), .s(n16781), .op(
        n3738) );
  mux2_1 U15185 ( .ip1(n15718), .ip2(\ANSWER/mem[6][5][1] ), .s(n16782), .op(
        n3737) );
  mux2_1 U15186 ( .ip1(n15718), .ip2(\ANSWER/mem[6][6][1] ), .s(n16783), .op(
        n3736) );
  mux2_1 U15187 ( .ip1(n15716), .ip2(\ANSWER/mem[6][7][1] ), .s(n16784), .op(
        n3735) );
  mux2_1 U15188 ( .ip1(n15717), .ip2(\ANSWER/mem[6][8][1] ), .s(n16785), .op(
        n3734) );
  mux2_1 U15189 ( .ip1(n15718), .ip2(\ANSWER/mem[6][9][1] ), .s(n16786), .op(
        n3733) );
  mux2_1 U15190 ( .ip1(n15716), .ip2(\ANSWER/mem[7][0][1] ), .s(n16787), .op(
        n3732) );
  mux2_1 U15191 ( .ip1(n15718), .ip2(\ANSWER/mem[7][1][1] ), .s(n16788), .op(
        n3731) );
  mux2_1 U15192 ( .ip1(n15716), .ip2(\ANSWER/mem[7][2][1] ), .s(n16790), .op(
        n3730) );
  mux2_1 U15193 ( .ip1(n15718), .ip2(\ANSWER/mem[7][3][1] ), .s(n16791), .op(
        n3729) );
  mux2_1 U15194 ( .ip1(n15716), .ip2(\ANSWER/mem[7][4][1] ), .s(n16792), .op(
        n3728) );
  mux2_1 U15195 ( .ip1(n15717), .ip2(\ANSWER/mem[7][5][1] ), .s(n16793), .op(
        n3727) );
  mux2_1 U15196 ( .ip1(n15717), .ip2(\ANSWER/mem[7][6][1] ), .s(n16794), .op(
        n3726) );
  mux2_1 U15197 ( .ip1(n15716), .ip2(\ANSWER/mem[7][7][1] ), .s(n16795), .op(
        n3725) );
  mux2_1 U15198 ( .ip1(n15716), .ip2(\ANSWER/mem[7][8][1] ), .s(n16796), .op(
        n3724) );
  mux2_1 U15199 ( .ip1(n15716), .ip2(\ANSWER/mem[7][9][1] ), .s(n16797), .op(
        n3723) );
  mux2_1 U15200 ( .ip1(n15717), .ip2(\ANSWER/mem[8][0][1] ), .s(n16798), .op(
        n3722) );
  mux2_1 U15201 ( .ip1(n15718), .ip2(\ANSWER/mem[8][1][1] ), .s(n16799), .op(
        n3721) );
  mux2_1 U15202 ( .ip1(n15717), .ip2(\ANSWER/mem[8][2][1] ), .s(n16800), .op(
        n3720) );
  mux2_1 U15203 ( .ip1(n15718), .ip2(\ANSWER/mem[8][3][1] ), .s(n16801), .op(
        n3719) );
  mux2_1 U15204 ( .ip1(n15717), .ip2(\ANSWER/mem[8][4][1] ), .s(n16803), .op(
        n3718) );
  mux2_1 U15205 ( .ip1(n15717), .ip2(\ANSWER/mem[8][5][1] ), .s(n16804), .op(
        n3717) );
  mux2_1 U15206 ( .ip1(n15717), .ip2(\ANSWER/mem[8][6][1] ), .s(n16805), .op(
        n3716) );
  mux2_1 U15207 ( .ip1(n15717), .ip2(\ANSWER/mem[8][7][1] ), .s(n16806), .op(
        n3715) );
  mux2_1 U15208 ( .ip1(n15717), .ip2(\ANSWER/mem[8][8][1] ), .s(n16807), .op(
        n3714) );
  mux2_1 U15209 ( .ip1(n15717), .ip2(\ANSWER/mem[8][9][1] ), .s(n16808), .op(
        n3713) );
  mux2_1 U15210 ( .ip1(n15717), .ip2(\ANSWER/mem[9][0][1] ), .s(n16809), .op(
        n3712) );
  mux2_1 U15211 ( .ip1(n15717), .ip2(\ANSWER/mem[9][1][1] ), .s(n16810), .op(
        n3711) );
  mux2_1 U15212 ( .ip1(n15717), .ip2(\ANSWER/mem[9][2][1] ), .s(n16811), .op(
        n3710) );
  mux2_1 U15213 ( .ip1(n15717), .ip2(\ANSWER/mem[9][3][1] ), .s(n16812), .op(
        n3709) );
  mux2_1 U15214 ( .ip1(n15717), .ip2(\ANSWER/mem[9][4][1] ), .s(n16813), .op(
        n3708) );
  mux2_1 U15215 ( .ip1(n15717), .ip2(\ANSWER/mem[9][5][1] ), .s(n16814), .op(
        n3707) );
  mux2_1 U15216 ( .ip1(n15718), .ip2(\ANSWER/mem[9][6][1] ), .s(n16815), .op(
        n3706) );
  mux2_1 U15217 ( .ip1(n15718), .ip2(\ANSWER/mem[9][7][1] ), .s(n16816), .op(
        n3705) );
  mux2_1 U15218 ( .ip1(n15718), .ip2(\ANSWER/mem[9][8][1] ), .s(n16817), .op(
        n3704) );
  mux2_1 U15219 ( .ip1(n15718), .ip2(\ANSWER/mem[9][9][1] ), .s(n16818), .op(
        n3703) );
  fulladder U15220 ( .a(n15721), .b(n15720), .ci(n15719), .co(n15786), .s(
        n15709) );
  inv_1 U15221 ( .ip(n15786), .op(n15776) );
  fulladder U15222 ( .a(n15724), .b(n15723), .ci(n15722), .co(n15774), .s(
        n15715) );
  nand2_1 U15223 ( .ip1(m2DataIn[7]), .ip2(q_w2[4]), .op(n15803) );
  nor3_1 U15224 ( .ip1(n16273), .ip2(n16177), .ip3(n15803), .op(n15820) );
  inv_1 U15225 ( .ip(n15820), .op(n15728) );
  nand2_1 U15226 ( .ip1(m2DataIn[7]), .ip2(q_w2[3]), .op(n15726) );
  nand2_1 U15227 ( .ip1(m2DataIn[6]), .ip2(q_w2[4]), .op(n15725) );
  nand2_1 U15228 ( .ip1(n15726), .ip2(n15725), .op(n15727) );
  nand2_1 U15229 ( .ip1(n15728), .ip2(n15727), .op(n15729) );
  nor3_1 U15230 ( .ip1(n16624), .ip2(n16308), .ip3(n15729), .op(n15819) );
  or2_1 U15231 ( .ip1(n15729), .ip2(n15819), .op(n15732) );
  nand2_1 U15232 ( .ip1(m2DataIn[8]), .ip2(q_w2[2]), .op(n15730) );
  or2_1 U15233 ( .ip1(n15730), .ip2(n15819), .op(n15731) );
  nand2_1 U15234 ( .ip1(n15732), .ip2(n15731), .op(n15834) );
  nand2_1 U15235 ( .ip1(m2DataIn[5]), .ip2(q_w2[6]), .op(n15799) );
  nor3_1 U15236 ( .ip1(n16445), .ip2(n16497), .ip3(n15799), .op(n15813) );
  inv_1 U15237 ( .ip(n15813), .op(n15736) );
  nand2_1 U15238 ( .ip1(m2DataIn[4]), .ip2(q_w2[6]), .op(n15734) );
  nand2_1 U15239 ( .ip1(n15734), .ip2(n15733), .op(n15735) );
  nand2_1 U15240 ( .ip1(n15736), .ip2(n15735), .op(n15737) );
  nor3_1 U15241 ( .ip1(n16690), .ip2(n16144), .ip3(n15737), .op(n15812) );
  or2_1 U15242 ( .ip1(n15737), .ip2(n15812), .op(n15740) );
  nand2_1 U15243 ( .ip1(m2DataIn[9]), .ip2(q_w2[1]), .op(n15738) );
  or2_1 U15244 ( .ip1(n15738), .ip2(n15812), .op(n15739) );
  nand2_1 U15245 ( .ip1(n15740), .ip2(n15739), .op(n15833) );
  nand3_1 U15246 ( .ip1(m2DataIn[9]), .ip2(q_w2[0]), .ip3(n15741), .op(n15742)
         );
  nand2_1 U15247 ( .ip1(n15743), .ip2(n15742), .op(n15832) );
  inv_1 U15248 ( .ip(n15744), .op(n15841) );
  nor2_1 U15249 ( .ip1(n15746), .ip2(n15745), .op(n15747) );
  nor2_1 U15250 ( .ip1(n15748), .ip2(n15747), .op(n15838) );
  inv_1 U15251 ( .ip(rdata[2]), .op(n15825) );
  nand2_1 U15252 ( .ip1(m2DataIn[2]), .ip2(q_w2[9]), .op(n15814) );
  nor3_1 U15253 ( .ip1(n16222), .ip2(n16596), .ip3(n15814), .op(n15827) );
  inv_1 U15254 ( .ip(n15827), .op(n15752) );
  nand2_1 U15255 ( .ip1(m2DataIn[1]), .ip2(q_w2[9]), .op(n15750) );
  nand2_1 U15256 ( .ip1(n15750), .ip2(n15749), .op(n15751) );
  nand2_1 U15257 ( .ip1(n15752), .ip2(n15751), .op(n15824) );
  mux2_1 U15258 ( .ip1(rdata[2]), .ip2(n15825), .s(n15824), .op(n15837) );
  nor3_1 U15259 ( .ip1(n16624), .ip2(n16144), .ip3(n15753), .op(n15754) );
  nor2_1 U15260 ( .ip1(n15755), .ip2(n15754), .op(n15836) );
  fulladder U15261 ( .a(n15758), .b(n15757), .ci(n15756), .co(n15839), .s(
        n15720) );
  inv_1 U15262 ( .ip(n15759), .op(n15785) );
  nor2_1 U15263 ( .ip1(n15761), .ip2(n15760), .op(n15823) );
  nor2_1 U15264 ( .ip1(n16600), .ip2(n15973), .op(n15765) );
  inv_1 U15265 ( .ip(q_w2[10]), .op(n16622) );
  nor2_1 U15266 ( .ip1(n16369), .ip2(n16622), .op(n15968) );
  nand3_1 U15267 ( .ip1(m2DataIn[0]), .ip2(q_w2[7]), .ip3(n15968), .op(n15828)
         );
  nand2_1 U15268 ( .ip1(m2DataIn[0]), .ip2(q_w2[10]), .op(n15763) );
  nand2_1 U15269 ( .ip1(n15763), .ip2(n15762), .op(n15764) );
  nand2_1 U15270 ( .ip1(n15828), .ip2(n15764), .op(n15829) );
  xor2_1 U15271 ( .ip1(n15765), .ip2(n15829), .op(n15822) );
  fulladder U15272 ( .a(n15768), .b(n15767), .ci(n15766), .co(n15821), .s(
        n15676) );
  inv_1 U15273 ( .ip(n15769), .op(n15784) );
  fulladder U15274 ( .a(n15772), .b(n15771), .ci(n15770), .co(n15783), .s(
        n15690) );
  and2_1 U15275 ( .ip1(n15774), .ip2(n15773), .op(n15789) );
  nor2_1 U15276 ( .ip1(n15774), .ip2(n15773), .op(n15787) );
  nor2_1 U15277 ( .ip1(n15789), .ip2(n15787), .op(n15775) );
  mux2_1 U15278 ( .ip1(n15776), .ip2(n15786), .s(n15775), .op(n15779) );
  nor2_1 U15279 ( .ip1(\SIGMOID/lut_out [1]), .ip2(\SIGMOID/N64 ), .op(n15777)
         );
  nor2_1 U15280 ( .ip1(\SIGMOID/sign_bit ), .ip2(n15777), .op(n15778) );
  xor2_1 U15281 ( .ip1(\SIGMOID/lut_out [2]), .ip2(n15778), .op(n17071) );
  mux2_1 U15282 ( .ip1(n15779), .ip2(n17071), .s(n16714), .op(n15781) );
  buf_1 U15283 ( .ip(n15781), .op(n15780) );
  mux2_1 U15284 ( .ip1(n15780), .ip2(\ANSWER/mem[0][0][2] ), .s(n16717), .op(
        n3702) );
  mux2_1 U15285 ( .ip1(n15780), .ip2(\ANSWER/mem[0][1][2] ), .s(n16718), .op(
        n3701) );
  mux2_1 U15286 ( .ip1(n15780), .ip2(\ANSWER/mem[0][2][2] ), .s(n16719), .op(
        n3700) );
  mux2_1 U15287 ( .ip1(n15780), .ip2(\ANSWER/mem[0][3][2] ), .s(n16720), .op(
        n3699) );
  mux2_1 U15288 ( .ip1(n15780), .ip2(\ANSWER/mem[0][4][2] ), .s(n16721), .op(
        n3698) );
  mux2_1 U15289 ( .ip1(n15780), .ip2(\ANSWER/mem[0][5][2] ), .s(n16722), .op(
        n3697) );
  mux2_1 U15290 ( .ip1(n15780), .ip2(\ANSWER/mem[0][6][2] ), .s(n16723), .op(
        n3696) );
  mux2_1 U15291 ( .ip1(n15780), .ip2(\ANSWER/mem[0][7][2] ), .s(n16724), .op(
        n3695) );
  mux2_1 U15292 ( .ip1(n15780), .ip2(\ANSWER/mem[0][8][2] ), .s(n16725), .op(
        n3694) );
  mux2_1 U15293 ( .ip1(n15780), .ip2(\ANSWER/mem[0][9][2] ), .s(n16726), .op(
        n3693) );
  mux2_1 U15294 ( .ip1(n15780), .ip2(\ANSWER/mem[1][0][2] ), .s(n16727), .op(
        n3692) );
  mux2_1 U15295 ( .ip1(n15780), .ip2(\ANSWER/mem[1][1][2] ), .s(n16728), .op(
        n3691) );
  mux2_1 U15296 ( .ip1(n15780), .ip2(\ANSWER/mem[1][2][2] ), .s(n16729), .op(
        n3690) );
  mux2_1 U15297 ( .ip1(n15780), .ip2(\ANSWER/mem[1][3][2] ), .s(n16730), .op(
        n3689) );
  mux2_1 U15298 ( .ip1(n15780), .ip2(\ANSWER/mem[1][4][2] ), .s(n16731), .op(
        n3688) );
  mux2_1 U15299 ( .ip1(n15780), .ip2(\ANSWER/mem[1][5][2] ), .s(n16732), .op(
        n3687) );
  mux2_1 U15300 ( .ip1(n15780), .ip2(\ANSWER/mem[1][6][2] ), .s(n16733), .op(
        n3686) );
  mux2_1 U15301 ( .ip1(n15780), .ip2(\ANSWER/mem[1][7][2] ), .s(n16734), .op(
        n3685) );
  mux2_1 U15302 ( .ip1(n15780), .ip2(\ANSWER/mem[1][8][2] ), .s(n16735), .op(
        n3684) );
  mux2_1 U15303 ( .ip1(n15780), .ip2(\ANSWER/mem[1][9][2] ), .s(n16736), .op(
        n3683) );
  mux2_1 U15304 ( .ip1(n15780), .ip2(\ANSWER/mem[2][0][2] ), .s(n16737), .op(
        n3682) );
  mux2_1 U15305 ( .ip1(n15780), .ip2(\ANSWER/mem[2][1][2] ), .s(n16738), .op(
        n3681) );
  mux2_1 U15306 ( .ip1(n15780), .ip2(\ANSWER/mem[2][2][2] ), .s(n16739), .op(
        n3680) );
  mux2_1 U15307 ( .ip1(n15780), .ip2(\ANSWER/mem[2][3][2] ), .s(n16740), .op(
        n3679) );
  mux2_1 U15308 ( .ip1(n15780), .ip2(\ANSWER/mem[2][4][2] ), .s(n16741), .op(
        n3678) );
  mux2_1 U15309 ( .ip1(n15780), .ip2(\ANSWER/mem[2][5][2] ), .s(n16742), .op(
        n3677) );
  mux2_1 U15310 ( .ip1(n15780), .ip2(\ANSWER/mem[2][6][2] ), .s(n16743), .op(
        n3676) );
  mux2_1 U15311 ( .ip1(n15780), .ip2(\ANSWER/mem[2][7][2] ), .s(n16744), .op(
        n3675) );
  mux2_1 U15312 ( .ip1(n15780), .ip2(\ANSWER/mem[2][8][2] ), .s(n16745), .op(
        n3674) );
  mux2_1 U15313 ( .ip1(n15780), .ip2(\ANSWER/mem[2][9][2] ), .s(n16746), .op(
        n3673) );
  mux2_1 U15314 ( .ip1(n15780), .ip2(\ANSWER/mem[3][0][2] ), .s(n16747), .op(
        n3672) );
  mux2_1 U15315 ( .ip1(n15780), .ip2(\ANSWER/mem[3][1][2] ), .s(n16748), .op(
        n3671) );
  mux2_1 U15316 ( .ip1(n15780), .ip2(\ANSWER/mem[3][2][2] ), .s(n16749), .op(
        n3670) );
  mux2_1 U15317 ( .ip1(n15780), .ip2(\ANSWER/mem[3][3][2] ), .s(n16750), .op(
        n3669) );
  mux2_1 U15318 ( .ip1(n15780), .ip2(\ANSWER/mem[3][4][2] ), .s(n16751), .op(
        n3668) );
  mux2_1 U15319 ( .ip1(n15780), .ip2(\ANSWER/mem[3][5][2] ), .s(n16752), .op(
        n3667) );
  mux2_1 U15320 ( .ip1(n15782), .ip2(\ANSWER/mem[3][6][2] ), .s(n16753), .op(
        n3666) );
  mux2_1 U15321 ( .ip1(n15782), .ip2(\ANSWER/mem[3][7][2] ), .s(n16754), .op(
        n3665) );
  mux2_1 U15322 ( .ip1(n15782), .ip2(\ANSWER/mem[3][8][2] ), .s(n16755), .op(
        n3664) );
  mux2_1 U15323 ( .ip1(n15782), .ip2(\ANSWER/mem[3][9][2] ), .s(n16756), .op(
        n3663) );
  mux2_1 U15324 ( .ip1(n15781), .ip2(\ANSWER/mem[4][0][2] ), .s(n16757), .op(
        n3662) );
  mux2_1 U15325 ( .ip1(n15781), .ip2(\ANSWER/mem[4][1][2] ), .s(n16758), .op(
        n3661) );
  mux2_1 U15326 ( .ip1(n15781), .ip2(\ANSWER/mem[4][2][2] ), .s(n16759), .op(
        n3660) );
  mux2_1 U15327 ( .ip1(n15781), .ip2(\ANSWER/mem[4][3][2] ), .s(n16760), .op(
        n3659) );
  mux2_1 U15328 ( .ip1(n15782), .ip2(\ANSWER/mem[4][4][2] ), .s(n16761), .op(
        n3658) );
  mux2_1 U15329 ( .ip1(n15782), .ip2(\ANSWER/mem[4][5][2] ), .s(n16762), .op(
        n3657) );
  mux2_1 U15330 ( .ip1(n15782), .ip2(\ANSWER/mem[4][6][2] ), .s(n16763), .op(
        n3656) );
  mux2_1 U15331 ( .ip1(n15782), .ip2(\ANSWER/mem[4][7][2] ), .s(n16764), .op(
        n3655) );
  mux2_1 U15332 ( .ip1(n15782), .ip2(\ANSWER/mem[4][8][2] ), .s(n16765), .op(
        n3654) );
  mux2_1 U15333 ( .ip1(n15782), .ip2(\ANSWER/mem[4][9][2] ), .s(n16766), .op(
        n3653) );
  mux2_1 U15334 ( .ip1(n15782), .ip2(\ANSWER/mem[5][0][2] ), .s(n16767), .op(
        n3652) );
  mux2_1 U15335 ( .ip1(n15781), .ip2(\ANSWER/mem[5][1][2] ), .s(n16768), .op(
        n3651) );
  mux2_1 U15336 ( .ip1(n15782), .ip2(\ANSWER/mem[5][2][2] ), .s(n16769), .op(
        n3650) );
  mux2_1 U15337 ( .ip1(n15781), .ip2(\ANSWER/mem[5][3][2] ), .s(n16770), .op(
        n3649) );
  mux2_1 U15338 ( .ip1(n15782), .ip2(\ANSWER/mem[5][4][2] ), .s(n16771), .op(
        n3648) );
  mux2_1 U15339 ( .ip1(n15781), .ip2(\ANSWER/mem[5][5][2] ), .s(n16772), .op(
        n3647) );
  mux2_1 U15340 ( .ip1(n15781), .ip2(\ANSWER/mem[5][6][2] ), .s(n16773), .op(
        n3646) );
  mux2_1 U15341 ( .ip1(n15781), .ip2(\ANSWER/mem[5][7][2] ), .s(n16774), .op(
        n3645) );
  mux2_1 U15342 ( .ip1(n15781), .ip2(\ANSWER/mem[5][8][2] ), .s(n16775), .op(
        n3644) );
  mux2_1 U15343 ( .ip1(n15781), .ip2(\ANSWER/mem[5][9][2] ), .s(n16776), .op(
        n3643) );
  mux2_1 U15344 ( .ip1(n15781), .ip2(\ANSWER/mem[6][0][2] ), .s(n16777), .op(
        n3642) );
  mux2_1 U15345 ( .ip1(n15781), .ip2(\ANSWER/mem[6][1][2] ), .s(n16778), .op(
        n3641) );
  mux2_1 U15346 ( .ip1(n15781), .ip2(\ANSWER/mem[6][2][2] ), .s(n16779), .op(
        n3640) );
  mux2_1 U15347 ( .ip1(n15781), .ip2(\ANSWER/mem[6][3][2] ), .s(n16780), .op(
        n3639) );
  mux2_1 U15348 ( .ip1(n15781), .ip2(\ANSWER/mem[6][4][2] ), .s(n16781), .op(
        n3638) );
  mux2_1 U15349 ( .ip1(n15781), .ip2(\ANSWER/mem[6][5][2] ), .s(n16782), .op(
        n3637) );
  mux2_1 U15350 ( .ip1(n15781), .ip2(\ANSWER/mem[6][6][2] ), .s(n16783), .op(
        n3636) );
  mux2_1 U15351 ( .ip1(n15781), .ip2(\ANSWER/mem[6][7][2] ), .s(n16784), .op(
        n3635) );
  mux2_1 U15352 ( .ip1(n15781), .ip2(\ANSWER/mem[6][8][2] ), .s(n16785), .op(
        n3634) );
  mux2_1 U15353 ( .ip1(n15781), .ip2(\ANSWER/mem[6][9][2] ), .s(n16786), .op(
        n3633) );
  mux2_1 U15354 ( .ip1(n15781), .ip2(\ANSWER/mem[7][0][2] ), .s(n16787), .op(
        n3632) );
  mux2_1 U15355 ( .ip1(n15781), .ip2(\ANSWER/mem[7][1][2] ), .s(n16788), .op(
        n3631) );
  buf_1 U15356 ( .ip(n15781), .op(n15782) );
  mux2_1 U15357 ( .ip1(n15782), .ip2(\ANSWER/mem[7][2][2] ), .s(n16790), .op(
        n3630) );
  mux2_1 U15358 ( .ip1(n15782), .ip2(\ANSWER/mem[7][3][2] ), .s(n16791), .op(
        n3629) );
  mux2_1 U15359 ( .ip1(n15781), .ip2(\ANSWER/mem[7][4][2] ), .s(n16792), .op(
        n3628) );
  mux2_1 U15360 ( .ip1(n15781), .ip2(\ANSWER/mem[7][5][2] ), .s(n16793), .op(
        n3627) );
  mux2_1 U15361 ( .ip1(n15782), .ip2(\ANSWER/mem[7][6][2] ), .s(n16794), .op(
        n3626) );
  mux2_1 U15362 ( .ip1(n15782), .ip2(\ANSWER/mem[7][7][2] ), .s(n16795), .op(
        n3625) );
  mux2_1 U15363 ( .ip1(n15782), .ip2(\ANSWER/mem[7][8][2] ), .s(n16796), .op(
        n3624) );
  mux2_1 U15364 ( .ip1(n15782), .ip2(\ANSWER/mem[7][9][2] ), .s(n16797), .op(
        n3623) );
  mux2_1 U15365 ( .ip1(n15782), .ip2(\ANSWER/mem[8][0][2] ), .s(n16798), .op(
        n3622) );
  mux2_1 U15366 ( .ip1(n15782), .ip2(\ANSWER/mem[8][1][2] ), .s(n16799), .op(
        n3621) );
  mux2_1 U15367 ( .ip1(n15782), .ip2(\ANSWER/mem[8][2][2] ), .s(n16800), .op(
        n3620) );
  mux2_1 U15368 ( .ip1(n15782), .ip2(\ANSWER/mem[8][3][2] ), .s(n16801), .op(
        n3619) );
  mux2_1 U15369 ( .ip1(n15781), .ip2(\ANSWER/mem[8][4][2] ), .s(n16803), .op(
        n3618) );
  mux2_1 U15370 ( .ip1(n15781), .ip2(\ANSWER/mem[8][5][2] ), .s(n16804), .op(
        n3617) );
  mux2_1 U15371 ( .ip1(n15781), .ip2(\ANSWER/mem[8][6][2] ), .s(n16805), .op(
        n3616) );
  mux2_1 U15372 ( .ip1(n15781), .ip2(\ANSWER/mem[8][7][2] ), .s(n16806), .op(
        n3615) );
  mux2_1 U15373 ( .ip1(n15781), .ip2(\ANSWER/mem[8][8][2] ), .s(n16807), .op(
        n3614) );
  mux2_1 U15374 ( .ip1(n15781), .ip2(\ANSWER/mem[8][9][2] ), .s(n16808), .op(
        n3613) );
  mux2_1 U15375 ( .ip1(n15781), .ip2(\ANSWER/mem[9][0][2] ), .s(n16809), .op(
        n3612) );
  mux2_1 U15376 ( .ip1(n15781), .ip2(\ANSWER/mem[9][1][2] ), .s(n16810), .op(
        n3611) );
  mux2_1 U15377 ( .ip1(n15781), .ip2(\ANSWER/mem[9][2][2] ), .s(n16811), .op(
        n3610) );
  mux2_1 U15378 ( .ip1(n15781), .ip2(\ANSWER/mem[9][3][2] ), .s(n16812), .op(
        n3609) );
  mux2_1 U15379 ( .ip1(n15781), .ip2(\ANSWER/mem[9][4][2] ), .s(n16813), .op(
        n3608) );
  mux2_1 U15380 ( .ip1(n15781), .ip2(\ANSWER/mem[9][5][2] ), .s(n16814), .op(
        n3607) );
  mux2_1 U15381 ( .ip1(n15782), .ip2(\ANSWER/mem[9][6][2] ), .s(n16815), .op(
        n3606) );
  mux2_1 U15382 ( .ip1(n15782), .ip2(\ANSWER/mem[9][7][2] ), .s(n16816), .op(
        n3605) );
  mux2_1 U15383 ( .ip1(n15782), .ip2(\ANSWER/mem[9][8][2] ), .s(n16817), .op(
        n3604) );
  mux2_1 U15384 ( .ip1(n15782), .ip2(\ANSWER/mem[9][9][2] ), .s(n16818), .op(
        n3603) );
  fulladder U15385 ( .a(n15785), .b(n15784), .ci(n15783), .co(n15856), .s(
        n15773) );
  nor2_1 U15386 ( .ip1(n15787), .ip2(n15786), .op(n15788) );
  nor2_1 U15387 ( .ip1(n15789), .ip2(n15788), .op(n15843) );
  inv_1 U15388 ( .ip(q_w2[11]), .op(n16599) );
  nor2_1 U15389 ( .ip1(n16369), .ip2(n16599), .op(n16055) );
  nand3_1 U15390 ( .ip1(m2DataIn[0]), .ip2(q_w2[8]), .ip3(n16055), .op(n15905)
         );
  nand2_1 U15391 ( .ip1(m2DataIn[0]), .ip2(q_w2[11]), .op(n15791) );
  nand2_1 U15392 ( .ip1(n15791), .ip2(n15790), .op(n15792) );
  nand2_1 U15393 ( .ip1(n15905), .ip2(n15792), .op(n15793) );
  inv_1 U15394 ( .ip(m2DataIn[11]), .op(n16679) );
  nor3_1 U15395 ( .ip1(n16679), .ip2(n15973), .ip3(n15793), .op(n15906) );
  or2_1 U15396 ( .ip1(n15793), .ip2(n15906), .op(n15796) );
  nand2_1 U15397 ( .ip1(m2DataIn[11]), .ip2(q_w2[0]), .op(n15794) );
  or2_1 U15398 ( .ip1(n15794), .ip2(n15906), .op(n15795) );
  nand2_1 U15399 ( .ip1(n15796), .ip2(n15795), .op(n15912) );
  nand2_1 U15400 ( .ip1(m2DataIn[4]), .ip2(q_w2[7]), .op(n15797) );
  nand4_1 U15401 ( .ip1(m2DataIn[5]), .ip2(m2DataIn[4]), .ip3(q_w2[6]), .ip4(
        q_w2[7]), .op(n15877) );
  inv_1 U15402 ( .ip(n15877), .op(n15798) );
  or2_1 U15403 ( .ip1(n15797), .ip2(n15798), .op(n15801) );
  or2_1 U15404 ( .ip1(n15799), .ip2(n15798), .op(n15800) );
  nand2_1 U15405 ( .ip1(n15801), .ip2(n15800), .op(n15875) );
  nor2_1 U15406 ( .ip1(n16600), .ip2(n16144), .op(n15802) );
  xor2_1 U15407 ( .ip1(n15875), .ip2(n15802), .op(n15911) );
  nand2_1 U15408 ( .ip1(m2DataIn[7]), .ip2(q_w2[5]), .op(n15867) );
  nor3_1 U15409 ( .ip1(n16273), .ip2(n16447), .ip3(n15867), .op(n15909) );
  inv_1 U15410 ( .ip(n15909), .op(n15806) );
  nand2_1 U15411 ( .ip1(m2DataIn[6]), .ip2(q_w2[5]), .op(n15804) );
  nand2_1 U15412 ( .ip1(n15804), .ip2(n15803), .op(n15805) );
  nand2_1 U15413 ( .ip1(n15806), .ip2(n15805), .op(n15807) );
  nor3_1 U15414 ( .ip1(n16690), .ip2(n16308), .ip3(n15807), .op(n15908) );
  or2_1 U15415 ( .ip1(n15807), .ip2(n15908), .op(n15810) );
  nand2_1 U15416 ( .ip1(m2DataIn[9]), .ip2(q_w2[2]), .op(n15808) );
  or2_1 U15417 ( .ip1(n15808), .ip2(n15908), .op(n15809) );
  nand2_1 U15418 ( .ip1(n15810), .ip2(n15809), .op(n15910) );
  inv_1 U15419 ( .ip(n15811), .op(n15919) );
  nor2_1 U15420 ( .ip1(n15813), .ip2(n15812), .op(n15916) );
  inv_1 U15421 ( .ip(rdata[3]), .op(n15818) );
  nand4_1 U15422 ( .ip1(m2DataIn[2]), .ip2(m2DataIn[1]), .ip3(q_w2[9]), .ip4(
        q_w2[10]), .op(n15890) );
  inv_1 U15423 ( .ip(n15890), .op(n15815) );
  or2_1 U15424 ( .ip1(n15814), .ip2(n15815), .op(n15817) );
  nand2_1 U15425 ( .ip1(m2DataIn[1]), .ip2(q_w2[10]), .op(n15900) );
  or2_1 U15426 ( .ip1(n15900), .ip2(n15815), .op(n15816) );
  nand2_1 U15427 ( .ip1(n15817), .ip2(n15816), .op(n15888) );
  mux2_1 U15428 ( .ip1(n15818), .ip2(rdata[3]), .s(n15888), .op(n15915) );
  nor2_1 U15429 ( .ip1(n15820), .ip2(n15819), .op(n15914) );
  fulladder U15430 ( .a(n15823), .b(n15822), .ci(n15821), .co(n15917), .s(
        n15769) );
  nand2_1 U15431 ( .ip1(m2DataIn[8]), .ip2(q_w2[3]), .op(n15896) );
  nor2_1 U15432 ( .ip1(n15825), .ip2(n15824), .op(n15826) );
  nor2_1 U15433 ( .ip1(n15827), .ip2(n15826), .op(n15895) );
  inv_1 U15434 ( .ip(n15828), .op(n15831) );
  nor3_1 U15435 ( .ip1(n16600), .ip2(n15973), .ip3(n15829), .op(n15830) );
  nor2_1 U15436 ( .ip1(n15831), .ip2(n15830), .op(n15894) );
  fulladder U15437 ( .a(n15834), .b(n15833), .ci(n15832), .co(n15835), .s(
        n15744) );
  inv_1 U15438 ( .ip(n15835), .op(n15898) );
  fulladder U15439 ( .a(n15838), .b(n15837), .ci(n15836), .co(n15897), .s(
        n15840) );
  fulladder U15440 ( .a(n15841), .b(n15840), .ci(n15839), .co(n15852), .s(
        n15759) );
  nor2_1 U15441 ( .ip1(n15843), .ip2(n15842), .op(n15855) );
  nand2_1 U15442 ( .ip1(n15843), .ip2(n15842), .op(n15857) );
  inv_1 U15443 ( .ip(n15857), .op(n15844) );
  nor2_1 U15444 ( .ip1(n15855), .ip2(n15844), .op(n15845) );
  xor2_1 U15445 ( .ip1(n15856), .ip2(n15845), .op(n15848) );
  nor3_1 U15446 ( .ip1(\SIGMOID/lut_out [2]), .ip2(\SIGMOID/lut_out [1]), 
        .ip3(\SIGMOID/N64 ), .op(n15846) );
  nor2_1 U15447 ( .ip1(\SIGMOID/sign_bit ), .ip2(n15846), .op(n15847) );
  xor2_1 U15448 ( .ip1(\SIGMOID/lut_out [3]), .ip2(n15847), .op(n17104) );
  mux2_1 U15449 ( .ip1(n15848), .ip2(n17104), .s(n16714), .op(n15849) );
  buf_1 U15450 ( .ip(n15849), .op(n15851) );
  mux2_1 U15451 ( .ip1(n15851), .ip2(\ANSWER/mem[0][0][3] ), .s(n16717), .op(
        n3602) );
  mux2_1 U15452 ( .ip1(n15851), .ip2(\ANSWER/mem[0][1][3] ), .s(n16718), .op(
        n3601) );
  mux2_1 U15453 ( .ip1(n15851), .ip2(\ANSWER/mem[0][2][3] ), .s(n16719), .op(
        n3600) );
  mux2_1 U15454 ( .ip1(n15851), .ip2(\ANSWER/mem[0][3][3] ), .s(n16720), .op(
        n3599) );
  mux2_1 U15455 ( .ip1(n15851), .ip2(\ANSWER/mem[0][4][3] ), .s(n16721), .op(
        n3598) );
  mux2_1 U15456 ( .ip1(n15851), .ip2(\ANSWER/mem[0][5][3] ), .s(n16722), .op(
        n3597) );
  mux2_1 U15457 ( .ip1(n15851), .ip2(\ANSWER/mem[0][6][3] ), .s(n16723), .op(
        n3596) );
  mux2_1 U15458 ( .ip1(n15851), .ip2(\ANSWER/mem[0][7][3] ), .s(n16724), .op(
        n3595) );
  mux2_1 U15459 ( .ip1(n15851), .ip2(\ANSWER/mem[0][8][3] ), .s(n16725), .op(
        n3594) );
  mux2_1 U15460 ( .ip1(n15851), .ip2(\ANSWER/mem[0][9][3] ), .s(n16726), .op(
        n3593) );
  mux2_1 U15461 ( .ip1(n15851), .ip2(\ANSWER/mem[1][0][3] ), .s(n16727), .op(
        n3592) );
  mux2_1 U15462 ( .ip1(n15851), .ip2(\ANSWER/mem[1][1][3] ), .s(n16728), .op(
        n3591) );
  mux2_1 U15463 ( .ip1(n15851), .ip2(\ANSWER/mem[1][2][3] ), .s(n16729), .op(
        n3590) );
  mux2_1 U15464 ( .ip1(n15849), .ip2(\ANSWER/mem[1][3][3] ), .s(n16730), .op(
        n3589) );
  mux2_1 U15465 ( .ip1(n15849), .ip2(\ANSWER/mem[1][4][3] ), .s(n16731), .op(
        n3588) );
  mux2_1 U15466 ( .ip1(n15849), .ip2(\ANSWER/mem[1][5][3] ), .s(n16732), .op(
        n3587) );
  mux2_1 U15467 ( .ip1(n15849), .ip2(\ANSWER/mem[1][6][3] ), .s(n16733), .op(
        n3586) );
  mux2_1 U15468 ( .ip1(n15849), .ip2(\ANSWER/mem[1][7][3] ), .s(n16734), .op(
        n3585) );
  mux2_1 U15469 ( .ip1(n15849), .ip2(\ANSWER/mem[1][8][3] ), .s(n16735), .op(
        n3584) );
  mux2_1 U15470 ( .ip1(n15849), .ip2(\ANSWER/mem[1][9][3] ), .s(n16736), .op(
        n3583) );
  mux2_1 U15471 ( .ip1(n15849), .ip2(\ANSWER/mem[2][0][3] ), .s(n16737), .op(
        n3582) );
  mux2_1 U15472 ( .ip1(n15849), .ip2(\ANSWER/mem[2][1][3] ), .s(n16738), .op(
        n3581) );
  mux2_1 U15473 ( .ip1(n15849), .ip2(\ANSWER/mem[2][2][3] ), .s(n16739), .op(
        n3580) );
  mux2_1 U15474 ( .ip1(n15849), .ip2(\ANSWER/mem[2][3][3] ), .s(n16740), .op(
        n3579) );
  mux2_1 U15475 ( .ip1(n15851), .ip2(\ANSWER/mem[2][4][3] ), .s(n16741), .op(
        n3578) );
  mux2_1 U15476 ( .ip1(n15849), .ip2(\ANSWER/mem[2][5][3] ), .s(n16742), .op(
        n3577) );
  mux2_1 U15477 ( .ip1(n15851), .ip2(\ANSWER/mem[2][6][3] ), .s(n16743), .op(
        n3576) );
  mux2_1 U15478 ( .ip1(n15849), .ip2(\ANSWER/mem[2][7][3] ), .s(n16744), .op(
        n3575) );
  mux2_1 U15479 ( .ip1(n15849), .ip2(\ANSWER/mem[2][8][3] ), .s(n16745), .op(
        n3574) );
  mux2_1 U15480 ( .ip1(n15849), .ip2(\ANSWER/mem[2][9][3] ), .s(n16746), .op(
        n3573) );
  mux2_1 U15481 ( .ip1(n15851), .ip2(\ANSWER/mem[3][0][3] ), .s(n16747), .op(
        n3572) );
  mux2_1 U15482 ( .ip1(n15851), .ip2(\ANSWER/mem[3][1][3] ), .s(n16748), .op(
        n3571) );
  mux2_1 U15483 ( .ip1(n15851), .ip2(\ANSWER/mem[3][2][3] ), .s(n16749), .op(
        n3570) );
  mux2_1 U15484 ( .ip1(n15851), .ip2(\ANSWER/mem[3][3][3] ), .s(n16750), .op(
        n3569) );
  mux2_1 U15485 ( .ip1(n15851), .ip2(\ANSWER/mem[3][4][3] ), .s(n16751), .op(
        n3568) );
  mux2_1 U15486 ( .ip1(n15851), .ip2(\ANSWER/mem[3][5][3] ), .s(n16752), .op(
        n3567) );
  buf_1 U15487 ( .ip(n15849), .op(n15850) );
  mux2_1 U15488 ( .ip1(n15850), .ip2(\ANSWER/mem[3][6][3] ), .s(n16753), .op(
        n3566) );
  mux2_1 U15489 ( .ip1(n15849), .ip2(\ANSWER/mem[3][7][3] ), .s(n16754), .op(
        n3565) );
  mux2_1 U15490 ( .ip1(n15849), .ip2(\ANSWER/mem[3][8][3] ), .s(n16755), .op(
        n3564) );
  mux2_1 U15491 ( .ip1(n15849), .ip2(\ANSWER/mem[3][9][3] ), .s(n16756), .op(
        n3563) );
  mux2_1 U15492 ( .ip1(n15850), .ip2(\ANSWER/mem[4][0][3] ), .s(n16757), .op(
        n3562) );
  mux2_1 U15493 ( .ip1(n15850), .ip2(\ANSWER/mem[4][1][3] ), .s(n16758), .op(
        n3561) );
  mux2_1 U15494 ( .ip1(n15850), .ip2(\ANSWER/mem[4][2][3] ), .s(n16759), .op(
        n3560) );
  mux2_1 U15495 ( .ip1(n15850), .ip2(\ANSWER/mem[4][3][3] ), .s(n16760), .op(
        n3559) );
  mux2_1 U15496 ( .ip1(n15850), .ip2(\ANSWER/mem[4][4][3] ), .s(n16761), .op(
        n3558) );
  mux2_1 U15497 ( .ip1(n15850), .ip2(\ANSWER/mem[4][5][3] ), .s(n16762), .op(
        n3557) );
  mux2_1 U15498 ( .ip1(n15850), .ip2(\ANSWER/mem[4][6][3] ), .s(n16763), .op(
        n3556) );
  mux2_1 U15499 ( .ip1(n15850), .ip2(\ANSWER/mem[4][7][3] ), .s(n16764), .op(
        n3555) );
  mux2_1 U15500 ( .ip1(n15851), .ip2(\ANSWER/mem[4][8][3] ), .s(n16765), .op(
        n3554) );
  mux2_1 U15501 ( .ip1(n15849), .ip2(\ANSWER/mem[4][9][3] ), .s(n16766), .op(
        n3553) );
  mux2_1 U15502 ( .ip1(n15849), .ip2(\ANSWER/mem[5][0][3] ), .s(n16767), .op(
        n3552) );
  mux2_1 U15503 ( .ip1(n15849), .ip2(\ANSWER/mem[5][1][3] ), .s(n16768), .op(
        n3551) );
  mux2_1 U15504 ( .ip1(n15849), .ip2(\ANSWER/mem[5][2][3] ), .s(n16769), .op(
        n3550) );
  mux2_1 U15505 ( .ip1(n15849), .ip2(\ANSWER/mem[5][3][3] ), .s(n16770), .op(
        n3549) );
  mux2_1 U15506 ( .ip1(n15849), .ip2(\ANSWER/mem[5][4][3] ), .s(n16771), .op(
        n3548) );
  mux2_1 U15507 ( .ip1(n15849), .ip2(\ANSWER/mem[5][5][3] ), .s(n16772), .op(
        n3547) );
  mux2_1 U15508 ( .ip1(n15849), .ip2(\ANSWER/mem[5][6][3] ), .s(n16773), .op(
        n3546) );
  mux2_1 U15509 ( .ip1(n15849), .ip2(\ANSWER/mem[5][7][3] ), .s(n16774), .op(
        n3545) );
  mux2_1 U15510 ( .ip1(n15849), .ip2(\ANSWER/mem[5][8][3] ), .s(n16775), .op(
        n3544) );
  mux2_1 U15511 ( .ip1(n15849), .ip2(\ANSWER/mem[5][9][3] ), .s(n16776), .op(
        n3543) );
  mux2_1 U15512 ( .ip1(n15850), .ip2(\ANSWER/mem[6][0][3] ), .s(n16777), .op(
        n3542) );
  mux2_1 U15513 ( .ip1(n15850), .ip2(\ANSWER/mem[6][1][3] ), .s(n16778), .op(
        n3541) );
  mux2_1 U15514 ( .ip1(n15850), .ip2(\ANSWER/mem[6][2][3] ), .s(n16779), .op(
        n3540) );
  mux2_1 U15515 ( .ip1(n15850), .ip2(\ANSWER/mem[6][3][3] ), .s(n16780), .op(
        n3539) );
  mux2_1 U15516 ( .ip1(n15849), .ip2(\ANSWER/mem[6][4][3] ), .s(n16781), .op(
        n3538) );
  mux2_1 U15517 ( .ip1(n15849), .ip2(\ANSWER/mem[6][5][3] ), .s(n16782), .op(
        n3537) );
  mux2_1 U15518 ( .ip1(n15849), .ip2(\ANSWER/mem[6][6][3] ), .s(n16783), .op(
        n3536) );
  mux2_1 U15519 ( .ip1(n15849), .ip2(\ANSWER/mem[6][7][3] ), .s(n16784), .op(
        n3535) );
  mux2_1 U15520 ( .ip1(n15849), .ip2(\ANSWER/mem[6][8][3] ), .s(n16785), .op(
        n3534) );
  mux2_1 U15521 ( .ip1(n15849), .ip2(\ANSWER/mem[6][9][3] ), .s(n16786), .op(
        n3533) );
  mux2_1 U15522 ( .ip1(n15849), .ip2(\ANSWER/mem[7][0][3] ), .s(n16787), .op(
        n3532) );
  mux2_1 U15523 ( .ip1(n15849), .ip2(\ANSWER/mem[7][1][3] ), .s(n16788), .op(
        n3531) );
  mux2_1 U15524 ( .ip1(n15850), .ip2(\ANSWER/mem[7][2][3] ), .s(n16790), .op(
        n3530) );
  mux2_1 U15525 ( .ip1(n15850), .ip2(\ANSWER/mem[7][3][3] ), .s(n16791), .op(
        n3529) );
  mux2_1 U15526 ( .ip1(n15850), .ip2(\ANSWER/mem[7][4][3] ), .s(n16792), .op(
        n3528) );
  mux2_1 U15527 ( .ip1(n15850), .ip2(\ANSWER/mem[7][5][3] ), .s(n16793), .op(
        n3527) );
  mux2_1 U15528 ( .ip1(n15850), .ip2(\ANSWER/mem[7][6][3] ), .s(n16794), .op(
        n3526) );
  mux2_1 U15529 ( .ip1(n15850), .ip2(\ANSWER/mem[7][7][3] ), .s(n16795), .op(
        n3525) );
  mux2_1 U15530 ( .ip1(n15850), .ip2(\ANSWER/mem[7][8][3] ), .s(n16796), .op(
        n3524) );
  mux2_1 U15531 ( .ip1(n15850), .ip2(\ANSWER/mem[7][9][3] ), .s(n16797), .op(
        n3523) );
  mux2_1 U15532 ( .ip1(n15850), .ip2(\ANSWER/mem[8][0][3] ), .s(n16798), .op(
        n3522) );
  mux2_1 U15533 ( .ip1(n15850), .ip2(\ANSWER/mem[8][1][3] ), .s(n16799), .op(
        n3521) );
  mux2_1 U15534 ( .ip1(n15850), .ip2(\ANSWER/mem[8][2][3] ), .s(n16800), .op(
        n3520) );
  mux2_1 U15535 ( .ip1(n15850), .ip2(\ANSWER/mem[8][3][3] ), .s(n16801), .op(
        n3519) );
  mux2_1 U15536 ( .ip1(n15850), .ip2(\ANSWER/mem[8][4][3] ), .s(n16803), .op(
        n3518) );
  mux2_1 U15537 ( .ip1(n15849), .ip2(\ANSWER/mem[8][5][3] ), .s(n16804), .op(
        n3517) );
  mux2_1 U15538 ( .ip1(n15851), .ip2(\ANSWER/mem[8][6][3] ), .s(n16805), .op(
        n3516) );
  mux2_1 U15539 ( .ip1(n15850), .ip2(\ANSWER/mem[8][7][3] ), .s(n16806), .op(
        n3515) );
  mux2_1 U15540 ( .ip1(n15851), .ip2(\ANSWER/mem[8][8][3] ), .s(n16807), .op(
        n3514) );
  mux2_1 U15541 ( .ip1(n15850), .ip2(\ANSWER/mem[8][9][3] ), .s(n16808), .op(
        n3513) );
  mux2_1 U15542 ( .ip1(n15851), .ip2(\ANSWER/mem[9][0][3] ), .s(n16809), .op(
        n3512) );
  mux2_1 U15543 ( .ip1(n15850), .ip2(\ANSWER/mem[9][1][3] ), .s(n16810), .op(
        n3511) );
  mux2_1 U15544 ( .ip1(n15851), .ip2(\ANSWER/mem[9][2][3] ), .s(n16811), .op(
        n3510) );
  mux2_1 U15545 ( .ip1(n15850), .ip2(\ANSWER/mem[9][3][3] ), .s(n16812), .op(
        n3509) );
  mux2_1 U15546 ( .ip1(n15851), .ip2(\ANSWER/mem[9][4][3] ), .s(n16813), .op(
        n3508) );
  mux2_1 U15547 ( .ip1(n15850), .ip2(\ANSWER/mem[9][5][3] ), .s(n16814), .op(
        n3507) );
  mux2_1 U15548 ( .ip1(n15851), .ip2(\ANSWER/mem[9][6][3] ), .s(n16815), .op(
        n3506) );
  mux2_1 U15549 ( .ip1(n15851), .ip2(\ANSWER/mem[9][7][3] ), .s(n16816), .op(
        n3505) );
  mux2_1 U15550 ( .ip1(n15851), .ip2(\ANSWER/mem[9][8][3] ), .s(n16817), .op(
        n3504) );
  mux2_1 U15551 ( .ip1(n15851), .ip2(\ANSWER/mem[9][9][3] ), .s(n16818), .op(
        n3503) );
  fulladder U15552 ( .a(n15854), .b(n15853), .ci(n15852), .co(n15924), .s(
        n15842) );
  inv_1 U15553 ( .ip(n15924), .op(n15996) );
  or2_1 U15554 ( .ip1(n15856), .ip2(n15855), .op(n15858) );
  nand2_1 U15555 ( .ip1(n15858), .ip2(n15857), .op(n15921) );
  nand2_1 U15556 ( .ip1(m2DataIn[5]), .ip2(q_w2[8]), .op(n15961) );
  nor3_1 U15557 ( .ip1(n16445), .ip2(n16561), .ip3(n15961), .op(n15960) );
  inv_1 U15558 ( .ip(n15960), .op(n15862) );
  nand2_1 U15559 ( .ip1(m2DataIn[4]), .ip2(q_w2[8]), .op(n15860) );
  nand2_1 U15560 ( .ip1(m2DataIn[5]), .ip2(q_w2[7]), .op(n15859) );
  nand2_1 U15561 ( .ip1(n15860), .ip2(n15859), .op(n15861) );
  nand2_1 U15562 ( .ip1(n15862), .ip2(n15861), .op(n15863) );
  nor3_1 U15563 ( .ip1(n16679), .ip2(n16144), .ip3(n15863), .op(n15959) );
  or2_1 U15564 ( .ip1(n15863), .ip2(n15959), .op(n15866) );
  nand2_1 U15565 ( .ip1(m2DataIn[11]), .ip2(q_w2[1]), .op(n15864) );
  or2_1 U15566 ( .ip1(n15864), .ip2(n15959), .op(n15865) );
  nand2_1 U15567 ( .ip1(n15866), .ip2(n15865), .op(n15945) );
  nand2_1 U15568 ( .ip1(m2DataIn[7]), .ip2(q_w2[6]), .op(n15975) );
  nor3_1 U15569 ( .ip1(n16273), .ip2(n16497), .ip3(n15975), .op(n15983) );
  inv_1 U15570 ( .ip(n15983), .op(n15870) );
  nand2_1 U15571 ( .ip1(m2DataIn[6]), .ip2(q_w2[6]), .op(n15868) );
  nand2_1 U15572 ( .ip1(n15868), .ip2(n15867), .op(n15869) );
  nand2_1 U15573 ( .ip1(n15870), .ip2(n15869), .op(n15871) );
  nor3_1 U15574 ( .ip1(n16600), .ip2(n16308), .ip3(n15871), .op(n15982) );
  or2_1 U15575 ( .ip1(n15871), .ip2(n15982), .op(n15874) );
  nand2_1 U15576 ( .ip1(m2DataIn[10]), .ip2(q_w2[2]), .op(n15872) );
  or2_1 U15577 ( .ip1(n15872), .ip2(n15982), .op(n15873) );
  nand2_1 U15578 ( .ip1(n15874), .ip2(n15873), .op(n15944) );
  nand3_1 U15579 ( .ip1(m2DataIn[10]), .ip2(q_w2[1]), .ip3(n15875), .op(n15876) );
  nand2_1 U15580 ( .ip1(n15877), .ip2(n15876), .op(n15943) );
  inv_1 U15581 ( .ip(n15878), .op(n15994) );
  inv_1 U15582 ( .ip(m2DataIn[12]), .op(n16623) );
  nor2_1 U15583 ( .ip1(n16623), .ip2(n15973), .op(n15883) );
  nand2_1 U15584 ( .ip1(m2DataIn[3]), .ip2(q_w2[12]), .op(n16197) );
  nor3_1 U15585 ( .ip1(n16145), .ip2(n16552), .ip3(n16197), .op(n15958) );
  or2_1 U15586 ( .ip1(q_w2[12]), .ip2(n15879), .op(n15881) );
  or2_1 U15587 ( .ip1(m2DataIn[0]), .ip2(n15879), .op(n15880) );
  nand2_1 U15588 ( .ip1(n15881), .ip2(n15880), .op(n15882) );
  or2_1 U15589 ( .ip1(n15958), .ip2(n15882), .op(n15956) );
  xor2_1 U15590 ( .ip1(n15883), .ip2(n15956), .op(n15936) );
  nand2_1 U15591 ( .ip1(m2DataIn[8]), .ip2(q_w2[4]), .op(n15952) );
  nand4_1 U15592 ( .ip1(m2DataIn[8]), .ip2(m2DataIn[9]), .ip3(q_w2[3]), .ip4(
        q_w2[4]), .op(n15942) );
  inv_1 U15593 ( .ip(n15942), .op(n15884) );
  or2_1 U15594 ( .ip1(n15952), .ip2(n15884), .op(n15887) );
  nand2_1 U15595 ( .ip1(m2DataIn[9]), .ip2(q_w2[3]), .op(n15885) );
  or2_1 U15596 ( .ip1(n15885), .ip2(n15884), .op(n15886) );
  nand2_1 U15597 ( .ip1(n15887), .ip2(n15886), .op(n15892) );
  nand2_1 U15598 ( .ip1(rdata[3]), .ip2(n15888), .op(n15889) );
  nand2_1 U15599 ( .ip1(n15890), .ip2(n15889), .op(n15891) );
  nand2_1 U15600 ( .ip1(n15892), .ip2(n15891), .op(n15941) );
  or2_1 U15601 ( .ip1(n15892), .ip2(n15891), .op(n15893) );
  nand2_1 U15602 ( .ip1(n15941), .ip2(n15893), .op(n15935) );
  fulladder U15603 ( .a(n15896), .b(n15895), .ci(n15894), .co(n15934), .s(
        n15899) );
  fulladder U15604 ( .a(n15899), .b(n15898), .ci(n15897), .co(n15992), .s(
        n15853) );
  nand2_1 U15605 ( .ip1(m2DataIn[2]), .ip2(q_w2[11]), .op(n15984) );
  nor2_1 U15606 ( .ip1(n15900), .ip2(n15984), .op(n15991) );
  inv_1 U15607 ( .ip(n15991), .op(n15904) );
  nand2_1 U15608 ( .ip1(m2DataIn[2]), .ip2(q_w2[10]), .op(n15902) );
  nand2_1 U15609 ( .ip1(m2DataIn[1]), .ip2(q_w2[11]), .op(n15901) );
  nand2_1 U15610 ( .ip1(n15902), .ip2(n15901), .op(n15903) );
  nand2_1 U15611 ( .ip1(n15904), .ip2(n15903), .op(n15988) );
  mux2_1 U15612 ( .ip1(rdata[4]), .ip2(n15989), .s(n15988), .op(n15939) );
  inv_1 U15613 ( .ip(n15905), .op(n15907) );
  nor2_1 U15614 ( .ip1(n15907), .ip2(n15906), .op(n15938) );
  nor2_1 U15615 ( .ip1(n15909), .ip2(n15908), .op(n15937) );
  fulladder U15616 ( .a(n15912), .b(n15911), .ci(n15910), .co(n15913), .s(
        n15811) );
  inv_1 U15617 ( .ip(n15913), .op(n15948) );
  fulladder U15618 ( .a(n15916), .b(n15915), .ci(n15914), .co(n15947), .s(
        n15918) );
  fulladder U15619 ( .a(n15919), .b(n15918), .ci(n15917), .co(n15931), .s(
        n15854) );
  nor2_1 U15620 ( .ip1(n15921), .ip2(n15920), .op(n15995) );
  nand2_1 U15621 ( .ip1(n15921), .ip2(n15920), .op(n15998) );
  inv_1 U15622 ( .ip(n15998), .op(n15922) );
  nor2_1 U15623 ( .ip1(n15995), .ip2(n15922), .op(n15923) );
  mux2_1 U15624 ( .ip1(n15996), .ip2(n15924), .s(n15923), .op(n15927) );
  inv_1 U15625 ( .ip(\SIGMOID/lut_out [4]), .op(n15926) );
  or4_1 U15626 ( .ip1(\SIGMOID/lut_out [3]), .ip2(\SIGMOID/lut_out [2]), .ip3(
        \SIGMOID/lut_out [1]), .ip4(\SIGMOID/N64 ), .op(n16002) );
  nand2_1 U15627 ( .ip1(n16164), .ip2(n16002), .op(n15925) );
  mux2_1 U15628 ( .ip1(n15926), .ip2(\SIGMOID/lut_out [4]), .s(n15925), .op(
        n17137) );
  mux2_1 U15629 ( .ip1(n15927), .ip2(n17137), .s(n16714), .op(n15928) );
  mux2_1 U15630 ( .ip1(n15928), .ip2(\ANSWER/mem[0][0][4] ), .s(n16717), .op(
        n3502) );
  buf_1 U15631 ( .ip(n15928), .op(n15930) );
  mux2_1 U15632 ( .ip1(n15930), .ip2(\ANSWER/mem[0][1][4] ), .s(n16718), .op(
        n3501) );
  mux2_1 U15633 ( .ip1(n15930), .ip2(\ANSWER/mem[0][2][4] ), .s(n16719), .op(
        n3500) );
  buf_1 U15634 ( .ip(n15928), .op(n15929) );
  mux2_1 U15635 ( .ip1(n15929), .ip2(\ANSWER/mem[0][3][4] ), .s(n16720), .op(
        n3499) );
  mux2_1 U15636 ( .ip1(n15930), .ip2(\ANSWER/mem[0][4][4] ), .s(n16721), .op(
        n3498) );
  mux2_1 U15637 ( .ip1(n15929), .ip2(\ANSWER/mem[0][5][4] ), .s(n16722), .op(
        n3497) );
  mux2_1 U15638 ( .ip1(n15930), .ip2(\ANSWER/mem[0][6][4] ), .s(n16723), .op(
        n3496) );
  mux2_1 U15639 ( .ip1(n15929), .ip2(\ANSWER/mem[0][7][4] ), .s(n16724), .op(
        n3495) );
  mux2_1 U15640 ( .ip1(n15930), .ip2(\ANSWER/mem[0][8][4] ), .s(n16725), .op(
        n3494) );
  mux2_1 U15641 ( .ip1(n15929), .ip2(\ANSWER/mem[0][9][4] ), .s(n16726), .op(
        n3493) );
  mux2_1 U15642 ( .ip1(n15930), .ip2(\ANSWER/mem[1][0][4] ), .s(n16727), .op(
        n3492) );
  mux2_1 U15643 ( .ip1(n15929), .ip2(\ANSWER/mem[1][1][4] ), .s(n16728), .op(
        n3491) );
  mux2_1 U15644 ( .ip1(n15928), .ip2(\ANSWER/mem[1][2][4] ), .s(n16729), .op(
        n3490) );
  mux2_1 U15645 ( .ip1(n15928), .ip2(\ANSWER/mem[1][3][4] ), .s(n16730), .op(
        n3489) );
  mux2_1 U15646 ( .ip1(n15928), .ip2(\ANSWER/mem[1][4][4] ), .s(n16731), .op(
        n3488) );
  mux2_1 U15647 ( .ip1(n15928), .ip2(\ANSWER/mem[1][5][4] ), .s(n16732), .op(
        n3487) );
  mux2_1 U15648 ( .ip1(n15930), .ip2(\ANSWER/mem[1][6][4] ), .s(n16733), .op(
        n3486) );
  mux2_1 U15649 ( .ip1(n15930), .ip2(\ANSWER/mem[1][7][4] ), .s(n16734), .op(
        n3485) );
  mux2_1 U15650 ( .ip1(n15929), .ip2(\ANSWER/mem[1][8][4] ), .s(n16735), .op(
        n3484) );
  mux2_1 U15651 ( .ip1(n15929), .ip2(\ANSWER/mem[1][9][4] ), .s(n16736), .op(
        n3483) );
  mux2_1 U15652 ( .ip1(n15928), .ip2(\ANSWER/mem[2][0][4] ), .s(n16737), .op(
        n3482) );
  mux2_1 U15653 ( .ip1(n15928), .ip2(\ANSWER/mem[2][1][4] ), .s(n16738), .op(
        n3481) );
  mux2_1 U15654 ( .ip1(n15928), .ip2(\ANSWER/mem[2][2][4] ), .s(n16739), .op(
        n3480) );
  mux2_1 U15655 ( .ip1(n15928), .ip2(\ANSWER/mem[2][3][4] ), .s(n16740), .op(
        n3479) );
  mux2_1 U15656 ( .ip1(n15928), .ip2(\ANSWER/mem[2][4][4] ), .s(n16741), .op(
        n3478) );
  mux2_1 U15657 ( .ip1(n15928), .ip2(\ANSWER/mem[2][5][4] ), .s(n16742), .op(
        n3477) );
  mux2_1 U15658 ( .ip1(n15928), .ip2(\ANSWER/mem[2][6][4] ), .s(n16743), .op(
        n3476) );
  mux2_1 U15659 ( .ip1(n15928), .ip2(\ANSWER/mem[2][7][4] ), .s(n16744), .op(
        n3475) );
  mux2_1 U15660 ( .ip1(n15928), .ip2(\ANSWER/mem[2][8][4] ), .s(n16745), .op(
        n3474) );
  mux2_1 U15661 ( .ip1(n15928), .ip2(\ANSWER/mem[2][9][4] ), .s(n16746), .op(
        n3473) );
  mux2_1 U15662 ( .ip1(n15928), .ip2(\ANSWER/mem[3][0][4] ), .s(n16747), .op(
        n3472) );
  mux2_1 U15663 ( .ip1(n15928), .ip2(\ANSWER/mem[3][1][4] ), .s(n16748), .op(
        n3471) );
  mux2_1 U15664 ( .ip1(n15928), .ip2(\ANSWER/mem[3][2][4] ), .s(n16749), .op(
        n3470) );
  mux2_1 U15665 ( .ip1(n15928), .ip2(\ANSWER/mem[3][3][4] ), .s(n16750), .op(
        n3469) );
  mux2_1 U15666 ( .ip1(n15928), .ip2(\ANSWER/mem[3][4][4] ), .s(n16751), .op(
        n3468) );
  mux2_1 U15667 ( .ip1(n15928), .ip2(\ANSWER/mem[3][5][4] ), .s(n16752), .op(
        n3467) );
  mux2_1 U15668 ( .ip1(n15928), .ip2(\ANSWER/mem[3][6][4] ), .s(n16753), .op(
        n3466) );
  mux2_1 U15669 ( .ip1(n15928), .ip2(\ANSWER/mem[3][7][4] ), .s(n16754), .op(
        n3465) );
  mux2_1 U15670 ( .ip1(n15928), .ip2(\ANSWER/mem[3][8][4] ), .s(n16755), .op(
        n3464) );
  mux2_1 U15671 ( .ip1(n15928), .ip2(\ANSWER/mem[3][9][4] ), .s(n16756), .op(
        n3463) );
  mux2_1 U15672 ( .ip1(n15929), .ip2(\ANSWER/mem[4][0][4] ), .s(n16757), .op(
        n3462) );
  mux2_1 U15673 ( .ip1(n15930), .ip2(\ANSWER/mem[4][1][4] ), .s(n16758), .op(
        n3461) );
  mux2_1 U15674 ( .ip1(n15930), .ip2(\ANSWER/mem[4][2][4] ), .s(n16759), .op(
        n3460) );
  mux2_1 U15675 ( .ip1(n15929), .ip2(\ANSWER/mem[4][3][4] ), .s(n16760), .op(
        n3459) );
  mux2_1 U15676 ( .ip1(n15929), .ip2(\ANSWER/mem[4][4][4] ), .s(n16761), .op(
        n3458) );
  mux2_1 U15677 ( .ip1(n15928), .ip2(\ANSWER/mem[4][5][4] ), .s(n16762), .op(
        n3457) );
  mux2_1 U15678 ( .ip1(n15928), .ip2(\ANSWER/mem[4][6][4] ), .s(n16763), .op(
        n3456) );
  mux2_1 U15679 ( .ip1(n15928), .ip2(\ANSWER/mem[4][7][4] ), .s(n16764), .op(
        n3455) );
  mux2_1 U15680 ( .ip1(n15930), .ip2(\ANSWER/mem[4][8][4] ), .s(n16765), .op(
        n3454) );
  mux2_1 U15681 ( .ip1(n15930), .ip2(\ANSWER/mem[4][9][4] ), .s(n16766), .op(
        n3453) );
  mux2_1 U15682 ( .ip1(n15930), .ip2(\ANSWER/mem[5][0][4] ), .s(n16767), .op(
        n3452) );
  mux2_1 U15683 ( .ip1(n15930), .ip2(\ANSWER/mem[5][1][4] ), .s(n16768), .op(
        n3451) );
  mux2_1 U15684 ( .ip1(n15929), .ip2(\ANSWER/mem[5][2][4] ), .s(n16769), .op(
        n3450) );
  mux2_1 U15685 ( .ip1(n15928), .ip2(\ANSWER/mem[5][3][4] ), .s(n16770), .op(
        n3449) );
  mux2_1 U15686 ( .ip1(n15930), .ip2(\ANSWER/mem[5][4][4] ), .s(n16771), .op(
        n3448) );
  mux2_1 U15687 ( .ip1(n15929), .ip2(\ANSWER/mem[5][5][4] ), .s(n16772), .op(
        n3447) );
  mux2_1 U15688 ( .ip1(n15928), .ip2(\ANSWER/mem[5][6][4] ), .s(n16773), .op(
        n3446) );
  mux2_1 U15689 ( .ip1(n15930), .ip2(\ANSWER/mem[5][7][4] ), .s(n16774), .op(
        n3445) );
  mux2_1 U15690 ( .ip1(n15929), .ip2(\ANSWER/mem[5][8][4] ), .s(n16775), .op(
        n3444) );
  mux2_1 U15691 ( .ip1(n15928), .ip2(\ANSWER/mem[5][9][4] ), .s(n16776), .op(
        n3443) );
  mux2_1 U15692 ( .ip1(n15930), .ip2(\ANSWER/mem[6][0][4] ), .s(n16777), .op(
        n3442) );
  mux2_1 U15693 ( .ip1(n15929), .ip2(\ANSWER/mem[6][1][4] ), .s(n16778), .op(
        n3441) );
  mux2_1 U15694 ( .ip1(n15930), .ip2(\ANSWER/mem[6][2][4] ), .s(n16779), .op(
        n3440) );
  mux2_1 U15695 ( .ip1(n15930), .ip2(\ANSWER/mem[6][3][4] ), .s(n16780), .op(
        n3439) );
  mux2_1 U15696 ( .ip1(n15930), .ip2(\ANSWER/mem[6][4][4] ), .s(n16781), .op(
        n3438) );
  mux2_1 U15697 ( .ip1(n15930), .ip2(\ANSWER/mem[6][5][4] ), .s(n16782), .op(
        n3437) );
  mux2_1 U15698 ( .ip1(n15930), .ip2(\ANSWER/mem[6][6][4] ), .s(n16783), .op(
        n3436) );
  mux2_1 U15699 ( .ip1(n15928), .ip2(\ANSWER/mem[6][7][4] ), .s(n16784), .op(
        n3435) );
  mux2_1 U15700 ( .ip1(n15929), .ip2(\ANSWER/mem[6][8][4] ), .s(n16785), .op(
        n3434) );
  mux2_1 U15701 ( .ip1(n15930), .ip2(\ANSWER/mem[6][9][4] ), .s(n16786), .op(
        n3433) );
  mux2_1 U15702 ( .ip1(n15928), .ip2(\ANSWER/mem[7][0][4] ), .s(n16787), .op(
        n3432) );
  mux2_1 U15703 ( .ip1(n15930), .ip2(\ANSWER/mem[7][1][4] ), .s(n16788), .op(
        n3431) );
  mux2_1 U15704 ( .ip1(n15928), .ip2(\ANSWER/mem[7][2][4] ), .s(n16790), .op(
        n3430) );
  mux2_1 U15705 ( .ip1(n15930), .ip2(\ANSWER/mem[7][3][4] ), .s(n16791), .op(
        n3429) );
  mux2_1 U15706 ( .ip1(n15928), .ip2(\ANSWER/mem[7][4][4] ), .s(n16792), .op(
        n3428) );
  mux2_1 U15707 ( .ip1(n15929), .ip2(\ANSWER/mem[7][5][4] ), .s(n16793), .op(
        n3427) );
  mux2_1 U15708 ( .ip1(n15929), .ip2(\ANSWER/mem[7][6][4] ), .s(n16794), .op(
        n3426) );
  mux2_1 U15709 ( .ip1(n15928), .ip2(\ANSWER/mem[7][7][4] ), .s(n16795), .op(
        n3425) );
  mux2_1 U15710 ( .ip1(n15928), .ip2(\ANSWER/mem[7][8][4] ), .s(n16796), .op(
        n3424) );
  mux2_1 U15711 ( .ip1(n15928), .ip2(\ANSWER/mem[7][9][4] ), .s(n16797), .op(
        n3423) );
  mux2_1 U15712 ( .ip1(n15929), .ip2(\ANSWER/mem[8][0][4] ), .s(n16798), .op(
        n3422) );
  mux2_1 U15713 ( .ip1(n15930), .ip2(\ANSWER/mem[8][1][4] ), .s(n16799), .op(
        n3421) );
  mux2_1 U15714 ( .ip1(n15929), .ip2(\ANSWER/mem[8][2][4] ), .s(n16800), .op(
        n3420) );
  mux2_1 U15715 ( .ip1(n15930), .ip2(\ANSWER/mem[8][3][4] ), .s(n16801), .op(
        n3419) );
  mux2_1 U15716 ( .ip1(n15929), .ip2(\ANSWER/mem[8][4][4] ), .s(n16803), .op(
        n3418) );
  mux2_1 U15717 ( .ip1(n15929), .ip2(\ANSWER/mem[8][5][4] ), .s(n16804), .op(
        n3417) );
  mux2_1 U15718 ( .ip1(n15929), .ip2(\ANSWER/mem[8][6][4] ), .s(n16805), .op(
        n3416) );
  mux2_1 U15719 ( .ip1(n15929), .ip2(\ANSWER/mem[8][7][4] ), .s(n16806), .op(
        n3415) );
  mux2_1 U15720 ( .ip1(n15929), .ip2(\ANSWER/mem[8][8][4] ), .s(n16807), .op(
        n3414) );
  mux2_1 U15721 ( .ip1(n15929), .ip2(\ANSWER/mem[8][9][4] ), .s(n16808), .op(
        n3413) );
  mux2_1 U15722 ( .ip1(n15929), .ip2(\ANSWER/mem[9][0][4] ), .s(n16809), .op(
        n3412) );
  mux2_1 U15723 ( .ip1(n15929), .ip2(\ANSWER/mem[9][1][4] ), .s(n16810), .op(
        n3411) );
  mux2_1 U15724 ( .ip1(n15929), .ip2(\ANSWER/mem[9][2][4] ), .s(n16811), .op(
        n3410) );
  mux2_1 U15725 ( .ip1(n15929), .ip2(\ANSWER/mem[9][3][4] ), .s(n16812), .op(
        n3409) );
  mux2_1 U15726 ( .ip1(n15929), .ip2(\ANSWER/mem[9][4][4] ), .s(n16813), .op(
        n3408) );
  mux2_1 U15727 ( .ip1(n15929), .ip2(\ANSWER/mem[9][5][4] ), .s(n16814), .op(
        n3407) );
  mux2_1 U15728 ( .ip1(n15930), .ip2(\ANSWER/mem[9][6][4] ), .s(n16815), .op(
        n3406) );
  mux2_1 U15729 ( .ip1(n15930), .ip2(\ANSWER/mem[9][7][4] ), .s(n16816), .op(
        n3405) );
  mux2_1 U15730 ( .ip1(n15930), .ip2(\ANSWER/mem[9][8][4] ), .s(n16817), .op(
        n3404) );
  mux2_1 U15731 ( .ip1(n15930), .ip2(\ANSWER/mem[9][9][4] ), .s(n16818), .op(
        n3403) );
  fulladder U15732 ( .a(n15933), .b(n15932), .ci(n15931), .co(n16071), .s(
        n15920) );
  fulladder U15733 ( .a(n15936), .b(n15935), .ci(n15934), .co(n16069), .s(
        n15993) );
  fulladder U15734 ( .a(n15939), .b(n15938), .ci(n15937), .co(n15940), .s(
        n15949) );
  inv_1 U15735 ( .ip(n15940), .op(n16039) );
  nand2_1 U15736 ( .ip1(n15942), .ip2(n15941), .op(n16038) );
  fulladder U15737 ( .a(n15945), .b(n15944), .ci(n15943), .co(n16037), .s(
        n15878) );
  inv_1 U15738 ( .ip(n15946), .op(n16068) );
  fulladder U15739 ( .a(n15949), .b(n15948), .ci(n15947), .co(n16067), .s(
        n15932) );
  nor2_1 U15740 ( .ip1(n16600), .ip2(n16177), .op(n15955) );
  nand2_1 U15741 ( .ip1(q_w2[5]), .ip2(m2DataIn[8]), .op(n15951) );
  nand2_1 U15742 ( .ip1(m2DataIn[9]), .ip2(q_w2[4]), .op(n15950) );
  nand2_1 U15743 ( .ip1(n15951), .ip2(n15950), .op(n15954) );
  nor3_1 U15744 ( .ip1(n16690), .ip2(n16497), .ip3(n15952), .op(n16018) );
  inv_1 U15745 ( .ip(n16018), .op(n15953) );
  nand2_1 U15746 ( .ip1(n15954), .ip2(n15953), .op(n16016) );
  xor2_1 U15747 ( .ip1(n15955), .ip2(n16016), .op(n16035) );
  nor3_1 U15748 ( .ip1(n16623), .ip2(n15973), .ip3(n15956), .op(n15957) );
  nor2_1 U15749 ( .ip1(n15958), .ip2(n15957), .op(n16034) );
  nor2_1 U15750 ( .ip1(n15960), .ip2(n15959), .op(n16033) );
  nor4_1 U15751 ( .ip1(n16496), .ip2(n16445), .ip3(n16596), .ip4(n16552), .op(
        n16029) );
  inv_1 U15752 ( .ip(n16029), .op(n15963) );
  nand2_1 U15753 ( .ip1(m2DataIn[4]), .ip2(q_w2[9]), .op(n16140) );
  nand2_1 U15754 ( .ip1(n16140), .ip2(n15961), .op(n15962) );
  nand2_1 U15755 ( .ip1(n15963), .ip2(n15962), .op(n15964) );
  nor3_1 U15756 ( .ip1(n16623), .ip2(n16144), .ip3(n15964), .op(n16028) );
  or2_1 U15757 ( .ip1(n15964), .ip2(n16028), .op(n15967) );
  nand2_1 U15758 ( .ip1(m2DataIn[12]), .ip2(q_w2[1]), .op(n15965) );
  or2_1 U15759 ( .ip1(n15965), .ip2(n16028), .op(n15966) );
  nand2_1 U15760 ( .ip1(n15967), .ip2(n15966), .op(n16065) );
  nand4_1 U15761 ( .ip1(m2DataIn[3]), .ip2(m2DataIn[0]), .ip3(q_w2[10]), .ip4(
        q_w2[13]), .op(n16050) );
  inv_1 U15762 ( .ip(n16050), .op(n15972) );
  or2_1 U15763 ( .ip1(q_w2[13]), .ip2(n15968), .op(n15970) );
  or2_1 U15764 ( .ip1(m2DataIn[0]), .ip2(n15968), .op(n15969) );
  nand2_1 U15765 ( .ip1(n15970), .ip2(n15969), .op(n15971) );
  nor2_1 U15766 ( .ip1(n15972), .ip2(n15971), .op(n16048) );
  inv_1 U15767 ( .ip(m2DataIn[13]), .op(n16510) );
  nor2_1 U15768 ( .ip1(n16510), .ip2(n15973), .op(n15974) );
  xor2_1 U15769 ( .ip1(n16048), .ip2(n15974), .op(n16064) );
  nor2_1 U15770 ( .ip1(n16550), .ip2(n16561), .op(n16104) );
  nand3_1 U15771 ( .ip1(m2DataIn[6]), .ip2(q_w2[6]), .ip3(n16104), .op(n16030)
         );
  nand2_1 U15772 ( .ip1(m2DataIn[6]), .ip2(q_w2[7]), .op(n16347) );
  nand2_1 U15773 ( .ip1(n16347), .ip2(n15975), .op(n15976) );
  nand2_1 U15774 ( .ip1(n16030), .ip2(n15976), .op(n15977) );
  nor3_1 U15775 ( .ip1(n16679), .ip2(n16308), .ip3(n15977), .op(n16031) );
  or2_1 U15776 ( .ip1(n15977), .ip2(n16031), .op(n15980) );
  nand2_1 U15777 ( .ip1(m2DataIn[11]), .ip2(q_w2[2]), .op(n15978) );
  or2_1 U15778 ( .ip1(n15978), .ip2(n16031), .op(n15979) );
  nand2_1 U15779 ( .ip1(n15980), .ip2(n15979), .op(n16063) );
  inv_1 U15780 ( .ip(n15981), .op(n16013) );
  nor2_1 U15781 ( .ip1(n15983), .ip2(n15982), .op(n16061) );
  inv_1 U15782 ( .ip(rdata[5]), .op(n16020) );
  nand2_1 U15783 ( .ip1(m2DataIn[2]), .ip2(q_w2[12]), .op(n16024) );
  nor3_1 U15784 ( .ip1(n16222), .ip2(n16599), .ip3(n16024), .op(n16022) );
  inv_1 U15785 ( .ip(n16022), .op(n15987) );
  nand2_1 U15786 ( .ip1(m2DataIn[1]), .ip2(q_w2[12]), .op(n15985) );
  nand2_1 U15787 ( .ip1(n15985), .ip2(n15984), .op(n15986) );
  nand2_1 U15788 ( .ip1(n15987), .ip2(n15986), .op(n16019) );
  mux2_1 U15789 ( .ip1(rdata[5]), .ip2(n16020), .s(n16019), .op(n16060) );
  nor2_1 U15790 ( .ip1(n15989), .ip2(n15988), .op(n15990) );
  nor2_1 U15791 ( .ip1(n15991), .ip2(n15990), .op(n16059) );
  fulladder U15792 ( .a(n15994), .b(n15993), .ci(n15992), .co(n16009), .s(
        n15933) );
  or2_1 U15793 ( .ip1(n15996), .ip2(n15995), .op(n15997) );
  nand2_1 U15794 ( .ip1(n15998), .ip2(n15997), .op(n15999) );
  nand2_1 U15795 ( .ip1(n16000), .ip2(n15999), .op(n16073) );
  or2_1 U15796 ( .ip1(n16000), .ip2(n15999), .op(n16070) );
  nand2_1 U15797 ( .ip1(n16073), .ip2(n16070), .op(n16001) );
  xor2_1 U15798 ( .ip1(n16071), .ip2(n16001), .op(n16005) );
  inv_1 U15799 ( .ip(\SIGMOID/lut_out [5]), .op(n16004) );
  or2_1 U15800 ( .ip1(\SIGMOID/lut_out [4]), .ip2(n16002), .op(n16078) );
  nand2_1 U15801 ( .ip1(n16164), .ip2(n16078), .op(n16003) );
  mux2_1 U15802 ( .ip1(n16004), .ip2(\SIGMOID/lut_out [5]), .s(n16003), .op(
        n17169) );
  mux2_1 U15803 ( .ip1(n16005), .ip2(n17169), .s(n16714), .op(n16007) );
  buf_1 U15804 ( .ip(n16007), .op(n16006) );
  mux2_1 U15805 ( .ip1(n16006), .ip2(\ANSWER/mem[0][0][5] ), .s(n16717), .op(
        n3402) );
  mux2_1 U15806 ( .ip1(n16006), .ip2(\ANSWER/mem[0][1][5] ), .s(n16718), .op(
        n3401) );
  mux2_1 U15807 ( .ip1(n16006), .ip2(\ANSWER/mem[0][2][5] ), .s(n16719), .op(
        n3400) );
  mux2_1 U15808 ( .ip1(n16006), .ip2(\ANSWER/mem[0][3][5] ), .s(n16720), .op(
        n3399) );
  mux2_1 U15809 ( .ip1(n16006), .ip2(\ANSWER/mem[0][4][5] ), .s(n16721), .op(
        n3398) );
  mux2_1 U15810 ( .ip1(n16006), .ip2(\ANSWER/mem[0][5][5] ), .s(n16722), .op(
        n3397) );
  mux2_1 U15811 ( .ip1(n16006), .ip2(\ANSWER/mem[0][6][5] ), .s(n16723), .op(
        n3396) );
  mux2_1 U15812 ( .ip1(n16006), .ip2(\ANSWER/mem[0][7][5] ), .s(n16724), .op(
        n3395) );
  mux2_1 U15813 ( .ip1(n16006), .ip2(\ANSWER/mem[0][8][5] ), .s(n16725), .op(
        n3394) );
  mux2_1 U15814 ( .ip1(n16006), .ip2(\ANSWER/mem[0][9][5] ), .s(n16726), .op(
        n3393) );
  mux2_1 U15815 ( .ip1(n16006), .ip2(\ANSWER/mem[1][0][5] ), .s(n16727), .op(
        n3392) );
  mux2_1 U15816 ( .ip1(n16006), .ip2(\ANSWER/mem[1][1][5] ), .s(n16728), .op(
        n3391) );
  mux2_1 U15817 ( .ip1(n16006), .ip2(\ANSWER/mem[1][2][5] ), .s(n16729), .op(
        n3390) );
  mux2_1 U15818 ( .ip1(n16006), .ip2(\ANSWER/mem[1][3][5] ), .s(n16730), .op(
        n3389) );
  mux2_1 U15819 ( .ip1(n16006), .ip2(\ANSWER/mem[1][4][5] ), .s(n16731), .op(
        n3388) );
  mux2_1 U15820 ( .ip1(n16006), .ip2(\ANSWER/mem[1][5][5] ), .s(n16732), .op(
        n3387) );
  mux2_1 U15821 ( .ip1(n16006), .ip2(\ANSWER/mem[1][6][5] ), .s(n16733), .op(
        n3386) );
  mux2_1 U15822 ( .ip1(n16006), .ip2(\ANSWER/mem[1][7][5] ), .s(n16734), .op(
        n3385) );
  mux2_1 U15823 ( .ip1(n16006), .ip2(\ANSWER/mem[1][8][5] ), .s(n16735), .op(
        n3384) );
  mux2_1 U15824 ( .ip1(n16006), .ip2(\ANSWER/mem[1][9][5] ), .s(n16736), .op(
        n3383) );
  mux2_1 U15825 ( .ip1(n16006), .ip2(\ANSWER/mem[2][0][5] ), .s(n16737), .op(
        n3382) );
  mux2_1 U15826 ( .ip1(n16006), .ip2(\ANSWER/mem[2][1][5] ), .s(n16738), .op(
        n3381) );
  mux2_1 U15827 ( .ip1(n16006), .ip2(\ANSWER/mem[2][2][5] ), .s(n16739), .op(
        n3380) );
  mux2_1 U15828 ( .ip1(n16006), .ip2(\ANSWER/mem[2][3][5] ), .s(n16740), .op(
        n3379) );
  mux2_1 U15829 ( .ip1(n16006), .ip2(\ANSWER/mem[2][4][5] ), .s(n16741), .op(
        n3378) );
  mux2_1 U15830 ( .ip1(n16006), .ip2(\ANSWER/mem[2][5][5] ), .s(n16742), .op(
        n3377) );
  mux2_1 U15831 ( .ip1(n16006), .ip2(\ANSWER/mem[2][6][5] ), .s(n16743), .op(
        n3376) );
  mux2_1 U15832 ( .ip1(n16006), .ip2(\ANSWER/mem[2][7][5] ), .s(n16744), .op(
        n3375) );
  mux2_1 U15833 ( .ip1(n16006), .ip2(\ANSWER/mem[2][8][5] ), .s(n16745), .op(
        n3374) );
  mux2_1 U15834 ( .ip1(n16006), .ip2(\ANSWER/mem[2][9][5] ), .s(n16746), .op(
        n3373) );
  mux2_1 U15835 ( .ip1(n16006), .ip2(\ANSWER/mem[3][0][5] ), .s(n16747), .op(
        n3372) );
  mux2_1 U15836 ( .ip1(n16006), .ip2(\ANSWER/mem[3][1][5] ), .s(n16748), .op(
        n3371) );
  mux2_1 U15837 ( .ip1(n16006), .ip2(\ANSWER/mem[3][2][5] ), .s(n16749), .op(
        n3370) );
  mux2_1 U15838 ( .ip1(n16006), .ip2(\ANSWER/mem[3][3][5] ), .s(n16750), .op(
        n3369) );
  mux2_1 U15839 ( .ip1(n16006), .ip2(\ANSWER/mem[3][4][5] ), .s(n16751), .op(
        n3368) );
  mux2_1 U15840 ( .ip1(n16006), .ip2(\ANSWER/mem[3][5][5] ), .s(n16752), .op(
        n3367) );
  mux2_1 U15841 ( .ip1(n16008), .ip2(\ANSWER/mem[3][6][5] ), .s(n16753), .op(
        n3366) );
  mux2_1 U15842 ( .ip1(n16008), .ip2(\ANSWER/mem[3][7][5] ), .s(n16754), .op(
        n3365) );
  mux2_1 U15843 ( .ip1(n16008), .ip2(\ANSWER/mem[3][8][5] ), .s(n16755), .op(
        n3364) );
  mux2_1 U15844 ( .ip1(n16008), .ip2(\ANSWER/mem[3][9][5] ), .s(n16756), .op(
        n3363) );
  mux2_1 U15845 ( .ip1(n16007), .ip2(\ANSWER/mem[4][0][5] ), .s(n16757), .op(
        n3362) );
  mux2_1 U15846 ( .ip1(n16007), .ip2(\ANSWER/mem[4][1][5] ), .s(n16758), .op(
        n3361) );
  mux2_1 U15847 ( .ip1(n16007), .ip2(\ANSWER/mem[4][2][5] ), .s(n16759), .op(
        n3360) );
  mux2_1 U15848 ( .ip1(n16007), .ip2(\ANSWER/mem[4][3][5] ), .s(n16760), .op(
        n3359) );
  mux2_1 U15849 ( .ip1(n16007), .ip2(\ANSWER/mem[4][4][5] ), .s(n16761), .op(
        n3358) );
  mux2_1 U15850 ( .ip1(n16007), .ip2(\ANSWER/mem[4][5][5] ), .s(n16762), .op(
        n3357) );
  mux2_1 U15851 ( .ip1(n16008), .ip2(\ANSWER/mem[4][6][5] ), .s(n16763), .op(
        n3356) );
  mux2_1 U15852 ( .ip1(n16008), .ip2(\ANSWER/mem[4][7][5] ), .s(n16764), .op(
        n3355) );
  mux2_1 U15853 ( .ip1(n16008), .ip2(\ANSWER/mem[4][8][5] ), .s(n16765), .op(
        n3354) );
  mux2_1 U15854 ( .ip1(n16008), .ip2(\ANSWER/mem[4][9][5] ), .s(n16766), .op(
        n3353) );
  mux2_1 U15855 ( .ip1(n16008), .ip2(\ANSWER/mem[5][0][5] ), .s(n16767), .op(
        n3352) );
  mux2_1 U15856 ( .ip1(n16007), .ip2(\ANSWER/mem[5][1][5] ), .s(n16768), .op(
        n3351) );
  mux2_1 U15857 ( .ip1(n16008), .ip2(\ANSWER/mem[5][2][5] ), .s(n16769), .op(
        n3350) );
  mux2_1 U15858 ( .ip1(n16007), .ip2(\ANSWER/mem[5][3][5] ), .s(n16770), .op(
        n3349) );
  mux2_1 U15859 ( .ip1(n16008), .ip2(\ANSWER/mem[5][4][5] ), .s(n16771), .op(
        n3348) );
  mux2_1 U15860 ( .ip1(n16007), .ip2(\ANSWER/mem[5][5][5] ), .s(n16772), .op(
        n3347) );
  mux2_1 U15861 ( .ip1(n16007), .ip2(\ANSWER/mem[5][6][5] ), .s(n16773), .op(
        n3346) );
  mux2_1 U15862 ( .ip1(n16007), .ip2(\ANSWER/mem[5][7][5] ), .s(n16774), .op(
        n3345) );
  mux2_1 U15863 ( .ip1(n16007), .ip2(\ANSWER/mem[5][8][5] ), .s(n16775), .op(
        n3344) );
  mux2_1 U15864 ( .ip1(n16007), .ip2(\ANSWER/mem[5][9][5] ), .s(n16776), .op(
        n3343) );
  mux2_1 U15865 ( .ip1(n16007), .ip2(\ANSWER/mem[6][0][5] ), .s(n16777), .op(
        n3342) );
  mux2_1 U15866 ( .ip1(n16007), .ip2(\ANSWER/mem[6][1][5] ), .s(n16778), .op(
        n3341) );
  mux2_1 U15867 ( .ip1(n16007), .ip2(\ANSWER/mem[6][2][5] ), .s(n16779), .op(
        n3340) );
  mux2_1 U15868 ( .ip1(n16007), .ip2(\ANSWER/mem[6][3][5] ), .s(n16780), .op(
        n3339) );
  mux2_1 U15869 ( .ip1(n16007), .ip2(\ANSWER/mem[6][4][5] ), .s(n16781), .op(
        n3338) );
  mux2_1 U15870 ( .ip1(n16007), .ip2(\ANSWER/mem[6][5][5] ), .s(n16782), .op(
        n3337) );
  mux2_1 U15871 ( .ip1(n16007), .ip2(\ANSWER/mem[6][6][5] ), .s(n16783), .op(
        n3336) );
  mux2_1 U15872 ( .ip1(n16007), .ip2(\ANSWER/mem[6][7][5] ), .s(n16784), .op(
        n3335) );
  mux2_1 U15873 ( .ip1(n16007), .ip2(\ANSWER/mem[6][8][5] ), .s(n16785), .op(
        n3334) );
  mux2_1 U15874 ( .ip1(n16007), .ip2(\ANSWER/mem[6][9][5] ), .s(n16786), .op(
        n3333) );
  mux2_1 U15875 ( .ip1(n16007), .ip2(\ANSWER/mem[7][0][5] ), .s(n16787), .op(
        n3332) );
  mux2_1 U15876 ( .ip1(n16007), .ip2(\ANSWER/mem[7][1][5] ), .s(n16788), .op(
        n3331) );
  buf_1 U15877 ( .ip(n16007), .op(n16008) );
  mux2_1 U15878 ( .ip1(n16008), .ip2(\ANSWER/mem[7][2][5] ), .s(n16790), .op(
        n3330) );
  mux2_1 U15879 ( .ip1(n16008), .ip2(\ANSWER/mem[7][3][5] ), .s(n16791), .op(
        n3329) );
  mux2_1 U15880 ( .ip1(n16008), .ip2(\ANSWER/mem[7][4][5] ), .s(n16792), .op(
        n3328) );
  mux2_1 U15881 ( .ip1(n16008), .ip2(\ANSWER/mem[7][5][5] ), .s(n16793), .op(
        n3327) );
  mux2_1 U15882 ( .ip1(n16008), .ip2(\ANSWER/mem[7][6][5] ), .s(n16794), .op(
        n3326) );
  mux2_1 U15883 ( .ip1(n16008), .ip2(\ANSWER/mem[7][7][5] ), .s(n16795), .op(
        n3325) );
  mux2_1 U15884 ( .ip1(n16008), .ip2(\ANSWER/mem[7][8][5] ), .s(n16796), .op(
        n3324) );
  mux2_1 U15885 ( .ip1(n16008), .ip2(\ANSWER/mem[7][9][5] ), .s(n16797), .op(
        n3323) );
  mux2_1 U15886 ( .ip1(n16008), .ip2(\ANSWER/mem[8][0][5] ), .s(n16798), .op(
        n3322) );
  mux2_1 U15887 ( .ip1(n16008), .ip2(\ANSWER/mem[8][1][5] ), .s(n16799), .op(
        n3321) );
  mux2_1 U15888 ( .ip1(n16008), .ip2(\ANSWER/mem[8][2][5] ), .s(n16800), .op(
        n3320) );
  mux2_1 U15889 ( .ip1(n16008), .ip2(\ANSWER/mem[8][3][5] ), .s(n16801), .op(
        n3319) );
  mux2_1 U15890 ( .ip1(n16007), .ip2(\ANSWER/mem[8][4][5] ), .s(n16803), .op(
        n3318) );
  mux2_1 U15891 ( .ip1(n16007), .ip2(\ANSWER/mem[8][5][5] ), .s(n16804), .op(
        n3317) );
  mux2_1 U15892 ( .ip1(n16007), .ip2(\ANSWER/mem[8][6][5] ), .s(n16805), .op(
        n3316) );
  mux2_1 U15893 ( .ip1(n16007), .ip2(\ANSWER/mem[8][7][5] ), .s(n16806), .op(
        n3315) );
  mux2_1 U15894 ( .ip1(n16007), .ip2(\ANSWER/mem[8][8][5] ), .s(n16807), .op(
        n3314) );
  mux2_1 U15895 ( .ip1(n16007), .ip2(\ANSWER/mem[8][9][5] ), .s(n16808), .op(
        n3313) );
  mux2_1 U15896 ( .ip1(n16007), .ip2(\ANSWER/mem[9][0][5] ), .s(n16809), .op(
        n3312) );
  mux2_1 U15897 ( .ip1(n16007), .ip2(\ANSWER/mem[9][1][5] ), .s(n16810), .op(
        n3311) );
  mux2_1 U15898 ( .ip1(n16007), .ip2(\ANSWER/mem[9][2][5] ), .s(n16811), .op(
        n3310) );
  mux2_1 U15899 ( .ip1(n16007), .ip2(\ANSWER/mem[9][3][5] ), .s(n16812), .op(
        n3309) );
  mux2_1 U15900 ( .ip1(n16007), .ip2(\ANSWER/mem[9][4][5] ), .s(n16813), .op(
        n3308) );
  mux2_1 U15901 ( .ip1(n16007), .ip2(\ANSWER/mem[9][5][5] ), .s(n16814), .op(
        n3307) );
  mux2_1 U15902 ( .ip1(n16008), .ip2(\ANSWER/mem[9][6][5] ), .s(n16815), .op(
        n3306) );
  mux2_1 U15903 ( .ip1(n16008), .ip2(\ANSWER/mem[9][7][5] ), .s(n16816), .op(
        n3305) );
  mux2_1 U15904 ( .ip1(n16008), .ip2(\ANSWER/mem[9][8][5] ), .s(n16817), .op(
        n3304) );
  mux2_1 U15905 ( .ip1(n16008), .ip2(\ANSWER/mem[9][9][5] ), .s(n16818), .op(
        n3303) );
  fulladder U15906 ( .a(n16011), .b(n16010), .ci(n16009), .co(n16077), .s(
        n16000) );
  inv_1 U15907 ( .ip(n16077), .op(n16155) );
  fulladder U15908 ( .a(n16014), .b(n16013), .ci(n16012), .co(n16015), .s(
        n16010) );
  inv_1 U15909 ( .ip(n16015), .op(n16154) );
  nor3_1 U15910 ( .ip1(n16600), .ip2(n16177), .ip3(n16016), .op(n16017) );
  nor2_1 U15911 ( .ip1(n16018), .ip2(n16017), .op(n16132) );
  nand2_1 U15912 ( .ip1(m2DataIn[11]), .ip2(q_w2[3]), .op(n16224) );
  nor2_1 U15913 ( .ip1(n16020), .ip2(n16019), .op(n16021) );
  nor2_1 U15914 ( .ip1(n16022), .ip2(n16021), .op(n16131) );
  nand2_1 U15915 ( .ip1(m2DataIn[1]), .ip2(q_w2[13]), .op(n16092) );
  nand4_1 U15916 ( .ip1(m2DataIn[2]), .ip2(m2DataIn[1]), .ip3(q_w2[12]), .ip4(
        q_w2[13]), .op(n16125) );
  inv_1 U15917 ( .ip(n16125), .op(n16023) );
  or2_1 U15918 ( .ip1(n16092), .ip2(n16023), .op(n16026) );
  or2_1 U15919 ( .ip1(n16024), .ip2(n16023), .op(n16025) );
  nand2_1 U15920 ( .ip1(n16026), .ip2(n16025), .op(n16123) );
  mux2_1 U15921 ( .ip1(n16027), .ip2(rdata[6]), .s(n16123), .op(n16130) );
  nor2_1 U15922 ( .ip1(n16029), .ip2(n16028), .op(n16129) );
  inv_1 U15923 ( .ip(n16030), .op(n16032) );
  nor2_1 U15924 ( .ip1(n16032), .ip2(n16031), .op(n16128) );
  fulladder U15925 ( .a(n16035), .b(n16034), .ci(n16033), .co(n16137), .s(
        n16014) );
  inv_1 U15926 ( .ip(n16036), .op(n16153) );
  fulladder U15927 ( .a(n16039), .b(n16038), .ci(n16037), .co(n16152), .s(
        n15946) );
  inv_1 U15928 ( .ip(n16040), .op(n16087) );
  nor2_1 U15929 ( .ip1(n16600), .ip2(n16497), .op(n16185) );
  and3_1 U15930 ( .ip1(m2DataIn[9]), .ip2(q_w2[4]), .ip3(n16185), .op(n16099)
         );
  nor2_1 U15931 ( .ip1(n16690), .ip2(n16497), .op(n16041) );
  or2_1 U15932 ( .ip1(q_w2[4]), .ip2(n16041), .op(n16043) );
  or2_1 U15933 ( .ip1(m2DataIn[10]), .ip2(n16041), .op(n16042) );
  nand2_1 U15934 ( .ip1(n16043), .ip2(n16042), .op(n16044) );
  nor2_1 U15935 ( .ip1(n16099), .ip2(n16044), .op(n16098) );
  nor2_1 U15936 ( .ip1(n16623), .ip2(n16308), .op(n16100) );
  xor2_1 U15937 ( .ip1(n16098), .ip2(n16100), .op(n16122) );
  nor4_1 U15938 ( .ip1(n16550), .ip2(n16273), .ip3(n16561), .ip4(n16596), .op(
        n16115) );
  or2_1 U15939 ( .ip1(q_w2[8]), .ip2(n16104), .op(n16046) );
  or2_1 U15940 ( .ip1(m2DataIn[6]), .ip2(n16104), .op(n16045) );
  nand2_1 U15941 ( .ip1(n16046), .ip2(n16045), .op(n16047) );
  nor2_1 U15942 ( .ip1(n16115), .ip2(n16047), .op(n16114) );
  nor2_1 U15943 ( .ip1(n16510), .ip2(n16144), .op(n16116) );
  xor2_1 U15944 ( .ip1(n16114), .ip2(n16116), .op(n16121) );
  nand3_1 U15945 ( .ip1(m2DataIn[13]), .ip2(q_w2[0]), .ip3(n16048), .op(n16049) );
  nand2_1 U15946 ( .ip1(n16050), .ip2(n16049), .op(n16120) );
  nand2_1 U15947 ( .ip1(m2DataIn[5]), .ip2(q_w2[9]), .op(n16051) );
  nor3_1 U15948 ( .ip1(n16496), .ip2(n16622), .ip3(n16140), .op(n16110) );
  or2_1 U15949 ( .ip1(n16051), .ip2(n16110), .op(n16054) );
  nand2_1 U15950 ( .ip1(m2DataIn[4]), .ip2(q_w2[10]), .op(n16052) );
  or2_1 U15951 ( .ip1(n16052), .ip2(n16110), .op(n16053) );
  nand2_1 U15952 ( .ip1(n16054), .ip2(n16053), .op(n16109) );
  nor2_1 U15953 ( .ip1(n16624), .ip2(n16538), .op(n16111) );
  xnor2_1 U15954 ( .ip1(n16109), .ip2(n16111), .op(n16150) );
  nand2_1 U15955 ( .ip1(m2DataIn[3]), .ip2(q_w2[14]), .op(n16352) );
  nor3_1 U15956 ( .ip1(n16145), .ip2(n16599), .ip3(n16352), .op(n16091) );
  or2_1 U15957 ( .ip1(q_w2[14]), .ip2(n16055), .op(n16057) );
  or2_1 U15958 ( .ip1(m2DataIn[0]), .ip2(n16055), .op(n16056) );
  nand2_1 U15959 ( .ip1(n16057), .ip2(n16056), .op(n16089) );
  nor2_1 U15960 ( .ip1(n16091), .ip2(n16089), .op(n16058) );
  nand2_1 U15961 ( .ip1(m2DataIn[14]), .ip2(q_w2[0]), .op(n16088) );
  xor2_1 U15962 ( .ip1(n16058), .ip2(n16088), .op(n16149) );
  fulladder U15963 ( .a(n16061), .b(n16060), .ci(n16059), .co(n16148), .s(
        n16012) );
  inv_1 U15964 ( .ip(n16062), .op(n16135) );
  fulladder U15965 ( .a(n16065), .b(n16064), .ci(n16063), .co(n16134), .s(
        n15981) );
  inv_1 U15966 ( .ip(n16066), .op(n16086) );
  fulladder U15967 ( .a(n16069), .b(n16068), .ci(n16067), .co(n16085), .s(
        n16011) );
  nand2_1 U15968 ( .ip1(n16071), .ip2(n16070), .op(n16072) );
  nand2_1 U15969 ( .ip1(n16073), .ip2(n16072), .op(n16074) );
  or2_1 U15970 ( .ip1(n16075), .ip2(n16074), .op(n16158) );
  nand2_1 U15971 ( .ip1(n16075), .ip2(n16074), .op(n16156) );
  nand2_1 U15972 ( .ip1(n16158), .ip2(n16156), .op(n16076) );
  mux2_1 U15973 ( .ip1(n16077), .ip2(n16155), .s(n16076), .op(n16081) );
  inv_1 U15974 ( .ip(\SIGMOID/lut_out [6]), .op(n16080) );
  or2_1 U15975 ( .ip1(\SIGMOID/lut_out [5]), .ip2(n16078), .op(n16163) );
  nand2_1 U15976 ( .ip1(n16164), .ip2(n16163), .op(n16079) );
  mux2_1 U15977 ( .ip1(n16080), .ip2(\SIGMOID/lut_out [6]), .s(n16079), .op(
        n17201) );
  mux2_1 U15978 ( .ip1(n16081), .ip2(n17201), .s(n16714), .op(n16082) );
  buf_1 U15979 ( .ip(n16082), .op(n16083) );
  mux2_1 U15980 ( .ip1(n16083), .ip2(\ANSWER/mem[0][0][6] ), .s(n16717), .op(
        n3302) );
  mux2_1 U15981 ( .ip1(n16083), .ip2(\ANSWER/mem[0][1][6] ), .s(n16718), .op(
        n3301) );
  mux2_1 U15982 ( .ip1(n16083), .ip2(\ANSWER/mem[0][2][6] ), .s(n16719), .op(
        n3300) );
  mux2_1 U15983 ( .ip1(n16083), .ip2(\ANSWER/mem[0][3][6] ), .s(n16720), .op(
        n3299) );
  mux2_1 U15984 ( .ip1(n16083), .ip2(\ANSWER/mem[0][4][6] ), .s(n16721), .op(
        n3298) );
  mux2_1 U15985 ( .ip1(n16083), .ip2(\ANSWER/mem[0][5][6] ), .s(n16722), .op(
        n3297) );
  mux2_1 U15986 ( .ip1(n16083), .ip2(\ANSWER/mem[0][6][6] ), .s(n16723), .op(
        n3296) );
  mux2_1 U15987 ( .ip1(n16083), .ip2(\ANSWER/mem[0][7][6] ), .s(n16724), .op(
        n3295) );
  mux2_1 U15988 ( .ip1(n16083), .ip2(\ANSWER/mem[0][8][6] ), .s(n16725), .op(
        n3294) );
  mux2_1 U15989 ( .ip1(n16083), .ip2(\ANSWER/mem[0][9][6] ), .s(n16726), .op(
        n3293) );
  mux2_1 U15990 ( .ip1(n16083), .ip2(\ANSWER/mem[1][0][6] ), .s(n16727), .op(
        n3292) );
  mux2_1 U15991 ( .ip1(n16083), .ip2(\ANSWER/mem[1][1][6] ), .s(n16728), .op(
        n3291) );
  buf_1 U15992 ( .ip(n16082), .op(n16084) );
  mux2_1 U15993 ( .ip1(n16084), .ip2(\ANSWER/mem[1][2][6] ), .s(n16729), .op(
        n3290) );
  mux2_1 U15994 ( .ip1(n16084), .ip2(\ANSWER/mem[1][3][6] ), .s(n16730), .op(
        n3289) );
  mux2_1 U15995 ( .ip1(n16082), .ip2(\ANSWER/mem[1][4][6] ), .s(n16731), .op(
        n3288) );
  mux2_1 U15996 ( .ip1(n16082), .ip2(\ANSWER/mem[1][5][6] ), .s(n16732), .op(
        n3287) );
  mux2_1 U15997 ( .ip1(n16082), .ip2(\ANSWER/mem[1][6][6] ), .s(n16733), .op(
        n3286) );
  mux2_1 U15998 ( .ip1(n16082), .ip2(\ANSWER/mem[1][7][6] ), .s(n16734), .op(
        n3285) );
  mux2_1 U15999 ( .ip1(n16082), .ip2(\ANSWER/mem[1][8][6] ), .s(n16735), .op(
        n3284) );
  mux2_1 U16000 ( .ip1(n16082), .ip2(\ANSWER/mem[1][9][6] ), .s(n16736), .op(
        n3283) );
  mux2_1 U16001 ( .ip1(n16082), .ip2(\ANSWER/mem[2][0][6] ), .s(n16737), .op(
        n3282) );
  mux2_1 U16002 ( .ip1(n16082), .ip2(\ANSWER/mem[2][1][6] ), .s(n16738), .op(
        n3281) );
  mux2_1 U16003 ( .ip1(n16082), .ip2(\ANSWER/mem[2][2][6] ), .s(n16739), .op(
        n3280) );
  mux2_1 U16004 ( .ip1(n16082), .ip2(\ANSWER/mem[2][3][6] ), .s(n16740), .op(
        n3279) );
  mux2_1 U16005 ( .ip1(n16084), .ip2(\ANSWER/mem[2][4][6] ), .s(n16741), .op(
        n3278) );
  mux2_1 U16006 ( .ip1(n16083), .ip2(\ANSWER/mem[2][5][6] ), .s(n16742), .op(
        n3277) );
  mux2_1 U16007 ( .ip1(n16083), .ip2(\ANSWER/mem[2][6][6] ), .s(n16743), .op(
        n3276) );
  mux2_1 U16008 ( .ip1(n16082), .ip2(\ANSWER/mem[2][7][6] ), .s(n16744), .op(
        n3275) );
  mux2_1 U16009 ( .ip1(n16084), .ip2(\ANSWER/mem[2][8][6] ), .s(n16745), .op(
        n3274) );
  mux2_1 U16010 ( .ip1(n16083), .ip2(\ANSWER/mem[2][9][6] ), .s(n16746), .op(
        n3273) );
  mux2_1 U16011 ( .ip1(n16084), .ip2(\ANSWER/mem[3][0][6] ), .s(n16747), .op(
        n3272) );
  mux2_1 U16012 ( .ip1(n16082), .ip2(\ANSWER/mem[3][1][6] ), .s(n16748), .op(
        n3271) );
  mux2_1 U16013 ( .ip1(n16082), .ip2(\ANSWER/mem[3][2][6] ), .s(n16749), .op(
        n3270) );
  mux2_1 U16014 ( .ip1(n16082), .ip2(\ANSWER/mem[3][3][6] ), .s(n16750), .op(
        n3269) );
  mux2_1 U16015 ( .ip1(n16082), .ip2(\ANSWER/mem[3][4][6] ), .s(n16751), .op(
        n3268) );
  mux2_1 U16016 ( .ip1(n16082), .ip2(\ANSWER/mem[3][5][6] ), .s(n16752), .op(
        n3267) );
  mux2_1 U16017 ( .ip1(n16084), .ip2(\ANSWER/mem[3][6][6] ), .s(n16753), .op(
        n3266) );
  mux2_1 U16018 ( .ip1(n16084), .ip2(\ANSWER/mem[3][7][6] ), .s(n16754), .op(
        n3265) );
  mux2_1 U16019 ( .ip1(n16084), .ip2(\ANSWER/mem[3][8][6] ), .s(n16755), .op(
        n3264) );
  mux2_1 U16020 ( .ip1(n16084), .ip2(\ANSWER/mem[3][9][6] ), .s(n16756), .op(
        n3263) );
  mux2_1 U16021 ( .ip1(n16084), .ip2(\ANSWER/mem[4][0][6] ), .s(n16757), .op(
        n3262) );
  mux2_1 U16022 ( .ip1(n16084), .ip2(\ANSWER/mem[4][1][6] ), .s(n16758), .op(
        n3261) );
  mux2_1 U16023 ( .ip1(n16083), .ip2(\ANSWER/mem[4][2][6] ), .s(n16759), .op(
        n3260) );
  mux2_1 U16024 ( .ip1(n16082), .ip2(\ANSWER/mem[4][3][6] ), .s(n16760), .op(
        n3259) );
  mux2_1 U16025 ( .ip1(n16084), .ip2(\ANSWER/mem[4][4][6] ), .s(n16761), .op(
        n3258) );
  mux2_1 U16026 ( .ip1(n16084), .ip2(\ANSWER/mem[4][5][6] ), .s(n16762), .op(
        n3257) );
  mux2_1 U16027 ( .ip1(n16082), .ip2(\ANSWER/mem[4][6][6] ), .s(n16763), .op(
        n3256) );
  mux2_1 U16028 ( .ip1(n16084), .ip2(\ANSWER/mem[4][7][6] ), .s(n16764), .op(
        n3255) );
  mux2_1 U16029 ( .ip1(n16084), .ip2(\ANSWER/mem[4][8][6] ), .s(n16765), .op(
        n3254) );
  mux2_1 U16030 ( .ip1(n16082), .ip2(\ANSWER/mem[4][9][6] ), .s(n16766), .op(
        n3253) );
  mux2_1 U16031 ( .ip1(n16082), .ip2(\ANSWER/mem[5][0][6] ), .s(n16767), .op(
        n3252) );
  mux2_1 U16032 ( .ip1(n16084), .ip2(\ANSWER/mem[5][1][6] ), .s(n16768), .op(
        n3251) );
  mux2_1 U16033 ( .ip1(n16082), .ip2(\ANSWER/mem[5][2][6] ), .s(n16769), .op(
        n3250) );
  mux2_1 U16034 ( .ip1(n16082), .ip2(\ANSWER/mem[5][3][6] ), .s(n16770), .op(
        n3249) );
  mux2_1 U16035 ( .ip1(n16084), .ip2(\ANSWER/mem[5][4][6] ), .s(n16771), .op(
        n3248) );
  mux2_1 U16036 ( .ip1(n16082), .ip2(\ANSWER/mem[5][5][6] ), .s(n16772), .op(
        n3247) );
  mux2_1 U16037 ( .ip1(n16082), .ip2(\ANSWER/mem[5][6][6] ), .s(n16773), .op(
        n3246) );
  mux2_1 U16038 ( .ip1(n16084), .ip2(\ANSWER/mem[5][7][6] ), .s(n16774), .op(
        n3245) );
  mux2_1 U16039 ( .ip1(n16082), .ip2(\ANSWER/mem[5][8][6] ), .s(n16775), .op(
        n3244) );
  mux2_1 U16040 ( .ip1(n16082), .ip2(\ANSWER/mem[5][9][6] ), .s(n16776), .op(
        n3243) );
  mux2_1 U16041 ( .ip1(n16083), .ip2(\ANSWER/mem[6][0][6] ), .s(n16777), .op(
        n3242) );
  mux2_1 U16042 ( .ip1(n16083), .ip2(\ANSWER/mem[6][1][6] ), .s(n16778), .op(
        n3241) );
  mux2_1 U16043 ( .ip1(n16084), .ip2(\ANSWER/mem[6][2][6] ), .s(n16779), .op(
        n3240) );
  mux2_1 U16044 ( .ip1(n16082), .ip2(\ANSWER/mem[6][3][6] ), .s(n16780), .op(
        n3239) );
  mux2_1 U16045 ( .ip1(n16082), .ip2(\ANSWER/mem[6][4][6] ), .s(n16781), .op(
        n3238) );
  mux2_1 U16046 ( .ip1(n16084), .ip2(\ANSWER/mem[6][5][6] ), .s(n16782), .op(
        n3237) );
  mux2_1 U16047 ( .ip1(n16083), .ip2(\ANSWER/mem[6][6][6] ), .s(n16783), .op(
        n3236) );
  mux2_1 U16048 ( .ip1(n16083), .ip2(\ANSWER/mem[6][7][6] ), .s(n16784), .op(
        n3235) );
  mux2_1 U16049 ( .ip1(n16083), .ip2(\ANSWER/mem[6][8][6] ), .s(n16785), .op(
        n3234) );
  mux2_1 U16050 ( .ip1(n16084), .ip2(\ANSWER/mem[6][9][6] ), .s(n16786), .op(
        n3233) );
  mux2_1 U16051 ( .ip1(n16082), .ip2(\ANSWER/mem[7][0][6] ), .s(n16787), .op(
        n3232) );
  mux2_1 U16052 ( .ip1(n16082), .ip2(\ANSWER/mem[7][1][6] ), .s(n16788), .op(
        n3231) );
  mux2_1 U16053 ( .ip1(n16082), .ip2(\ANSWER/mem[7][2][6] ), .s(n16790), .op(
        n3230) );
  mux2_1 U16054 ( .ip1(n16082), .ip2(\ANSWER/mem[7][3][6] ), .s(n16791), .op(
        n3229) );
  mux2_1 U16055 ( .ip1(n16082), .ip2(\ANSWER/mem[7][4][6] ), .s(n16792), .op(
        n3228) );
  mux2_1 U16056 ( .ip1(n16082), .ip2(\ANSWER/mem[7][5][6] ), .s(n16793), .op(
        n3227) );
  mux2_1 U16057 ( .ip1(n16082), .ip2(\ANSWER/mem[7][6][6] ), .s(n16794), .op(
        n3226) );
  mux2_1 U16058 ( .ip1(n16082), .ip2(\ANSWER/mem[7][7][6] ), .s(n16795), .op(
        n3225) );
  mux2_1 U16059 ( .ip1(n16082), .ip2(\ANSWER/mem[7][8][6] ), .s(n16796), .op(
        n3224) );
  mux2_1 U16060 ( .ip1(n16083), .ip2(\ANSWER/mem[7][9][6] ), .s(n16797), .op(
        n3223) );
  mux2_1 U16061 ( .ip1(n16083), .ip2(\ANSWER/mem[8][0][6] ), .s(n16798), .op(
        n3222) );
  mux2_1 U16062 ( .ip1(n16084), .ip2(\ANSWER/mem[8][1][6] ), .s(n16799), .op(
        n3221) );
  mux2_1 U16063 ( .ip1(n16083), .ip2(\ANSWER/mem[8][2][6] ), .s(n16800), .op(
        n3220) );
  mux2_1 U16064 ( .ip1(n16084), .ip2(\ANSWER/mem[8][3][6] ), .s(n16801), .op(
        n3219) );
  mux2_1 U16065 ( .ip1(n16083), .ip2(\ANSWER/mem[8][4][6] ), .s(n16803), .op(
        n3218) );
  mux2_1 U16066 ( .ip1(n16082), .ip2(\ANSWER/mem[8][5][6] ), .s(n16804), .op(
        n3217) );
  mux2_1 U16067 ( .ip1(n16084), .ip2(\ANSWER/mem[8][6][6] ), .s(n16805), .op(
        n3216) );
  mux2_1 U16068 ( .ip1(n16083), .ip2(\ANSWER/mem[8][7][6] ), .s(n16806), .op(
        n3215) );
  mux2_1 U16069 ( .ip1(n16084), .ip2(\ANSWER/mem[8][8][6] ), .s(n16807), .op(
        n3214) );
  mux2_1 U16070 ( .ip1(n16083), .ip2(\ANSWER/mem[8][9][6] ), .s(n16808), .op(
        n3213) );
  mux2_1 U16071 ( .ip1(n16084), .ip2(\ANSWER/mem[9][0][6] ), .s(n16809), .op(
        n3212) );
  mux2_1 U16072 ( .ip1(n16083), .ip2(\ANSWER/mem[9][1][6] ), .s(n16810), .op(
        n3211) );
  mux2_1 U16073 ( .ip1(n16084), .ip2(\ANSWER/mem[9][2][6] ), .s(n16811), .op(
        n3210) );
  mux2_1 U16074 ( .ip1(n16083), .ip2(\ANSWER/mem[9][3][6] ), .s(n16812), .op(
        n3209) );
  mux2_1 U16075 ( .ip1(n16084), .ip2(\ANSWER/mem[9][4][6] ), .s(n16813), .op(
        n3208) );
  mux2_1 U16076 ( .ip1(n16083), .ip2(\ANSWER/mem[9][5][6] ), .s(n16814), .op(
        n3207) );
  mux2_1 U16077 ( .ip1(n16084), .ip2(\ANSWER/mem[9][6][6] ), .s(n16815), .op(
        n3206) );
  mux2_1 U16078 ( .ip1(n16084), .ip2(\ANSWER/mem[9][7][6] ), .s(n16816), .op(
        n3205) );
  mux2_1 U16079 ( .ip1(n16084), .ip2(\ANSWER/mem[9][8][6] ), .s(n16817), .op(
        n3204) );
  mux2_1 U16080 ( .ip1(n16084), .ip2(\ANSWER/mem[9][9][6] ), .s(n16818), .op(
        n3203) );
  fulladder U16081 ( .a(n16087), .b(n16086), .ci(n16085), .co(n16242), .s(
        n16075) );
  nor2_1 U16082 ( .ip1(n16089), .ip2(n16088), .op(n16090) );
  nor2_1 U16083 ( .ip1(n16091), .ip2(n16090), .op(n16217) );
  inv_1 U16084 ( .ip(rdata[7]), .op(n16097) );
  nand2_1 U16085 ( .ip1(m2DataIn[2]), .ip2(q_w2[13]), .op(n16093) );
  inv_1 U16086 ( .ip(q_w2[14]), .op(n16689) );
  nor3_1 U16087 ( .ip1(n16309), .ip2(n16689), .ip3(n16092), .op(n16208) );
  or2_1 U16088 ( .ip1(n16093), .ip2(n16208), .op(n16096) );
  nand2_1 U16089 ( .ip1(m2DataIn[1]), .ip2(q_w2[14]), .op(n16094) );
  or2_1 U16090 ( .ip1(n16094), .ip2(n16208), .op(n16095) );
  nand2_1 U16091 ( .ip1(n16096), .ip2(n16095), .op(n16209) );
  mux2_1 U16092 ( .ip1(n16097), .ip2(rdata[7]), .s(n16209), .op(n16216) );
  or2_1 U16093 ( .ip1(n16098), .ip2(n16099), .op(n16102) );
  or2_1 U16094 ( .ip1(n16100), .ip2(n16099), .op(n16101) );
  nand2_1 U16095 ( .ip1(n16102), .ip2(n16101), .op(n16215) );
  inv_1 U16096 ( .ip(n16103), .op(n16233) );
  nor2_1 U16097 ( .ip1(n16624), .ip2(n16596), .op(n16413) );
  and2_1 U16098 ( .ip1(n16104), .ip2(n16413), .op(n16207) );
  nor2_1 U16099 ( .ip1(n16550), .ip2(n16596), .op(n16105) );
  or2_1 U16100 ( .ip1(q_w2[7]), .ip2(n16105), .op(n16107) );
  or2_1 U16101 ( .ip1(m2DataIn[8]), .ip2(n16105), .op(n16106) );
  nand2_1 U16102 ( .ip1(n16107), .ip2(n16106), .op(n16205) );
  nor2_1 U16103 ( .ip1(n16207), .ip2(n16205), .op(n16108) );
  nand2_1 U16104 ( .ip1(m2DataIn[13]), .ip2(q_w2[2]), .op(n16204) );
  xor2_1 U16105 ( .ip1(n16108), .ip2(n16204), .op(n16214) );
  or2_1 U16106 ( .ip1(n16109), .ip2(n16110), .op(n16113) );
  or2_1 U16107 ( .ip1(n16111), .ip2(n16110), .op(n16112) );
  nand2_1 U16108 ( .ip1(n16113), .ip2(n16112), .op(n16213) );
  or2_1 U16109 ( .ip1(n16114), .ip2(n16115), .op(n16118) );
  or2_1 U16110 ( .ip1(n16116), .ip2(n16115), .op(n16117) );
  nand2_1 U16111 ( .ip1(n16118), .ip2(n16117), .op(n16212) );
  inv_1 U16112 ( .ip(n16119), .op(n16232) );
  fulladder U16113 ( .a(n16122), .b(n16121), .ci(n16120), .co(n16231), .s(
        n16136) );
  nand2_1 U16114 ( .ip1(rdata[6]), .ip2(n16123), .op(n16124) );
  nand2_1 U16115 ( .ip1(n16125), .ip2(n16124), .op(n16226) );
  nand2_1 U16116 ( .ip1(q_w2[4]), .ip2(m2DataIn[11]), .op(n16127) );
  nor2_1 U16117 ( .ip1(n16177), .ip2(n16623), .op(n16126) );
  xor2_1 U16118 ( .ip1(n16127), .ip2(n16126), .op(n16225) );
  xor2_1 U16119 ( .ip1(n16226), .ip2(n16225), .op(n16237) );
  fulladder U16120 ( .a(n16130), .b(n16129), .ci(n16128), .co(n16236), .s(
        n16138) );
  fulladder U16121 ( .a(n16132), .b(n16224), .ci(n16131), .co(n16235), .s(
        n16139) );
  inv_1 U16122 ( .ip(n16133), .op(n16240) );
  fulladder U16123 ( .a(n16136), .b(n16135), .ci(n16134), .co(n16239), .s(
        n16066) );
  fulladder U16124 ( .a(n16139), .b(n16138), .ci(n16137), .co(n16220), .s(
        n16036) );
  nor2_1 U16125 ( .ip1(n16496), .ip2(n16622), .op(n16184) );
  nand2_1 U16126 ( .ip1(m2DataIn[15]), .ip2(q_w2[0]), .op(n16183) );
  nor3_1 U16127 ( .ip1(n16273), .ip2(n16599), .ip3(n16140), .op(n16187) );
  nor2_1 U16128 ( .ip1(n16273), .ip2(n16552), .op(n16178) );
  or2_1 U16129 ( .ip1(q_w2[11]), .ip2(n16178), .op(n16142) );
  or2_1 U16130 ( .ip1(m2DataIn[4]), .ip2(n16178), .op(n16141) );
  nand2_1 U16131 ( .ip1(n16142), .ip2(n16141), .op(n16143) );
  nor2_1 U16132 ( .ip1(n16187), .ip2(n16143), .op(n16186) );
  inv_1 U16133 ( .ip(m2DataIn[14]), .op(n16597) );
  nor2_1 U16134 ( .ip1(n16597), .ip2(n16144), .op(n16188) );
  xor2_1 U16135 ( .ip1(n16186), .ip2(n16188), .op(n16201) );
  inv_1 U16136 ( .ip(q_w2[15]), .op(n16495) );
  nor2_1 U16137 ( .ip1(n16145), .ip2(n16495), .op(n16198) );
  nand2_1 U16138 ( .ip1(m2DataIn[9]), .ip2(q_w2[6]), .op(n16196) );
  inv_1 U16139 ( .ip(n16146), .op(n16200) );
  inv_1 U16140 ( .ip(n16147), .op(n16219) );
  fulladder U16141 ( .a(n16150), .b(n16149), .ci(n16148), .co(n16218), .s(
        n16062) );
  inv_1 U16142 ( .ip(n16151), .op(n16172) );
  fulladder U16143 ( .a(n16154), .b(n16153), .ci(n16152), .co(n16171), .s(
        n16040) );
  nand2_1 U16144 ( .ip1(n16156), .ip2(n16155), .op(n16157) );
  nand2_1 U16145 ( .ip1(n16158), .ip2(n16157), .op(n16159) );
  nand2_1 U16146 ( .ip1(n16160), .ip2(n16159), .op(n16245) );
  nor2_1 U16147 ( .ip1(n16160), .ip2(n16159), .op(n16243) );
  inv_1 U16148 ( .ip(n16243), .op(n16161) );
  nand2_1 U16149 ( .ip1(n16245), .ip2(n16161), .op(n16162) );
  xor2_1 U16150 ( .ip1(n16242), .ip2(n16162), .op(n16167) );
  inv_1 U16151 ( .ip(\SIGMOID/lut_out [7]), .op(n16166) );
  or2_1 U16152 ( .ip1(\SIGMOID/lut_out [6]), .ip2(n16163), .op(n16250) );
  nand2_1 U16153 ( .ip1(n16164), .ip2(n16250), .op(n16165) );
  mux2_1 U16154 ( .ip1(n16166), .ip2(\SIGMOID/lut_out [7]), .s(n16165), .op(
        n17242) );
  mux2_1 U16155 ( .ip1(n16167), .ip2(n17242), .s(n16714), .op(n16169) );
  buf_1 U16156 ( .ip(n16169), .op(n16168) );
  mux2_1 U16157 ( .ip1(n16168), .ip2(\ANSWER/mem[0][0][7] ), .s(n16717), .op(
        n3202) );
  mux2_1 U16158 ( .ip1(n16168), .ip2(\ANSWER/mem[0][1][7] ), .s(n16718), .op(
        n3201) );
  mux2_1 U16159 ( .ip1(n16168), .ip2(\ANSWER/mem[0][2][7] ), .s(n16719), .op(
        n3200) );
  mux2_1 U16160 ( .ip1(n16168), .ip2(\ANSWER/mem[0][3][7] ), .s(n16720), .op(
        n3199) );
  mux2_1 U16161 ( .ip1(n16168), .ip2(\ANSWER/mem[0][4][7] ), .s(n16721), .op(
        n3198) );
  mux2_1 U16162 ( .ip1(n16168), .ip2(\ANSWER/mem[0][5][7] ), .s(n16722), .op(
        n3197) );
  mux2_1 U16163 ( .ip1(n16168), .ip2(\ANSWER/mem[0][6][7] ), .s(n16723), .op(
        n3196) );
  mux2_1 U16164 ( .ip1(n16168), .ip2(\ANSWER/mem[0][7][7] ), .s(n16724), .op(
        n3195) );
  mux2_1 U16165 ( .ip1(n16168), .ip2(\ANSWER/mem[0][8][7] ), .s(n16725), .op(
        n3194) );
  mux2_1 U16166 ( .ip1(n16168), .ip2(\ANSWER/mem[0][9][7] ), .s(n16726), .op(
        n3193) );
  mux2_1 U16167 ( .ip1(n16168), .ip2(\ANSWER/mem[1][0][7] ), .s(n16727), .op(
        n3192) );
  mux2_1 U16168 ( .ip1(n16168), .ip2(\ANSWER/mem[1][1][7] ), .s(n16728), .op(
        n3191) );
  mux2_1 U16169 ( .ip1(n16168), .ip2(\ANSWER/mem[1][2][7] ), .s(n16729), .op(
        n3190) );
  mux2_1 U16170 ( .ip1(n16168), .ip2(\ANSWER/mem[1][3][7] ), .s(n16730), .op(
        n3189) );
  mux2_1 U16171 ( .ip1(n16168), .ip2(\ANSWER/mem[1][4][7] ), .s(n16731), .op(
        n3188) );
  mux2_1 U16172 ( .ip1(n16168), .ip2(\ANSWER/mem[1][5][7] ), .s(n16732), .op(
        n3187) );
  mux2_1 U16173 ( .ip1(n16168), .ip2(\ANSWER/mem[1][6][7] ), .s(n16733), .op(
        n3186) );
  mux2_1 U16174 ( .ip1(n16168), .ip2(\ANSWER/mem[1][7][7] ), .s(n16734), .op(
        n3185) );
  mux2_1 U16175 ( .ip1(n16168), .ip2(\ANSWER/mem[1][8][7] ), .s(n16735), .op(
        n3184) );
  mux2_1 U16176 ( .ip1(n16168), .ip2(\ANSWER/mem[1][9][7] ), .s(n16736), .op(
        n3183) );
  mux2_1 U16177 ( .ip1(n16168), .ip2(\ANSWER/mem[2][0][7] ), .s(n16737), .op(
        n3182) );
  mux2_1 U16178 ( .ip1(n16168), .ip2(\ANSWER/mem[2][1][7] ), .s(n16738), .op(
        n3181) );
  mux2_1 U16179 ( .ip1(n16168), .ip2(\ANSWER/mem[2][2][7] ), .s(n16739), .op(
        n3180) );
  mux2_1 U16180 ( .ip1(n16168), .ip2(\ANSWER/mem[2][3][7] ), .s(n16740), .op(
        n3179) );
  mux2_1 U16181 ( .ip1(n16168), .ip2(\ANSWER/mem[2][4][7] ), .s(n16741), .op(
        n3178) );
  mux2_1 U16182 ( .ip1(n16168), .ip2(\ANSWER/mem[2][5][7] ), .s(n16742), .op(
        n3177) );
  mux2_1 U16183 ( .ip1(n16168), .ip2(\ANSWER/mem[2][6][7] ), .s(n16743), .op(
        n3176) );
  mux2_1 U16184 ( .ip1(n16168), .ip2(\ANSWER/mem[2][7][7] ), .s(n16744), .op(
        n3175) );
  mux2_1 U16185 ( .ip1(n16168), .ip2(\ANSWER/mem[2][8][7] ), .s(n16745), .op(
        n3174) );
  mux2_1 U16186 ( .ip1(n16168), .ip2(\ANSWER/mem[2][9][7] ), .s(n16746), .op(
        n3173) );
  mux2_1 U16187 ( .ip1(n16168), .ip2(\ANSWER/mem[3][0][7] ), .s(n16747), .op(
        n3172) );
  mux2_1 U16188 ( .ip1(n16168), .ip2(\ANSWER/mem[3][1][7] ), .s(n16748), .op(
        n3171) );
  mux2_1 U16189 ( .ip1(n16168), .ip2(\ANSWER/mem[3][2][7] ), .s(n16749), .op(
        n3170) );
  mux2_1 U16190 ( .ip1(n16168), .ip2(\ANSWER/mem[3][3][7] ), .s(n16750), .op(
        n3169) );
  mux2_1 U16191 ( .ip1(n16168), .ip2(\ANSWER/mem[3][4][7] ), .s(n16751), .op(
        n3168) );
  mux2_1 U16192 ( .ip1(n16168), .ip2(\ANSWER/mem[3][5][7] ), .s(n16752), .op(
        n3167) );
  mux2_1 U16193 ( .ip1(n16170), .ip2(\ANSWER/mem[3][6][7] ), .s(n16753), .op(
        n3166) );
  mux2_1 U16194 ( .ip1(n16170), .ip2(\ANSWER/mem[3][7][7] ), .s(n16754), .op(
        n3165) );
  mux2_1 U16195 ( .ip1(n16170), .ip2(\ANSWER/mem[3][8][7] ), .s(n16755), .op(
        n3164) );
  mux2_1 U16196 ( .ip1(n16170), .ip2(\ANSWER/mem[3][9][7] ), .s(n16756), .op(
        n3163) );
  mux2_1 U16197 ( .ip1(n16169), .ip2(\ANSWER/mem[4][0][7] ), .s(n16757), .op(
        n3162) );
  mux2_1 U16198 ( .ip1(n16169), .ip2(\ANSWER/mem[4][1][7] ), .s(n16758), .op(
        n3161) );
  mux2_1 U16199 ( .ip1(n16169), .ip2(\ANSWER/mem[4][2][7] ), .s(n16759), .op(
        n3160) );
  mux2_1 U16200 ( .ip1(n16169), .ip2(\ANSWER/mem[4][3][7] ), .s(n16760), .op(
        n3159) );
  mux2_1 U16201 ( .ip1(n16170), .ip2(\ANSWER/mem[4][4][7] ), .s(n16761), .op(
        n3158) );
  mux2_1 U16202 ( .ip1(n16170), .ip2(\ANSWER/mem[4][5][7] ), .s(n16762), .op(
        n3157) );
  mux2_1 U16203 ( .ip1(n16170), .ip2(\ANSWER/mem[4][6][7] ), .s(n16763), .op(
        n3156) );
  mux2_1 U16204 ( .ip1(n16170), .ip2(\ANSWER/mem[4][7][7] ), .s(n16764), .op(
        n3155) );
  mux2_1 U16205 ( .ip1(n16170), .ip2(\ANSWER/mem[4][8][7] ), .s(n16765), .op(
        n3154) );
  mux2_1 U16206 ( .ip1(n16170), .ip2(\ANSWER/mem[4][9][7] ), .s(n16766), .op(
        n3153) );
  mux2_1 U16207 ( .ip1(n16170), .ip2(\ANSWER/mem[5][0][7] ), .s(n16767), .op(
        n3152) );
  mux2_1 U16208 ( .ip1(n16169), .ip2(\ANSWER/mem[5][1][7] ), .s(n16768), .op(
        n3151) );
  mux2_1 U16209 ( .ip1(n16170), .ip2(\ANSWER/mem[5][2][7] ), .s(n16769), .op(
        n3150) );
  mux2_1 U16210 ( .ip1(n16169), .ip2(\ANSWER/mem[5][3][7] ), .s(n16770), .op(
        n3149) );
  mux2_1 U16211 ( .ip1(n16170), .ip2(\ANSWER/mem[5][4][7] ), .s(n16771), .op(
        n3148) );
  mux2_1 U16212 ( .ip1(n16169), .ip2(\ANSWER/mem[5][5][7] ), .s(n16772), .op(
        n3147) );
  mux2_1 U16213 ( .ip1(n16169), .ip2(\ANSWER/mem[5][6][7] ), .s(n16773), .op(
        n3146) );
  mux2_1 U16214 ( .ip1(n16169), .ip2(\ANSWER/mem[5][7][7] ), .s(n16774), .op(
        n3145) );
  mux2_1 U16215 ( .ip1(n16169), .ip2(\ANSWER/mem[5][8][7] ), .s(n16775), .op(
        n3144) );
  mux2_1 U16216 ( .ip1(n16169), .ip2(\ANSWER/mem[5][9][7] ), .s(n16776), .op(
        n3143) );
  mux2_1 U16217 ( .ip1(n16169), .ip2(\ANSWER/mem[6][0][7] ), .s(n16777), .op(
        n3142) );
  mux2_1 U16218 ( .ip1(n16169), .ip2(\ANSWER/mem[6][1][7] ), .s(n16778), .op(
        n3141) );
  mux2_1 U16219 ( .ip1(n16169), .ip2(\ANSWER/mem[6][2][7] ), .s(n16779), .op(
        n3140) );
  mux2_1 U16220 ( .ip1(n16169), .ip2(\ANSWER/mem[6][3][7] ), .s(n16780), .op(
        n3139) );
  mux2_1 U16221 ( .ip1(n16169), .ip2(\ANSWER/mem[6][4][7] ), .s(n16781), .op(
        n3138) );
  mux2_1 U16222 ( .ip1(n16169), .ip2(\ANSWER/mem[6][5][7] ), .s(n16782), .op(
        n3137) );
  mux2_1 U16223 ( .ip1(n16169), .ip2(\ANSWER/mem[6][6][7] ), .s(n16783), .op(
        n3136) );
  mux2_1 U16224 ( .ip1(n16169), .ip2(\ANSWER/mem[6][7][7] ), .s(n16784), .op(
        n3135) );
  mux2_1 U16225 ( .ip1(n16169), .ip2(\ANSWER/mem[6][8][7] ), .s(n16785), .op(
        n3134) );
  mux2_1 U16226 ( .ip1(n16169), .ip2(\ANSWER/mem[6][9][7] ), .s(n16786), .op(
        n3133) );
  mux2_1 U16227 ( .ip1(n16169), .ip2(\ANSWER/mem[7][0][7] ), .s(n16787), .op(
        n3132) );
  mux2_1 U16228 ( .ip1(n16169), .ip2(\ANSWER/mem[7][1][7] ), .s(n16788), .op(
        n3131) );
  buf_1 U16229 ( .ip(n16169), .op(n16170) );
  mux2_1 U16230 ( .ip1(n16170), .ip2(\ANSWER/mem[7][2][7] ), .s(n16790), .op(
        n3130) );
  mux2_1 U16231 ( .ip1(n16170), .ip2(\ANSWER/mem[7][3][7] ), .s(n16791), .op(
        n3129) );
  mux2_1 U16232 ( .ip1(n16169), .ip2(\ANSWER/mem[7][4][7] ), .s(n16792), .op(
        n3128) );
  mux2_1 U16233 ( .ip1(n16169), .ip2(\ANSWER/mem[7][5][7] ), .s(n16793), .op(
        n3127) );
  mux2_1 U16234 ( .ip1(n16170), .ip2(\ANSWER/mem[7][6][7] ), .s(n16794), .op(
        n3126) );
  mux2_1 U16235 ( .ip1(n16170), .ip2(\ANSWER/mem[7][7][7] ), .s(n16795), .op(
        n3125) );
  mux2_1 U16236 ( .ip1(n16170), .ip2(\ANSWER/mem[7][8][7] ), .s(n16796), .op(
        n3124) );
  mux2_1 U16237 ( .ip1(n16170), .ip2(\ANSWER/mem[7][9][7] ), .s(n16797), .op(
        n3123) );
  mux2_1 U16238 ( .ip1(n16170), .ip2(\ANSWER/mem[8][0][7] ), .s(n16798), .op(
        n3122) );
  mux2_1 U16239 ( .ip1(n16170), .ip2(\ANSWER/mem[8][1][7] ), .s(n16799), .op(
        n3121) );
  mux2_1 U16240 ( .ip1(n16170), .ip2(\ANSWER/mem[8][2][7] ), .s(n16800), .op(
        n3120) );
  mux2_1 U16241 ( .ip1(n16170), .ip2(\ANSWER/mem[8][3][7] ), .s(n16801), .op(
        n3119) );
  mux2_1 U16242 ( .ip1(n16169), .ip2(\ANSWER/mem[8][4][7] ), .s(n16803), .op(
        n3118) );
  mux2_1 U16243 ( .ip1(n16169), .ip2(\ANSWER/mem[8][5][7] ), .s(n16804), .op(
        n3117) );
  mux2_1 U16244 ( .ip1(n16169), .ip2(\ANSWER/mem[8][6][7] ), .s(n16805), .op(
        n3116) );
  mux2_1 U16245 ( .ip1(n16169), .ip2(\ANSWER/mem[8][7][7] ), .s(n16806), .op(
        n3115) );
  mux2_1 U16246 ( .ip1(n16169), .ip2(\ANSWER/mem[8][8][7] ), .s(n16807), .op(
        n3114) );
  mux2_1 U16247 ( .ip1(n16169), .ip2(\ANSWER/mem[8][9][7] ), .s(n16808), .op(
        n3113) );
  mux2_1 U16248 ( .ip1(n16169), .ip2(\ANSWER/mem[9][0][7] ), .s(n16809), .op(
        n3112) );
  mux2_1 U16249 ( .ip1(n16169), .ip2(\ANSWER/mem[9][1][7] ), .s(n16810), .op(
        n3111) );
  mux2_1 U16250 ( .ip1(n16169), .ip2(\ANSWER/mem[9][2][7] ), .s(n16811), .op(
        n3110) );
  mux2_1 U16251 ( .ip1(n16169), .ip2(\ANSWER/mem[9][3][7] ), .s(n16812), .op(
        n3109) );
  mux2_1 U16252 ( .ip1(n16169), .ip2(\ANSWER/mem[9][4][7] ), .s(n16813), .op(
        n3108) );
  mux2_1 U16253 ( .ip1(n16169), .ip2(\ANSWER/mem[9][5][7] ), .s(n16814), .op(
        n3107) );
  mux2_1 U16254 ( .ip1(n16170), .ip2(\ANSWER/mem[9][6][7] ), .s(n16815), .op(
        n3106) );
  mux2_1 U16255 ( .ip1(n16170), .ip2(\ANSWER/mem[9][7][7] ), .s(n16816), .op(
        n3105) );
  mux2_1 U16256 ( .ip1(n16170), .ip2(\ANSWER/mem[9][8][7] ), .s(n16817), .op(
        n3104) );
  mux2_1 U16257 ( .ip1(n16170), .ip2(\ANSWER/mem[9][9][7] ), .s(n16818), .op(
        n3103) );
  fulladder U16258 ( .a(n16173), .b(n16172), .ci(n16171), .co(n16249), .s(
        n16160) );
  inv_1 U16259 ( .ip(n16249), .op(n16323) );
  and3_1 U16260 ( .ip1(m2DataIn[11]), .ip2(q_w2[6]), .ip3(n16185), .op(n16289)
         );
  nor2_1 U16261 ( .ip1(n16600), .ip2(n16538), .op(n16268) );
  or2_1 U16262 ( .ip1(q_w2[5]), .ip2(n16268), .op(n16175) );
  or2_1 U16263 ( .ip1(m2DataIn[11]), .ip2(n16268), .op(n16174) );
  nand2_1 U16264 ( .ip1(n16175), .ip2(n16174), .op(n16176) );
  nor2_1 U16265 ( .ip1(n16289), .ip2(n16176), .op(n16288) );
  nor2_1 U16266 ( .ip1(n16510), .ip2(n16177), .op(n16290) );
  xor2_1 U16267 ( .ip1(n16288), .ip2(n16290), .op(n16300) );
  and3_1 U16268 ( .ip1(m2DataIn[7]), .ip2(q_w2[10]), .ip3(n16178), .op(n16259)
         );
  nor2_1 U16269 ( .ip1(n16273), .ip2(n16622), .op(n16179) );
  or2_1 U16270 ( .ip1(q_w2[9]), .ip2(n16179), .op(n16181) );
  or2_1 U16271 ( .ip1(m2DataIn[7]), .ip2(n16179), .op(n16180) );
  nand2_1 U16272 ( .ip1(n16181), .ip2(n16180), .op(n16182) );
  nor2_1 U16273 ( .ip1(n16259), .ip2(n16182), .op(n16258) );
  nor2_1 U16274 ( .ip1(n16496), .ip2(n16599), .op(n16260) );
  xor2_1 U16275 ( .ip1(n16258), .ip2(n16260), .op(n16299) );
  fulladder U16276 ( .a(n16185), .b(n16184), .ci(n16183), .co(n16298), .s(
        n16202) );
  or2_1 U16277 ( .ip1(n16186), .ip2(n16187), .op(n16190) );
  or2_1 U16278 ( .ip1(n16188), .ip2(n16187), .op(n16189) );
  nand2_1 U16279 ( .ip1(n16190), .ip2(n16189), .op(n16304) );
  inv_1 U16280 ( .ip(rdata[8]), .op(n16295) );
  nor3_1 U16281 ( .ip1(n16690), .ip2(n16689), .ip3(n16191), .op(n16294) );
  nor2_1 U16282 ( .ip1(n16309), .ip2(n16689), .op(n16192) );
  or2_1 U16283 ( .ip1(q_w2[7]), .ip2(n16192), .op(n16194) );
  or2_1 U16284 ( .ip1(m2DataIn[9]), .ip2(n16192), .op(n16193) );
  nand2_1 U16285 ( .ip1(n16194), .ip2(n16193), .op(n16195) );
  nor2_1 U16286 ( .ip1(n16294), .ip2(n16195), .op(n16293) );
  mux2_1 U16287 ( .ip1(rdata[8]), .ip2(n16295), .s(n16293), .op(n16303) );
  fulladder U16288 ( .a(n16198), .b(n16197), .ci(n16196), .co(n16302), .s(
        n16146) );
  inv_1 U16289 ( .ip(n16199), .op(n16314) );
  fulladder U16290 ( .a(n16202), .b(n16201), .ci(n16200), .co(n16313), .s(
        n16147) );
  inv_1 U16291 ( .ip(n16203), .op(n16322) );
  nor2_1 U16292 ( .ip1(n16205), .ip2(n16204), .op(n16206) );
  nor2_1 U16293 ( .ip1(n16207), .ip2(n16206), .op(n16312) );
  nand2_1 U16294 ( .ip1(m2DataIn[12]), .ip2(q_w2[4]), .op(n16311) );
  or2_1 U16295 ( .ip1(rdata[7]), .ip2(n16208), .op(n16211) );
  or2_1 U16296 ( .ip1(n16209), .ip2(n16208), .op(n16210) );
  nand2_1 U16297 ( .ip1(n16211), .ip2(n16210), .op(n16310) );
  fulladder U16298 ( .a(n16214), .b(n16213), .ci(n16212), .co(n16318), .s(
        n16119) );
  fulladder U16299 ( .a(n16217), .b(n16216), .ci(n16215), .co(n16317), .s(
        n16103) );
  fulladder U16300 ( .a(n16220), .b(n16219), .ci(n16218), .co(n16320), .s(
        n16151) );
  inv_1 U16301 ( .ip(n16221), .op(n16257) );
  inv_1 U16302 ( .ip(q_w2[12]), .op(n16678) );
  nor2_1 U16303 ( .ip1(n16445), .ip2(n16678), .op(n16283) );
  nand2_1 U16304 ( .ip1(m2DataIn[15]), .ip2(q_w2[1]), .op(n16282) );
  nor2_1 U16305 ( .ip1(n16222), .ip2(n16495), .op(n16266) );
  nand2_1 U16306 ( .ip1(m2DataIn[3]), .ip2(q_w2[13]), .op(n16265) );
  nand2_1 U16307 ( .ip1(m2DataIn[14]), .ip2(q_w2[2]), .op(n16264) );
  inv_1 U16308 ( .ip(n16223), .op(n16285) );
  or2_1 U16309 ( .ip1(n16311), .ip2(n16224), .op(n16229) );
  inv_1 U16310 ( .ip(n16225), .op(n16227) );
  nand2_1 U16311 ( .ip1(n16227), .ip2(n16226), .op(n16228) );
  nand2_1 U16312 ( .ip1(n16229), .ip2(n16228), .op(n16284) );
  inv_1 U16313 ( .ip(n16230), .op(n16307) );
  fulladder U16314 ( .a(n16233), .b(n16232), .ci(n16231), .co(n16234), .s(
        n16241) );
  inv_1 U16315 ( .ip(n16234), .op(n16306) );
  fulladder U16316 ( .a(n16237), .b(n16236), .ci(n16235), .co(n16305), .s(
        n16133) );
  inv_1 U16317 ( .ip(n16238), .op(n16256) );
  fulladder U16318 ( .a(n16241), .b(n16240), .ci(n16239), .co(n16255), .s(
        n16173) );
  or2_1 U16319 ( .ip1(n16243), .ip2(n16242), .op(n16244) );
  nand2_1 U16320 ( .ip1(n16245), .ip2(n16244), .op(n16246) );
  or2_1 U16321 ( .ip1(n16247), .ip2(n16246), .op(n16326) );
  nand2_1 U16322 ( .ip1(n16247), .ip2(n16246), .op(n16324) );
  nand2_1 U16323 ( .ip1(n16326), .ip2(n16324), .op(n16248) );
  mux2_1 U16324 ( .ip1(n16323), .ip2(n16249), .s(n16248), .op(n16251) );
  nor3_1 U16325 ( .ip1(\SIGMOID/lut_out [7]), .ip2(\SIGMOID/sign_bit ), .ip3(
        n16250), .op(n16827) );
  mux2_1 U16326 ( .ip1(n16251), .ip2(n16827), .s(n16714), .op(n16252) );
  buf_1 U16327 ( .ip(n16252), .op(n16253) );
  mux2_1 U16328 ( .ip1(n16253), .ip2(\ANSWER/mem[0][0][8] ), .s(n16717), .op(
        n3102) );
  mux2_1 U16329 ( .ip1(n16253), .ip2(\ANSWER/mem[0][1][8] ), .s(n16718), .op(
        n3101) );
  mux2_1 U16330 ( .ip1(n16253), .ip2(\ANSWER/mem[0][2][8] ), .s(n16719), .op(
        n3100) );
  mux2_1 U16331 ( .ip1(n16252), .ip2(\ANSWER/mem[0][3][8] ), .s(n16720), .op(
        n3099) );
  mux2_1 U16332 ( .ip1(n16253), .ip2(\ANSWER/mem[0][4][8] ), .s(n16721), .op(
        n3098) );
  buf_1 U16333 ( .ip(n16252), .op(n16254) );
  mux2_1 U16334 ( .ip1(n16254), .ip2(\ANSWER/mem[0][5][8] ), .s(n16722), .op(
        n3097) );
  mux2_1 U16335 ( .ip1(n16254), .ip2(\ANSWER/mem[0][6][8] ), .s(n16723), .op(
        n3096) );
  mux2_1 U16336 ( .ip1(n16253), .ip2(\ANSWER/mem[0][7][8] ), .s(n16724), .op(
        n3095) );
  mux2_1 U16337 ( .ip1(n16252), .ip2(\ANSWER/mem[0][8][8] ), .s(n16725), .op(
        n3094) );
  mux2_1 U16338 ( .ip1(n16253), .ip2(\ANSWER/mem[0][9][8] ), .s(n16726), .op(
        n3093) );
  mux2_1 U16339 ( .ip1(n16252), .ip2(\ANSWER/mem[1][0][8] ), .s(n16727), .op(
        n3092) );
  mux2_1 U16340 ( .ip1(n16254), .ip2(\ANSWER/mem[1][1][8] ), .s(n16728), .op(
        n3091) );
  mux2_1 U16341 ( .ip1(n16253), .ip2(\ANSWER/mem[1][2][8] ), .s(n16729), .op(
        n3090) );
  mux2_1 U16342 ( .ip1(n16254), .ip2(\ANSWER/mem[1][3][8] ), .s(n16730), .op(
        n3089) );
  mux2_1 U16343 ( .ip1(n16253), .ip2(\ANSWER/mem[1][4][8] ), .s(n16731), .op(
        n3088) );
  mux2_1 U16344 ( .ip1(n16254), .ip2(\ANSWER/mem[1][5][8] ), .s(n16732), .op(
        n3087) );
  mux2_1 U16345 ( .ip1(n16253), .ip2(\ANSWER/mem[1][6][8] ), .s(n16733), .op(
        n3086) );
  mux2_1 U16346 ( .ip1(n16254), .ip2(\ANSWER/mem[1][7][8] ), .s(n16734), .op(
        n3085) );
  mux2_1 U16347 ( .ip1(n16253), .ip2(\ANSWER/mem[1][8][8] ), .s(n16735), .op(
        n3084) );
  mux2_1 U16348 ( .ip1(n16254), .ip2(\ANSWER/mem[1][9][8] ), .s(n16736), .op(
        n3083) );
  mux2_1 U16349 ( .ip1(n16253), .ip2(\ANSWER/mem[2][0][8] ), .s(n16737), .op(
        n3082) );
  mux2_1 U16350 ( .ip1(n16254), .ip2(\ANSWER/mem[2][1][8] ), .s(n16738), .op(
        n3081) );
  mux2_1 U16351 ( .ip1(n16253), .ip2(\ANSWER/mem[2][2][8] ), .s(n16739), .op(
        n3080) );
  mux2_1 U16352 ( .ip1(n16254), .ip2(\ANSWER/mem[2][3][8] ), .s(n16740), .op(
        n3079) );
  mux2_1 U16353 ( .ip1(n16252), .ip2(\ANSWER/mem[2][4][8] ), .s(n16741), .op(
        n3078) );
  mux2_1 U16354 ( .ip1(n16252), .ip2(\ANSWER/mem[2][5][8] ), .s(n16742), .op(
        n3077) );
  mux2_1 U16355 ( .ip1(n16252), .ip2(\ANSWER/mem[2][6][8] ), .s(n16743), .op(
        n3076) );
  mux2_1 U16356 ( .ip1(n16252), .ip2(\ANSWER/mem[2][7][8] ), .s(n16744), .op(
        n3075) );
  mux2_1 U16357 ( .ip1(n16252), .ip2(\ANSWER/mem[2][8][8] ), .s(n16745), .op(
        n3074) );
  mux2_1 U16358 ( .ip1(n16252), .ip2(\ANSWER/mem[2][9][8] ), .s(n16746), .op(
        n3073) );
  mux2_1 U16359 ( .ip1(n16252), .ip2(\ANSWER/mem[3][0][8] ), .s(n16747), .op(
        n3072) );
  mux2_1 U16360 ( .ip1(n16252), .ip2(\ANSWER/mem[3][1][8] ), .s(n16748), .op(
        n3071) );
  mux2_1 U16361 ( .ip1(n16252), .ip2(\ANSWER/mem[3][2][8] ), .s(n16749), .op(
        n3070) );
  mux2_1 U16362 ( .ip1(n16253), .ip2(\ANSWER/mem[3][3][8] ), .s(n16750), .op(
        n3069) );
  mux2_1 U16363 ( .ip1(n16254), .ip2(\ANSWER/mem[3][4][8] ), .s(n16751), .op(
        n3068) );
  mux2_1 U16364 ( .ip1(n16254), .ip2(\ANSWER/mem[3][5][8] ), .s(n16752), .op(
        n3067) );
  mux2_1 U16365 ( .ip1(n16252), .ip2(\ANSWER/mem[3][6][8] ), .s(n16753), .op(
        n3066) );
  mux2_1 U16366 ( .ip1(n16252), .ip2(\ANSWER/mem[3][7][8] ), .s(n16754), .op(
        n3065) );
  mux2_1 U16367 ( .ip1(n16252), .ip2(\ANSWER/mem[3][8][8] ), .s(n16755), .op(
        n3064) );
  mux2_1 U16368 ( .ip1(n16252), .ip2(\ANSWER/mem[3][9][8] ), .s(n16756), .op(
        n3063) );
  mux2_1 U16369 ( .ip1(n16252), .ip2(\ANSWER/mem[4][0][8] ), .s(n16757), .op(
        n3062) );
  mux2_1 U16370 ( .ip1(n16252), .ip2(\ANSWER/mem[4][1][8] ), .s(n16758), .op(
        n3061) );
  mux2_1 U16371 ( .ip1(n16252), .ip2(\ANSWER/mem[4][2][8] ), .s(n16759), .op(
        n3060) );
  mux2_1 U16372 ( .ip1(n16252), .ip2(\ANSWER/mem[4][3][8] ), .s(n16760), .op(
        n3059) );
  mux2_1 U16373 ( .ip1(n16252), .ip2(\ANSWER/mem[4][4][8] ), .s(n16761), .op(
        n3058) );
  mux2_1 U16374 ( .ip1(n16252), .ip2(\ANSWER/mem[4][5][8] ), .s(n16762), .op(
        n3057) );
  mux2_1 U16375 ( .ip1(n16252), .ip2(\ANSWER/mem[4][6][8] ), .s(n16763), .op(
        n3056) );
  mux2_1 U16376 ( .ip1(n16252), .ip2(\ANSWER/mem[4][7][8] ), .s(n16764), .op(
        n3055) );
  mux2_1 U16377 ( .ip1(n16254), .ip2(\ANSWER/mem[4][8][8] ), .s(n16765), .op(
        n3054) );
  mux2_1 U16378 ( .ip1(n16253), .ip2(\ANSWER/mem[4][9][8] ), .s(n16766), .op(
        n3053) );
  mux2_1 U16379 ( .ip1(n16254), .ip2(\ANSWER/mem[5][0][8] ), .s(n16767), .op(
        n3052) );
  mux2_1 U16380 ( .ip1(n16252), .ip2(\ANSWER/mem[5][1][8] ), .s(n16768), .op(
        n3051) );
  mux2_1 U16381 ( .ip1(n16253), .ip2(\ANSWER/mem[5][2][8] ), .s(n16769), .op(
        n3050) );
  mux2_1 U16382 ( .ip1(n16253), .ip2(\ANSWER/mem[5][3][8] ), .s(n16770), .op(
        n3049) );
  mux2_1 U16383 ( .ip1(n16252), .ip2(\ANSWER/mem[5][4][8] ), .s(n16771), .op(
        n3048) );
  mux2_1 U16384 ( .ip1(n16252), .ip2(\ANSWER/mem[5][5][8] ), .s(n16772), .op(
        n3047) );
  mux2_1 U16385 ( .ip1(n16252), .ip2(\ANSWER/mem[5][6][8] ), .s(n16773), .op(
        n3046) );
  mux2_1 U16386 ( .ip1(n16252), .ip2(\ANSWER/mem[5][7][8] ), .s(n16774), .op(
        n3045) );
  mux2_1 U16387 ( .ip1(n16252), .ip2(\ANSWER/mem[5][8][8] ), .s(n16775), .op(
        n3044) );
  mux2_1 U16388 ( .ip1(n16252), .ip2(\ANSWER/mem[5][9][8] ), .s(n16776), .op(
        n3043) );
  mux2_1 U16389 ( .ip1(n16254), .ip2(\ANSWER/mem[6][0][8] ), .s(n16777), .op(
        n3042) );
  mux2_1 U16390 ( .ip1(n16254), .ip2(\ANSWER/mem[6][1][8] ), .s(n16778), .op(
        n3041) );
  mux2_1 U16391 ( .ip1(n16254), .ip2(\ANSWER/mem[6][2][8] ), .s(n16779), .op(
        n3040) );
  mux2_1 U16392 ( .ip1(n16254), .ip2(\ANSWER/mem[6][3][8] ), .s(n16780), .op(
        n3039) );
  mux2_1 U16393 ( .ip1(n16254), .ip2(\ANSWER/mem[6][4][8] ), .s(n16781), .op(
        n3038) );
  mux2_1 U16394 ( .ip1(n16254), .ip2(\ANSWER/mem[6][5][8] ), .s(n16782), .op(
        n3037) );
  mux2_1 U16395 ( .ip1(n16254), .ip2(\ANSWER/mem[6][6][8] ), .s(n16783), .op(
        n3036) );
  mux2_1 U16396 ( .ip1(n16253), .ip2(\ANSWER/mem[6][7][8] ), .s(n16784), .op(
        n3035) );
  mux2_1 U16397 ( .ip1(n16254), .ip2(\ANSWER/mem[6][8][8] ), .s(n16785), .op(
        n3034) );
  mux2_1 U16398 ( .ip1(n16252), .ip2(\ANSWER/mem[6][9][8] ), .s(n16786), .op(
        n3033) );
  mux2_1 U16399 ( .ip1(n16252), .ip2(\ANSWER/mem[7][0][8] ), .s(n16787), .op(
        n3032) );
  mux2_1 U16400 ( .ip1(n16254), .ip2(\ANSWER/mem[7][1][8] ), .s(n16788), .op(
        n3031) );
  mux2_1 U16401 ( .ip1(n16254), .ip2(\ANSWER/mem[7][2][8] ), .s(n16790), .op(
        n3030) );
  mux2_1 U16402 ( .ip1(n16252), .ip2(\ANSWER/mem[7][3][8] ), .s(n16791), .op(
        n3029) );
  mux2_1 U16403 ( .ip1(n16253), .ip2(\ANSWER/mem[7][4][8] ), .s(n16792), .op(
        n3028) );
  mux2_1 U16404 ( .ip1(n16253), .ip2(\ANSWER/mem[7][5][8] ), .s(n16793), .op(
        n3027) );
  mux2_1 U16405 ( .ip1(n16252), .ip2(\ANSWER/mem[7][6][8] ), .s(n16794), .op(
        n3026) );
  mux2_1 U16406 ( .ip1(n16252), .ip2(\ANSWER/mem[7][7][8] ), .s(n16795), .op(
        n3025) );
  mux2_1 U16407 ( .ip1(n16254), .ip2(\ANSWER/mem[7][8][8] ), .s(n16796), .op(
        n3024) );
  mux2_1 U16408 ( .ip1(n16252), .ip2(\ANSWER/mem[7][9][8] ), .s(n16797), .op(
        n3023) );
  mux2_1 U16409 ( .ip1(n16254), .ip2(\ANSWER/mem[8][0][8] ), .s(n16798), .op(
        n3022) );
  mux2_1 U16410 ( .ip1(n16254), .ip2(\ANSWER/mem[8][1][8] ), .s(n16799), .op(
        n3021) );
  mux2_1 U16411 ( .ip1(n16252), .ip2(\ANSWER/mem[8][2][8] ), .s(n16800), .op(
        n3020) );
  mux2_1 U16412 ( .ip1(n16254), .ip2(\ANSWER/mem[8][3][8] ), .s(n16801), .op(
        n3019) );
  mux2_1 U16413 ( .ip1(n16253), .ip2(\ANSWER/mem[8][4][8] ), .s(n16803), .op(
        n3018) );
  mux2_1 U16414 ( .ip1(n16253), .ip2(\ANSWER/mem[8][5][8] ), .s(n16804), .op(
        n3017) );
  mux2_1 U16415 ( .ip1(n16253), .ip2(\ANSWER/mem[8][6][8] ), .s(n16805), .op(
        n3016) );
  mux2_1 U16416 ( .ip1(n16253), .ip2(\ANSWER/mem[8][7][8] ), .s(n16806), .op(
        n3015) );
  mux2_1 U16417 ( .ip1(n16253), .ip2(\ANSWER/mem[8][8][8] ), .s(n16807), .op(
        n3014) );
  mux2_1 U16418 ( .ip1(n16253), .ip2(\ANSWER/mem[8][9][8] ), .s(n16808), .op(
        n3013) );
  mux2_1 U16419 ( .ip1(n16253), .ip2(\ANSWER/mem[9][0][8] ), .s(n16809), .op(
        n3012) );
  mux2_1 U16420 ( .ip1(n16253), .ip2(\ANSWER/mem[9][1][8] ), .s(n16810), .op(
        n3011) );
  mux2_1 U16421 ( .ip1(n16253), .ip2(\ANSWER/mem[9][2][8] ), .s(n16811), .op(
        n3010) );
  mux2_1 U16422 ( .ip1(n16253), .ip2(\ANSWER/mem[9][3][8] ), .s(n16812), .op(
        n3009) );
  mux2_1 U16423 ( .ip1(n16253), .ip2(\ANSWER/mem[9][4][8] ), .s(n16813), .op(
        n3008) );
  mux2_1 U16424 ( .ip1(n16253), .ip2(\ANSWER/mem[9][5][8] ), .s(n16814), .op(
        n3007) );
  mux2_1 U16425 ( .ip1(n16254), .ip2(\ANSWER/mem[9][6][8] ), .s(n16815), .op(
        n3006) );
  mux2_1 U16426 ( .ip1(n16254), .ip2(\ANSWER/mem[9][7][8] ), .s(n16816), .op(
        n3005) );
  mux2_1 U16427 ( .ip1(n16254), .ip2(\ANSWER/mem[9][8][8] ), .s(n16817), .op(
        n3004) );
  mux2_1 U16428 ( .ip1(n16254), .ip2(\ANSWER/mem[9][9][8] ), .s(n16818), .op(
        n3003) );
  fulladder U16429 ( .a(n16257), .b(n16256), .ci(n16255), .co(n16389), .s(
        n16247) );
  or2_1 U16430 ( .ip1(n16258), .ip2(n16259), .op(n16262) );
  or2_1 U16431 ( .ip1(n16260), .ip2(n16259), .op(n16261) );
  nand2_1 U16432 ( .ip1(n16262), .ip2(n16261), .op(n16382) );
  nor2_1 U16433 ( .ip1(n16690), .ip2(n16596), .op(n16372) );
  inv_1 U16434 ( .ip(n16263), .op(n16381) );
  fulladder U16435 ( .a(n16266), .b(n16265), .ci(n16264), .co(n16380), .s(
        n16223) );
  inv_1 U16436 ( .ip(n16267), .op(n16340) );
  and3_1 U16437 ( .ip1(m2DataIn[11]), .ip2(q_w2[7]), .ip3(n16268), .op(n16343)
         );
  nor2_1 U16438 ( .ip1(n16679), .ip2(n16538), .op(n16269) );
  or2_1 U16439 ( .ip1(q_w2[7]), .ip2(n16269), .op(n16271) );
  or2_1 U16440 ( .ip1(m2DataIn[10]), .ip2(n16269), .op(n16270) );
  nand2_1 U16441 ( .ip1(n16271), .ip2(n16270), .op(n16272) );
  nor2_1 U16442 ( .ip1(n16343), .ip2(n16272), .op(n16342) );
  nor2_1 U16443 ( .ip1(n16510), .ip2(n16447), .op(n16344) );
  xor2_1 U16444 ( .ip1(n16342), .ip2(n16344), .op(n16378) );
  nand2_1 U16445 ( .ip1(m2DataIn[7]), .ip2(q_w2[11]), .op(n16432) );
  nor3_1 U16446 ( .ip1(n16273), .ip2(n16622), .ip3(n16432), .op(n16355) );
  inv_1 U16447 ( .ip(n16355), .op(n16277) );
  nand2_1 U16448 ( .ip1(m2DataIn[6]), .ip2(q_w2[11]), .op(n16275) );
  nand2_1 U16449 ( .ip1(m2DataIn[7]), .ip2(q_w2[10]), .op(n16274) );
  nand2_1 U16450 ( .ip1(n16275), .ip2(n16274), .op(n16276) );
  nand2_1 U16451 ( .ip1(n16277), .ip2(n16276), .op(n16278) );
  nor3_1 U16452 ( .ip1(n16496), .ip2(n16678), .ip3(n16278), .op(n16354) );
  or2_1 U16453 ( .ip1(n16278), .ip2(n16354), .op(n16281) );
  nand2_1 U16454 ( .ip1(m2DataIn[5]), .ip2(q_w2[12]), .op(n16279) );
  or2_1 U16455 ( .ip1(n16279), .ip2(n16354), .op(n16280) );
  nand2_1 U16456 ( .ip1(n16281), .ip2(n16280), .op(n16377) );
  fulladder U16457 ( .a(n16413), .b(n16283), .ci(n16282), .co(n16376), .s(
        n16286) );
  fulladder U16458 ( .a(n16286), .b(n16285), .ci(n16284), .co(n16338), .s(
        n16230) );
  inv_1 U16459 ( .ip(n16287), .op(n16388) );
  nand2_1 U16460 ( .ip1(m2DataIn[12]), .ip2(q_w2[5]), .op(n16418) );
  or2_1 U16461 ( .ip1(n16288), .ip2(n16289), .op(n16292) );
  or2_1 U16462 ( .ip1(n16290), .ip2(n16289), .op(n16291) );
  nand2_1 U16463 ( .ip1(n16292), .ip2(n16291), .op(n16371) );
  or2_1 U16464 ( .ip1(n16293), .ip2(n16294), .op(n16297) );
  or2_1 U16465 ( .ip1(n16295), .ip2(n16294), .op(n16296) );
  nand2_1 U16466 ( .ip1(n16297), .ip2(n16296), .op(n16370) );
  fulladder U16467 ( .a(n16300), .b(n16299), .ci(n16298), .co(n16301), .s(
        n16315) );
  inv_1 U16468 ( .ip(n16301), .op(n16384) );
  fulladder U16469 ( .a(n16304), .b(n16303), .ci(n16302), .co(n16383), .s(
        n16199) );
  fulladder U16470 ( .a(n16307), .b(n16306), .ci(n16305), .co(n16386), .s(
        n16238) );
  inv_1 U16471 ( .ip(m2DataIn[15]), .op(n16498) );
  nor2_1 U16472 ( .ip1(n16498), .ip2(n16308), .op(n16361) );
  nand2_1 U16473 ( .ip1(m2DataIn[4]), .ip2(q_w2[13]), .op(n16360) );
  nand2_1 U16474 ( .ip1(m2DataIn[8]), .ip2(q_w2[9]), .op(n16359) );
  nor2_1 U16475 ( .ip1(n16309), .ip2(n16495), .op(n16353) );
  nand2_1 U16476 ( .ip1(m2DataIn[14]), .ip2(q_w2[3]), .op(n16351) );
  fulladder U16477 ( .a(n16312), .b(n16311), .ci(n16310), .co(n16362), .s(
        n16319) );
  fulladder U16478 ( .a(n16315), .b(n16314), .ci(n16313), .co(n16316), .s(
        n16203) );
  inv_1 U16479 ( .ip(n16316), .op(n16366) );
  fulladder U16480 ( .a(n16319), .b(n16318), .ci(n16317), .co(n16365), .s(
        n16321) );
  fulladder U16481 ( .a(n16322), .b(n16321), .ci(n16320), .co(n16335), .s(
        n16221) );
  nand2_1 U16482 ( .ip1(n16324), .ip2(n16323), .op(n16325) );
  nand2_1 U16483 ( .ip1(n16326), .ip2(n16325), .op(n16327) );
  nand2_1 U16484 ( .ip1(n16328), .ip2(n16327), .op(n16392) );
  inv_1 U16485 ( .ip(n16392), .op(n16329) );
  nor2_1 U16486 ( .ip1(n16328), .ip2(n16327), .op(n16390) );
  nor2_1 U16487 ( .ip1(n16329), .ip2(n16390), .op(n16331) );
  nor2_1 U16488 ( .ip1(n16389), .ip2(n16331), .op(n16330) );
  not_ab_or_c_or_d U16489 ( .ip1(n16389), .ip2(n16331), .ip3(n16714), .ip4(
        n16330), .op(n16332) );
  buf_1 U16490 ( .ip(n16332), .op(n16334) );
  mux2_1 U16491 ( .ip1(n16334), .ip2(\ANSWER/mem[0][0][9] ), .s(n16717), .op(
        n3002) );
  mux2_1 U16492 ( .ip1(n16334), .ip2(\ANSWER/mem[0][1][9] ), .s(n16718), .op(
        n3001) );
  mux2_1 U16493 ( .ip1(n16334), .ip2(\ANSWER/mem[0][2][9] ), .s(n16719), .op(
        n3000) );
  mux2_1 U16494 ( .ip1(n16334), .ip2(\ANSWER/mem[0][3][9] ), .s(n16720), .op(
        n2999) );
  mux2_1 U16495 ( .ip1(n16334), .ip2(\ANSWER/mem[0][4][9] ), .s(n16721), .op(
        n2998) );
  mux2_1 U16496 ( .ip1(n16334), .ip2(\ANSWER/mem[0][5][9] ), .s(n16722), .op(
        n2997) );
  mux2_1 U16497 ( .ip1(n16334), .ip2(\ANSWER/mem[0][6][9] ), .s(n16723), .op(
        n2996) );
  mux2_1 U16498 ( .ip1(n16334), .ip2(\ANSWER/mem[0][7][9] ), .s(n16724), .op(
        n2995) );
  mux2_1 U16499 ( .ip1(n16334), .ip2(\ANSWER/mem[0][8][9] ), .s(n16725), .op(
        n2994) );
  mux2_1 U16500 ( .ip1(n16334), .ip2(\ANSWER/mem[0][9][9] ), .s(n16726), .op(
        n2993) );
  mux2_1 U16501 ( .ip1(n16334), .ip2(\ANSWER/mem[1][0][9] ), .s(n16727), .op(
        n2992) );
  mux2_1 U16502 ( .ip1(n16334), .ip2(\ANSWER/mem[1][1][9] ), .s(n16728), .op(
        n2991) );
  mux2_1 U16503 ( .ip1(n16334), .ip2(\ANSWER/mem[1][2][9] ), .s(n16729), .op(
        n2990) );
  mux2_1 U16504 ( .ip1(n16332), .ip2(\ANSWER/mem[1][3][9] ), .s(n16730), .op(
        n2989) );
  mux2_1 U16505 ( .ip1(n16332), .ip2(\ANSWER/mem[1][4][9] ), .s(n16731), .op(
        n2988) );
  mux2_1 U16506 ( .ip1(n16332), .ip2(\ANSWER/mem[1][5][9] ), .s(n16732), .op(
        n2987) );
  mux2_1 U16507 ( .ip1(n16332), .ip2(\ANSWER/mem[1][6][9] ), .s(n16733), .op(
        n2986) );
  mux2_1 U16508 ( .ip1(n16332), .ip2(\ANSWER/mem[1][7][9] ), .s(n16734), .op(
        n2985) );
  mux2_1 U16509 ( .ip1(n16332), .ip2(\ANSWER/mem[1][8][9] ), .s(n16735), .op(
        n2984) );
  mux2_1 U16510 ( .ip1(n16332), .ip2(\ANSWER/mem[1][9][9] ), .s(n16736), .op(
        n2983) );
  mux2_1 U16511 ( .ip1(n16332), .ip2(\ANSWER/mem[2][0][9] ), .s(n16737), .op(
        n2982) );
  mux2_1 U16512 ( .ip1(n16332), .ip2(\ANSWER/mem[2][1][9] ), .s(n16738), .op(
        n2981) );
  mux2_1 U16513 ( .ip1(n16332), .ip2(\ANSWER/mem[2][2][9] ), .s(n16739), .op(
        n2980) );
  mux2_1 U16514 ( .ip1(n16332), .ip2(\ANSWER/mem[2][3][9] ), .s(n16740), .op(
        n2979) );
  mux2_1 U16515 ( .ip1(n16334), .ip2(\ANSWER/mem[2][4][9] ), .s(n16741), .op(
        n2978) );
  mux2_1 U16516 ( .ip1(n16332), .ip2(\ANSWER/mem[2][5][9] ), .s(n16742), .op(
        n2977) );
  mux2_1 U16517 ( .ip1(n16334), .ip2(\ANSWER/mem[2][6][9] ), .s(n16743), .op(
        n2976) );
  mux2_1 U16518 ( .ip1(n16332), .ip2(\ANSWER/mem[2][7][9] ), .s(n16744), .op(
        n2975) );
  mux2_1 U16519 ( .ip1(n16332), .ip2(\ANSWER/mem[2][8][9] ), .s(n16745), .op(
        n2974) );
  mux2_1 U16520 ( .ip1(n16332), .ip2(\ANSWER/mem[2][9][9] ), .s(n16746), .op(
        n2973) );
  mux2_1 U16521 ( .ip1(n16334), .ip2(\ANSWER/mem[3][0][9] ), .s(n16747), .op(
        n2972) );
  mux2_1 U16522 ( .ip1(n16334), .ip2(\ANSWER/mem[3][1][9] ), .s(n16748), .op(
        n2971) );
  mux2_1 U16523 ( .ip1(n16334), .ip2(\ANSWER/mem[3][2][9] ), .s(n16749), .op(
        n2970) );
  mux2_1 U16524 ( .ip1(n16334), .ip2(\ANSWER/mem[3][3][9] ), .s(n16750), .op(
        n2969) );
  mux2_1 U16525 ( .ip1(n16334), .ip2(\ANSWER/mem[3][4][9] ), .s(n16751), .op(
        n2968) );
  mux2_1 U16526 ( .ip1(n16334), .ip2(\ANSWER/mem[3][5][9] ), .s(n16752), .op(
        n2967) );
  buf_1 U16527 ( .ip(n16332), .op(n16333) );
  mux2_1 U16528 ( .ip1(n16333), .ip2(\ANSWER/mem[3][6][9] ), .s(n16753), .op(
        n2966) );
  mux2_1 U16529 ( .ip1(n16332), .ip2(\ANSWER/mem[3][7][9] ), .s(n16754), .op(
        n2965) );
  mux2_1 U16530 ( .ip1(n16332), .ip2(\ANSWER/mem[3][8][9] ), .s(n16755), .op(
        n2964) );
  mux2_1 U16531 ( .ip1(n16332), .ip2(\ANSWER/mem[3][9][9] ), .s(n16756), .op(
        n2963) );
  mux2_1 U16532 ( .ip1(n16333), .ip2(\ANSWER/mem[4][0][9] ), .s(n16757), .op(
        n2962) );
  mux2_1 U16533 ( .ip1(n16333), .ip2(\ANSWER/mem[4][1][9] ), .s(n16758), .op(
        n2961) );
  mux2_1 U16534 ( .ip1(n16333), .ip2(\ANSWER/mem[4][2][9] ), .s(n16759), .op(
        n2960) );
  mux2_1 U16535 ( .ip1(n16333), .ip2(\ANSWER/mem[4][3][9] ), .s(n16760), .op(
        n2959) );
  mux2_1 U16536 ( .ip1(n16333), .ip2(\ANSWER/mem[4][4][9] ), .s(n16761), .op(
        n2958) );
  mux2_1 U16537 ( .ip1(n16333), .ip2(\ANSWER/mem[4][5][9] ), .s(n16762), .op(
        n2957) );
  mux2_1 U16538 ( .ip1(n16333), .ip2(\ANSWER/mem[4][6][9] ), .s(n16763), .op(
        n2956) );
  mux2_1 U16539 ( .ip1(n16333), .ip2(\ANSWER/mem[4][7][9] ), .s(n16764), .op(
        n2955) );
  mux2_1 U16540 ( .ip1(n16334), .ip2(\ANSWER/mem[4][8][9] ), .s(n16765), .op(
        n2954) );
  mux2_1 U16541 ( .ip1(n16332), .ip2(\ANSWER/mem[4][9][9] ), .s(n16766), .op(
        n2953) );
  mux2_1 U16542 ( .ip1(n16332), .ip2(\ANSWER/mem[5][0][9] ), .s(n16767), .op(
        n2952) );
  mux2_1 U16543 ( .ip1(n16332), .ip2(\ANSWER/mem[5][1][9] ), .s(n16768), .op(
        n2951) );
  mux2_1 U16544 ( .ip1(n16332), .ip2(\ANSWER/mem[5][2][9] ), .s(n16769), .op(
        n2950) );
  mux2_1 U16545 ( .ip1(n16332), .ip2(\ANSWER/mem[5][3][9] ), .s(n16770), .op(
        n2949) );
  mux2_1 U16546 ( .ip1(n16332), .ip2(\ANSWER/mem[5][4][9] ), .s(n16771), .op(
        n2948) );
  mux2_1 U16547 ( .ip1(n16332), .ip2(\ANSWER/mem[5][5][9] ), .s(n16772), .op(
        n2947) );
  mux2_1 U16548 ( .ip1(n16332), .ip2(\ANSWER/mem[5][6][9] ), .s(n16773), .op(
        n2946) );
  mux2_1 U16549 ( .ip1(n16332), .ip2(\ANSWER/mem[5][7][9] ), .s(n16774), .op(
        n2945) );
  mux2_1 U16550 ( .ip1(n16332), .ip2(\ANSWER/mem[5][8][9] ), .s(n16775), .op(
        n2944) );
  mux2_1 U16551 ( .ip1(n16332), .ip2(\ANSWER/mem[5][9][9] ), .s(n16776), .op(
        n2943) );
  mux2_1 U16552 ( .ip1(n16333), .ip2(\ANSWER/mem[6][0][9] ), .s(n16777), .op(
        n2942) );
  mux2_1 U16553 ( .ip1(n16333), .ip2(\ANSWER/mem[6][1][9] ), .s(n16778), .op(
        n2941) );
  mux2_1 U16554 ( .ip1(n16333), .ip2(\ANSWER/mem[6][2][9] ), .s(n16779), .op(
        n2940) );
  mux2_1 U16555 ( .ip1(n16333), .ip2(\ANSWER/mem[6][3][9] ), .s(n16780), .op(
        n2939) );
  mux2_1 U16556 ( .ip1(n16332), .ip2(\ANSWER/mem[6][4][9] ), .s(n16781), .op(
        n2938) );
  mux2_1 U16557 ( .ip1(n16332), .ip2(\ANSWER/mem[6][5][9] ), .s(n16782), .op(
        n2937) );
  mux2_1 U16558 ( .ip1(n16332), .ip2(\ANSWER/mem[6][6][9] ), .s(n16783), .op(
        n2936) );
  mux2_1 U16559 ( .ip1(n16332), .ip2(\ANSWER/mem[6][7][9] ), .s(n16784), .op(
        n2935) );
  mux2_1 U16560 ( .ip1(n16332), .ip2(\ANSWER/mem[6][8][9] ), .s(n16785), .op(
        n2934) );
  mux2_1 U16561 ( .ip1(n16332), .ip2(\ANSWER/mem[6][9][9] ), .s(n16786), .op(
        n2933) );
  mux2_1 U16562 ( .ip1(n16332), .ip2(\ANSWER/mem[7][0][9] ), .s(n16787), .op(
        n2932) );
  mux2_1 U16563 ( .ip1(n16332), .ip2(\ANSWER/mem[7][1][9] ), .s(n16788), .op(
        n2931) );
  mux2_1 U16564 ( .ip1(n16333), .ip2(\ANSWER/mem[7][2][9] ), .s(n16790), .op(
        n2930) );
  mux2_1 U16565 ( .ip1(n16333), .ip2(\ANSWER/mem[7][3][9] ), .s(n16791), .op(
        n2929) );
  mux2_1 U16566 ( .ip1(n16333), .ip2(\ANSWER/mem[7][4][9] ), .s(n16792), .op(
        n2928) );
  mux2_1 U16567 ( .ip1(n16333), .ip2(\ANSWER/mem[7][5][9] ), .s(n16793), .op(
        n2927) );
  mux2_1 U16568 ( .ip1(n16333), .ip2(\ANSWER/mem[7][6][9] ), .s(n16794), .op(
        n2926) );
  mux2_1 U16569 ( .ip1(n16333), .ip2(\ANSWER/mem[7][7][9] ), .s(n16795), .op(
        n2925) );
  mux2_1 U16570 ( .ip1(n16333), .ip2(\ANSWER/mem[7][8][9] ), .s(n16796), .op(
        n2924) );
  mux2_1 U16571 ( .ip1(n16333), .ip2(\ANSWER/mem[7][9][9] ), .s(n16797), .op(
        n2923) );
  mux2_1 U16572 ( .ip1(n16333), .ip2(\ANSWER/mem[8][0][9] ), .s(n16798), .op(
        n2922) );
  mux2_1 U16573 ( .ip1(n16333), .ip2(\ANSWER/mem[8][1][9] ), .s(n16799), .op(
        n2921) );
  mux2_1 U16574 ( .ip1(n16333), .ip2(\ANSWER/mem[8][2][9] ), .s(n16800), .op(
        n2920) );
  mux2_1 U16575 ( .ip1(n16333), .ip2(\ANSWER/mem[8][3][9] ), .s(n16801), .op(
        n2919) );
  mux2_1 U16576 ( .ip1(n16333), .ip2(\ANSWER/mem[8][4][9] ), .s(n16803), .op(
        n2918) );
  mux2_1 U16577 ( .ip1(n16334), .ip2(\ANSWER/mem[8][5][9] ), .s(n16804), .op(
        n2917) );
  mux2_1 U16578 ( .ip1(n16333), .ip2(\ANSWER/mem[8][6][9] ), .s(n16805), .op(
        n2916) );
  mux2_1 U16579 ( .ip1(n16334), .ip2(\ANSWER/mem[8][7][9] ), .s(n16806), .op(
        n2915) );
  mux2_1 U16580 ( .ip1(n16333), .ip2(\ANSWER/mem[8][8][9] ), .s(n16807), .op(
        n2914) );
  mux2_1 U16581 ( .ip1(n16332), .ip2(\ANSWER/mem[8][9][9] ), .s(n16808), .op(
        n2913) );
  mux2_1 U16582 ( .ip1(n16334), .ip2(\ANSWER/mem[9][0][9] ), .s(n16809), .op(
        n2912) );
  mux2_1 U16583 ( .ip1(n16333), .ip2(\ANSWER/mem[9][1][9] ), .s(n16810), .op(
        n2911) );
  mux2_1 U16584 ( .ip1(n16334), .ip2(\ANSWER/mem[9][2][9] ), .s(n16811), .op(
        n2910) );
  mux2_1 U16585 ( .ip1(n16333), .ip2(\ANSWER/mem[9][3][9] ), .s(n16812), .op(
        n2909) );
  mux2_1 U16586 ( .ip1(n16334), .ip2(\ANSWER/mem[9][4][9] ), .s(n16813), .op(
        n2908) );
  mux2_1 U16587 ( .ip1(n16333), .ip2(\ANSWER/mem[9][5][9] ), .s(n16814), .op(
        n2907) );
  mux2_1 U16588 ( .ip1(n16334), .ip2(\ANSWER/mem[9][6][9] ), .s(n16815), .op(
        n2906) );
  mux2_1 U16589 ( .ip1(n16334), .ip2(\ANSWER/mem[9][7][9] ), .s(n16816), .op(
        n2905) );
  mux2_1 U16590 ( .ip1(n16334), .ip2(\ANSWER/mem[9][8][9] ), .s(n16817), .op(
        n2904) );
  mux2_1 U16591 ( .ip1(n16334), .ip2(\ANSWER/mem[9][9][9] ), .s(n16818), .op(
        n2903) );
  fulladder U16592 ( .a(n16337), .b(n16336), .ci(n16335), .co(n16401), .s(
        n16328) );
  fulladder U16593 ( .a(n16340), .b(n16339), .ci(n16338), .co(n16341), .s(
        n16287) );
  inv_1 U16594 ( .ip(n16341), .op(n16460) );
  or2_1 U16595 ( .ip1(n16342), .ip2(n16343), .op(n16346) );
  or2_1 U16596 ( .ip1(n16344), .ip2(n16343), .op(n16345) );
  nand2_1 U16597 ( .ip1(n16346), .ip2(n16345), .op(n16454) );
  nor3_1 U16598 ( .ip1(n16679), .ip2(n16678), .ip3(n16347), .op(n16412) );
  nor2_1 U16599 ( .ip1(n16679), .ip2(n16561), .op(n16511) );
  or2_1 U16600 ( .ip1(q_w2[12]), .ip2(n16511), .op(n16349) );
  or2_1 U16601 ( .ip1(m2DataIn[6]), .ip2(n16511), .op(n16348) );
  nand2_1 U16602 ( .ip1(n16349), .ip2(n16348), .op(n16410) );
  nor2_1 U16603 ( .ip1(n16412), .ip2(n16410), .op(n16350) );
  nand2_1 U16604 ( .ip1(m2DataIn[14]), .ip2(q_w2[4]), .op(n16409) );
  xor2_1 U16605 ( .ip1(n16350), .ip2(n16409), .op(n16453) );
  fulladder U16606 ( .a(n16353), .b(n16352), .ci(n16351), .co(n16452), .s(
        n16363) );
  nor2_1 U16607 ( .ip1(n16355), .ip2(n16354), .op(n16425) );
  nand2_1 U16608 ( .ip1(q_w2[8]), .ip2(m2DataIn[10]), .op(n16357) );
  nand2_1 U16609 ( .ip1(q_w2[10]), .ip2(m2DataIn[8]), .op(n16356) );
  xor2_1 U16610 ( .ip1(n16357), .ip2(n16356), .op(n16415) );
  mux2_1 U16611 ( .ip1(n16358), .ip2(rdata[10]), .s(n16415), .op(n16424) );
  fulladder U16612 ( .a(n16361), .b(n16360), .ci(n16359), .co(n16423), .s(
        n16364) );
  fulladder U16613 ( .a(n16364), .b(n16363), .ci(n16362), .co(n16429), .s(
        n16367) );
  fulladder U16614 ( .a(n16367), .b(n16366), .ci(n16365), .co(n16458), .s(
        n16336) );
  inv_1 U16615 ( .ip(q_w2[13]), .op(n16598) );
  nor2_1 U16616 ( .ip1(n16496), .ip2(n16598), .op(n16443) );
  nor2_1 U16617 ( .ip1(n16690), .ip2(n16552), .op(n16442) );
  nand2_1 U16618 ( .ip1(m2DataIn[15]), .ip2(q_w2[3]), .op(n16441) );
  inv_1 U16619 ( .ip(n16368), .op(n16408) );
  nand2_1 U16620 ( .ip1(m2DataIn[4]), .ip2(q_w2[14]), .op(n16434) );
  nor2_1 U16621 ( .ip1(n16369), .ip2(n16495), .op(n16433) );
  fulladder U16622 ( .a(n16418), .b(n16371), .ci(n16370), .co(n16406), .s(
        n16385) );
  fulladder U16623 ( .a(rdata[9]), .b(rdata[8]), .ci(n16372), .co(n16375), .s(
        n16263) );
  inv_1 U16624 ( .ip(n16375), .op(n16420) );
  nand2_1 U16625 ( .ip1(q_w2[6]), .ip2(m2DataIn[12]), .op(n16374) );
  nor2_1 U16626 ( .ip1(n16497), .ip2(n16510), .op(n16373) );
  xor2_1 U16627 ( .ip1(n16374), .ip2(n16373), .op(n16419) );
  mux2_1 U16628 ( .ip1(n16375), .ip2(n16420), .s(n16419), .op(n16428) );
  fulladder U16629 ( .a(n16378), .b(n16377), .ci(n16376), .co(n16379), .s(
        n16339) );
  inv_1 U16630 ( .ip(n16379), .op(n16427) );
  fulladder U16631 ( .a(n16382), .b(n16381), .ci(n16380), .co(n16426), .s(
        n16267) );
  fulladder U16632 ( .a(n16385), .b(n16384), .ci(n16383), .co(n16455), .s(
        n16387) );
  fulladder U16633 ( .a(n16388), .b(n16387), .ci(n16386), .co(n16461), .s(
        n16337) );
  or2_1 U16634 ( .ip1(n16390), .ip2(n16389), .op(n16391) );
  nand2_1 U16635 ( .ip1(n16392), .ip2(n16391), .op(n16393) );
  nor2_1 U16636 ( .ip1(n16394), .ip2(n16393), .op(n16402) );
  inv_1 U16637 ( .ip(n16402), .op(n16395) );
  nand2_1 U16638 ( .ip1(n16394), .ip2(n16393), .op(n16405) );
  nand2_1 U16639 ( .ip1(n16395), .ip2(n16405), .op(n16397) );
  nor2_1 U16640 ( .ip1(n16401), .ip2(n16397), .op(n16396) );
  not_ab_or_c_or_d U16641 ( .ip1(n16401), .ip2(n16397), .ip3(n16714), .ip4(
        n16396), .op(n16399) );
  buf_1 U16642 ( .ip(n16399), .op(n16398) );
  mux2_1 U16643 ( .ip1(n16398), .ip2(\ANSWER/mem[0][0][10] ), .s(n16717), .op(
        n2902) );
  mux2_1 U16644 ( .ip1(n16398), .ip2(\ANSWER/mem[0][1][10] ), .s(n16718), .op(
        n2901) );
  mux2_1 U16645 ( .ip1(n16398), .ip2(\ANSWER/mem[0][2][10] ), .s(n16719), .op(
        n2900) );
  mux2_1 U16646 ( .ip1(n16398), .ip2(\ANSWER/mem[0][3][10] ), .s(n16720), .op(
        n2899) );
  mux2_1 U16647 ( .ip1(n16398), .ip2(\ANSWER/mem[0][4][10] ), .s(n16721), .op(
        n2898) );
  mux2_1 U16648 ( .ip1(n16398), .ip2(\ANSWER/mem[0][5][10] ), .s(n16722), .op(
        n2897) );
  mux2_1 U16649 ( .ip1(n16398), .ip2(\ANSWER/mem[0][6][10] ), .s(n16723), .op(
        n2896) );
  mux2_1 U16650 ( .ip1(n16398), .ip2(\ANSWER/mem[0][7][10] ), .s(n16724), .op(
        n2895) );
  mux2_1 U16651 ( .ip1(n16398), .ip2(\ANSWER/mem[0][8][10] ), .s(n16725), .op(
        n2894) );
  mux2_1 U16652 ( .ip1(n16398), .ip2(\ANSWER/mem[0][9][10] ), .s(n16726), .op(
        n2893) );
  mux2_1 U16653 ( .ip1(n16398), .ip2(\ANSWER/mem[1][0][10] ), .s(n16727), .op(
        n2892) );
  mux2_1 U16654 ( .ip1(n16398), .ip2(\ANSWER/mem[1][1][10] ), .s(n16728), .op(
        n2891) );
  mux2_1 U16655 ( .ip1(n16398), .ip2(\ANSWER/mem[1][2][10] ), .s(n16729), .op(
        n2890) );
  mux2_1 U16656 ( .ip1(n16398), .ip2(\ANSWER/mem[1][3][10] ), .s(n16730), .op(
        n2889) );
  mux2_1 U16657 ( .ip1(n16398), .ip2(\ANSWER/mem[1][4][10] ), .s(n16731), .op(
        n2888) );
  mux2_1 U16658 ( .ip1(n16398), .ip2(\ANSWER/mem[1][5][10] ), .s(n16732), .op(
        n2887) );
  mux2_1 U16659 ( .ip1(n16398), .ip2(\ANSWER/mem[1][6][10] ), .s(n16733), .op(
        n2886) );
  mux2_1 U16660 ( .ip1(n16398), .ip2(\ANSWER/mem[1][7][10] ), .s(n16734), .op(
        n2885) );
  mux2_1 U16661 ( .ip1(n16398), .ip2(\ANSWER/mem[1][8][10] ), .s(n16735), .op(
        n2884) );
  mux2_1 U16662 ( .ip1(n16398), .ip2(\ANSWER/mem[1][9][10] ), .s(n16736), .op(
        n2883) );
  mux2_1 U16663 ( .ip1(n16398), .ip2(\ANSWER/mem[2][0][10] ), .s(n16737), .op(
        n2882) );
  mux2_1 U16664 ( .ip1(n16398), .ip2(\ANSWER/mem[2][1][10] ), .s(n16738), .op(
        n2881) );
  mux2_1 U16665 ( .ip1(n16398), .ip2(\ANSWER/mem[2][2][10] ), .s(n16739), .op(
        n2880) );
  mux2_1 U16666 ( .ip1(n16398), .ip2(\ANSWER/mem[2][3][10] ), .s(n16740), .op(
        n2879) );
  mux2_1 U16667 ( .ip1(n16398), .ip2(\ANSWER/mem[2][4][10] ), .s(n16741), .op(
        n2878) );
  mux2_1 U16668 ( .ip1(n16398), .ip2(\ANSWER/mem[2][5][10] ), .s(n16742), .op(
        n2877) );
  mux2_1 U16669 ( .ip1(n16398), .ip2(\ANSWER/mem[2][6][10] ), .s(n16743), .op(
        n2876) );
  mux2_1 U16670 ( .ip1(n16398), .ip2(\ANSWER/mem[2][7][10] ), .s(n16744), .op(
        n2875) );
  mux2_1 U16671 ( .ip1(n16398), .ip2(\ANSWER/mem[2][8][10] ), .s(n16745), .op(
        n2874) );
  mux2_1 U16672 ( .ip1(n16398), .ip2(\ANSWER/mem[2][9][10] ), .s(n16746), .op(
        n2873) );
  mux2_1 U16673 ( .ip1(n16398), .ip2(\ANSWER/mem[3][0][10] ), .s(n16747), .op(
        n2872) );
  mux2_1 U16674 ( .ip1(n16398), .ip2(\ANSWER/mem[3][1][10] ), .s(n16748), .op(
        n2871) );
  mux2_1 U16675 ( .ip1(n16398), .ip2(\ANSWER/mem[3][2][10] ), .s(n16749), .op(
        n2870) );
  mux2_1 U16676 ( .ip1(n16398), .ip2(\ANSWER/mem[3][3][10] ), .s(n16750), .op(
        n2869) );
  mux2_1 U16677 ( .ip1(n16398), .ip2(\ANSWER/mem[3][4][10] ), .s(n16751), .op(
        n2868) );
  mux2_1 U16678 ( .ip1(n16398), .ip2(\ANSWER/mem[3][5][10] ), .s(n16752), .op(
        n2867) );
  mux2_1 U16679 ( .ip1(n16400), .ip2(\ANSWER/mem[3][6][10] ), .s(n16753), .op(
        n2866) );
  mux2_1 U16680 ( .ip1(n16400), .ip2(\ANSWER/mem[3][7][10] ), .s(n16754), .op(
        n2865) );
  mux2_1 U16681 ( .ip1(n16400), .ip2(\ANSWER/mem[3][8][10] ), .s(n16755), .op(
        n2864) );
  mux2_1 U16682 ( .ip1(n16400), .ip2(\ANSWER/mem[3][9][10] ), .s(n16756), .op(
        n2863) );
  mux2_1 U16683 ( .ip1(n16399), .ip2(\ANSWER/mem[4][0][10] ), .s(n16757), .op(
        n2862) );
  mux2_1 U16684 ( .ip1(n16399), .ip2(\ANSWER/mem[4][1][10] ), .s(n16758), .op(
        n2861) );
  mux2_1 U16685 ( .ip1(n16399), .ip2(\ANSWER/mem[4][2][10] ), .s(n16759), .op(
        n2860) );
  mux2_1 U16686 ( .ip1(n16399), .ip2(\ANSWER/mem[4][3][10] ), .s(n16760), .op(
        n2859) );
  mux2_1 U16687 ( .ip1(n16400), .ip2(\ANSWER/mem[4][4][10] ), .s(n16761), .op(
        n2858) );
  mux2_1 U16688 ( .ip1(n16400), .ip2(\ANSWER/mem[4][5][10] ), .s(n16762), .op(
        n2857) );
  mux2_1 U16689 ( .ip1(n16400), .ip2(\ANSWER/mem[4][6][10] ), .s(n16763), .op(
        n2856) );
  mux2_1 U16690 ( .ip1(n16400), .ip2(\ANSWER/mem[4][7][10] ), .s(n16764), .op(
        n2855) );
  mux2_1 U16691 ( .ip1(n16400), .ip2(\ANSWER/mem[4][8][10] ), .s(n16765), .op(
        n2854) );
  mux2_1 U16692 ( .ip1(n16400), .ip2(\ANSWER/mem[4][9][10] ), .s(n16766), .op(
        n2853) );
  mux2_1 U16693 ( .ip1(n16400), .ip2(\ANSWER/mem[5][0][10] ), .s(n16767), .op(
        n2852) );
  mux2_1 U16694 ( .ip1(n16399), .ip2(\ANSWER/mem[5][1][10] ), .s(n16768), .op(
        n2851) );
  mux2_1 U16695 ( .ip1(n16400), .ip2(\ANSWER/mem[5][2][10] ), .s(n16769), .op(
        n2850) );
  mux2_1 U16696 ( .ip1(n16399), .ip2(\ANSWER/mem[5][3][10] ), .s(n16770), .op(
        n2849) );
  mux2_1 U16697 ( .ip1(n16400), .ip2(\ANSWER/mem[5][4][10] ), .s(n16771), .op(
        n2848) );
  mux2_1 U16698 ( .ip1(n16399), .ip2(\ANSWER/mem[5][5][10] ), .s(n16772), .op(
        n2847) );
  mux2_1 U16699 ( .ip1(n16399), .ip2(\ANSWER/mem[5][6][10] ), .s(n16773), .op(
        n2846) );
  mux2_1 U16700 ( .ip1(n16399), .ip2(\ANSWER/mem[5][7][10] ), .s(n16774), .op(
        n2845) );
  mux2_1 U16701 ( .ip1(n16399), .ip2(\ANSWER/mem[5][8][10] ), .s(n16775), .op(
        n2844) );
  mux2_1 U16702 ( .ip1(n16399), .ip2(\ANSWER/mem[5][9][10] ), .s(n16776), .op(
        n2843) );
  mux2_1 U16703 ( .ip1(n16399), .ip2(\ANSWER/mem[6][0][10] ), .s(n16777), .op(
        n2842) );
  mux2_1 U16704 ( .ip1(n16399), .ip2(\ANSWER/mem[6][1][10] ), .s(n16778), .op(
        n2841) );
  mux2_1 U16705 ( .ip1(n16399), .ip2(\ANSWER/mem[6][2][10] ), .s(n16779), .op(
        n2840) );
  mux2_1 U16706 ( .ip1(n16399), .ip2(\ANSWER/mem[6][3][10] ), .s(n16780), .op(
        n2839) );
  mux2_1 U16707 ( .ip1(n16399), .ip2(\ANSWER/mem[6][4][10] ), .s(n16781), .op(
        n2838) );
  mux2_1 U16708 ( .ip1(n16399), .ip2(\ANSWER/mem[6][5][10] ), .s(n16782), .op(
        n2837) );
  mux2_1 U16709 ( .ip1(n16399), .ip2(\ANSWER/mem[6][6][10] ), .s(n16783), .op(
        n2836) );
  mux2_1 U16710 ( .ip1(n16399), .ip2(\ANSWER/mem[6][7][10] ), .s(n16784), .op(
        n2835) );
  mux2_1 U16711 ( .ip1(n16399), .ip2(\ANSWER/mem[6][8][10] ), .s(n16785), .op(
        n2834) );
  mux2_1 U16712 ( .ip1(n16399), .ip2(\ANSWER/mem[6][9][10] ), .s(n16786), .op(
        n2833) );
  mux2_1 U16713 ( .ip1(n16399), .ip2(\ANSWER/mem[7][0][10] ), .s(n16787), .op(
        n2832) );
  mux2_1 U16714 ( .ip1(n16399), .ip2(\ANSWER/mem[7][1][10] ), .s(n16788), .op(
        n2831) );
  buf_1 U16715 ( .ip(n16399), .op(n16400) );
  mux2_1 U16716 ( .ip1(n16400), .ip2(\ANSWER/mem[7][2][10] ), .s(n16790), .op(
        n2830) );
  mux2_1 U16717 ( .ip1(n16400), .ip2(\ANSWER/mem[7][3][10] ), .s(n16791), .op(
        n2829) );
  mux2_1 U16718 ( .ip1(n16399), .ip2(\ANSWER/mem[7][4][10] ), .s(n16792), .op(
        n2828) );
  mux2_1 U16719 ( .ip1(n16399), .ip2(\ANSWER/mem[7][5][10] ), .s(n16793), .op(
        n2827) );
  mux2_1 U16720 ( .ip1(n16400), .ip2(\ANSWER/mem[7][6][10] ), .s(n16794), .op(
        n2826) );
  mux2_1 U16721 ( .ip1(n16400), .ip2(\ANSWER/mem[7][7][10] ), .s(n16795), .op(
        n2825) );
  mux2_1 U16722 ( .ip1(n16400), .ip2(\ANSWER/mem[7][8][10] ), .s(n16796), .op(
        n2824) );
  mux2_1 U16723 ( .ip1(n16400), .ip2(\ANSWER/mem[7][9][10] ), .s(n16797), .op(
        n2823) );
  mux2_1 U16724 ( .ip1(n16400), .ip2(\ANSWER/mem[8][0][10] ), .s(n16798), .op(
        n2822) );
  mux2_1 U16725 ( .ip1(n16400), .ip2(\ANSWER/mem[8][1][10] ), .s(n16799), .op(
        n2821) );
  mux2_1 U16726 ( .ip1(n16400), .ip2(\ANSWER/mem[8][2][10] ), .s(n16800), .op(
        n2820) );
  mux2_1 U16727 ( .ip1(n16400), .ip2(\ANSWER/mem[8][3][10] ), .s(n16801), .op(
        n2819) );
  mux2_1 U16728 ( .ip1(n16399), .ip2(\ANSWER/mem[8][4][10] ), .s(n16803), .op(
        n2818) );
  mux2_1 U16729 ( .ip1(n16399), .ip2(\ANSWER/mem[8][5][10] ), .s(n16804), .op(
        n2817) );
  mux2_1 U16730 ( .ip1(n16399), .ip2(\ANSWER/mem[8][6][10] ), .s(n16805), .op(
        n2816) );
  mux2_1 U16731 ( .ip1(n16399), .ip2(\ANSWER/mem[8][7][10] ), .s(n16806), .op(
        n2815) );
  mux2_1 U16732 ( .ip1(n16399), .ip2(\ANSWER/mem[8][8][10] ), .s(n16807), .op(
        n2814) );
  mux2_1 U16733 ( .ip1(n16399), .ip2(\ANSWER/mem[8][9][10] ), .s(n16808), .op(
        n2813) );
  mux2_1 U16734 ( .ip1(n16399), .ip2(\ANSWER/mem[9][0][10] ), .s(n16809), .op(
        n2812) );
  mux2_1 U16735 ( .ip1(n16399), .ip2(\ANSWER/mem[9][1][10] ), .s(n16810), .op(
        n2811) );
  mux2_1 U16736 ( .ip1(n16399), .ip2(\ANSWER/mem[9][2][10] ), .s(n16811), .op(
        n2810) );
  mux2_1 U16737 ( .ip1(n16399), .ip2(\ANSWER/mem[9][3][10] ), .s(n16812), .op(
        n2809) );
  mux2_1 U16738 ( .ip1(n16399), .ip2(\ANSWER/mem[9][4][10] ), .s(n16813), .op(
        n2808) );
  mux2_1 U16739 ( .ip1(n16399), .ip2(\ANSWER/mem[9][5][10] ), .s(n16814), .op(
        n2807) );
  mux2_1 U16740 ( .ip1(n16400), .ip2(\ANSWER/mem[9][6][10] ), .s(n16815), .op(
        n2806) );
  mux2_1 U16741 ( .ip1(n16400), .ip2(\ANSWER/mem[9][7][10] ), .s(n16816), .op(
        n2805) );
  mux2_1 U16742 ( .ip1(n16400), .ip2(\ANSWER/mem[9][8][10] ), .s(n16817), .op(
        n2804) );
  mux2_1 U16743 ( .ip1(n16400), .ip2(\ANSWER/mem[9][9][10] ), .s(n16818), .op(
        n2803) );
  inv_1 U16744 ( .ip(n16401), .op(n16403) );
  or2_1 U16745 ( .ip1(n16403), .ip2(n16402), .op(n16404) );
  nand2_1 U16746 ( .ip1(n16405), .ip2(n16404), .op(n16525) );
  fulladder U16747 ( .a(n16408), .b(n16407), .ci(n16406), .co(n16494), .s(
        n16457) );
  nor2_1 U16748 ( .ip1(n16410), .ip2(n16409), .op(n16411) );
  nor2_1 U16749 ( .ip1(n16412), .ip2(n16411), .op(n16501) );
  nand2_1 U16750 ( .ip1(m2DataIn[13]), .ip2(q_w2[6]), .op(n16500) );
  nor2_1 U16751 ( .ip1(n16600), .ip2(n16622), .op(n16541) );
  and2_1 U16752 ( .ip1(n16541), .ip2(n16413), .op(n16414) );
  or2_1 U16753 ( .ip1(rdata[10]), .ip2(n16414), .op(n16417) );
  or2_1 U16754 ( .ip1(n16415), .ip2(n16414), .op(n16416) );
  nand2_1 U16755 ( .ip1(n16417), .ip2(n16416), .op(n16499) );
  nor2_1 U16756 ( .ip1(n16500), .ip2(n16418), .op(n16422) );
  nor2_1 U16757 ( .ip1(n16420), .ip2(n16419), .op(n16421) );
  nor2_1 U16758 ( .ip1(n16422), .ip2(n16421), .op(n16518) );
  fulladder U16759 ( .a(n16425), .b(n16424), .ci(n16423), .co(n16517), .s(
        n16430) );
  fulladder U16760 ( .a(n16428), .b(n16427), .ci(n16426), .co(n16492), .s(
        n16456) );
  fulladder U16761 ( .a(n16431), .b(n16430), .ci(n16429), .co(n16522), .s(
        n16459) );
  fulladder U16762 ( .a(n16434), .b(n16433), .ci(n16432), .co(n16435), .s(
        n16407) );
  inv_1 U16763 ( .ip(n16435), .op(n16487) );
  inv_1 U16764 ( .ip(rdata[11]), .op(n16440) );
  nand2_1 U16765 ( .ip1(m2DataIn[9]), .ip2(q_w2[10]), .op(n16436) );
  and2_1 U16766 ( .ip1(n16541), .ip2(n16442), .op(n16477) );
  or2_1 U16767 ( .ip1(n16436), .ip2(n16477), .op(n16439) );
  nand2_1 U16768 ( .ip1(m2DataIn[10]), .ip2(q_w2[9]), .op(n16437) );
  or2_1 U16769 ( .ip1(n16437), .ip2(n16477), .op(n16438) );
  nand2_1 U16770 ( .ip1(n16439), .ip2(n16438), .op(n16478) );
  mux2_1 U16771 ( .ip1(rdata[11]), .ip2(n16440), .s(n16478), .op(n16486) );
  fulladder U16772 ( .a(n16443), .b(n16442), .ci(n16441), .co(n16485), .s(
        n16368) );
  inv_1 U16773 ( .ip(n16444), .op(n16491) );
  nor2_1 U16774 ( .ip1(n16445), .ip2(n16495), .op(n16516) );
  nand2_1 U16775 ( .ip1(m2DataIn[7]), .ip2(q_w2[12]), .op(n16515) );
  nand2_1 U16776 ( .ip1(m2DataIn[5]), .ip2(q_w2[14]), .op(n16514) );
  inv_1 U16777 ( .ip(n16446), .op(n16484) );
  nand2_1 U16778 ( .ip1(m2DataIn[6]), .ip2(q_w2[13]), .op(n16476) );
  nor2_1 U16779 ( .ip1(n16498), .ip2(n16447), .op(n16475) );
  nand2_1 U16780 ( .ip1(m2DataIn[8]), .ip2(q_w2[11]), .op(n16474) );
  inv_1 U16781 ( .ip(n16448), .op(n16483) );
  nand2_1 U16782 ( .ip1(q_w2[7]), .ip2(m2DataIn[12]), .op(n16450) );
  nand2_1 U16783 ( .ip1(q_w2[8]), .ip2(m2DataIn[11]), .op(n16449) );
  xor2_1 U16784 ( .ip1(n16450), .ip2(n16449), .op(n16503) );
  nor2_1 U16785 ( .ip1(n16597), .ip2(n16497), .op(n16505) );
  xor2_1 U16786 ( .ip1(n16503), .ip2(n16505), .op(n16482) );
  inv_1 U16787 ( .ip(n16451), .op(n16490) );
  fulladder U16788 ( .a(n16454), .b(n16453), .ci(n16452), .co(n16489), .s(
        n16431) );
  fulladder U16789 ( .a(n16457), .b(n16456), .ci(n16455), .co(n16520), .s(
        n16462) );
  fulladder U16790 ( .a(n16460), .b(n16459), .ci(n16458), .co(n16468), .s(
        n16463) );
  fulladder U16791 ( .a(n16463), .b(n16462), .ci(n16461), .co(n16523), .s(
        n16394) );
  nor2_1 U16792 ( .ip1(n16714), .ip2(n16464), .op(n16466) );
  buf_1 U16793 ( .ip(n16466), .op(n16465) );
  mux2_1 U16794 ( .ip1(n16465), .ip2(\ANSWER/mem[0][0][11] ), .s(n16717), .op(
        n2802) );
  mux2_1 U16795 ( .ip1(n16465), .ip2(\ANSWER/mem[0][1][11] ), .s(n16718), .op(
        n2801) );
  mux2_1 U16796 ( .ip1(n16465), .ip2(\ANSWER/mem[0][2][11] ), .s(n16719), .op(
        n2800) );
  mux2_1 U16797 ( .ip1(n16465), .ip2(\ANSWER/mem[0][3][11] ), .s(n16720), .op(
        n2799) );
  mux2_1 U16798 ( .ip1(n16465), .ip2(\ANSWER/mem[0][4][11] ), .s(n16721), .op(
        n2798) );
  mux2_1 U16799 ( .ip1(n16465), .ip2(\ANSWER/mem[0][5][11] ), .s(n16722), .op(
        n2797) );
  mux2_1 U16800 ( .ip1(n16465), .ip2(\ANSWER/mem[0][6][11] ), .s(n16723), .op(
        n2796) );
  mux2_1 U16801 ( .ip1(n16465), .ip2(\ANSWER/mem[0][7][11] ), .s(n16724), .op(
        n2795) );
  mux2_1 U16802 ( .ip1(n16465), .ip2(\ANSWER/mem[0][8][11] ), .s(n16725), .op(
        n2794) );
  mux2_1 U16803 ( .ip1(n16465), .ip2(\ANSWER/mem[0][9][11] ), .s(n16726), .op(
        n2793) );
  mux2_1 U16804 ( .ip1(n16465), .ip2(\ANSWER/mem[1][0][11] ), .s(n16727), .op(
        n2792) );
  mux2_1 U16805 ( .ip1(n16465), .ip2(\ANSWER/mem[1][1][11] ), .s(n16728), .op(
        n2791) );
  mux2_1 U16806 ( .ip1(n16465), .ip2(\ANSWER/mem[1][2][11] ), .s(n16729), .op(
        n2790) );
  mux2_1 U16807 ( .ip1(n16465), .ip2(\ANSWER/mem[1][3][11] ), .s(n16730), .op(
        n2789) );
  mux2_1 U16808 ( .ip1(n16465), .ip2(\ANSWER/mem[1][4][11] ), .s(n16731), .op(
        n2788) );
  mux2_1 U16809 ( .ip1(n16465), .ip2(\ANSWER/mem[1][5][11] ), .s(n16732), .op(
        n2787) );
  mux2_1 U16810 ( .ip1(n16465), .ip2(\ANSWER/mem[1][6][11] ), .s(n16733), .op(
        n2786) );
  mux2_1 U16811 ( .ip1(n16465), .ip2(\ANSWER/mem[1][7][11] ), .s(n16734), .op(
        n2785) );
  mux2_1 U16812 ( .ip1(n16465), .ip2(\ANSWER/mem[1][8][11] ), .s(n16735), .op(
        n2784) );
  mux2_1 U16813 ( .ip1(n16465), .ip2(\ANSWER/mem[1][9][11] ), .s(n16736), .op(
        n2783) );
  mux2_1 U16814 ( .ip1(n16465), .ip2(\ANSWER/mem[2][0][11] ), .s(n16737), .op(
        n2782) );
  mux2_1 U16815 ( .ip1(n16465), .ip2(\ANSWER/mem[2][1][11] ), .s(n16738), .op(
        n2781) );
  mux2_1 U16816 ( .ip1(n16465), .ip2(\ANSWER/mem[2][2][11] ), .s(n16739), .op(
        n2780) );
  mux2_1 U16817 ( .ip1(n16465), .ip2(\ANSWER/mem[2][3][11] ), .s(n16740), .op(
        n2779) );
  mux2_1 U16818 ( .ip1(n16465), .ip2(\ANSWER/mem[2][4][11] ), .s(n16741), .op(
        n2778) );
  mux2_1 U16819 ( .ip1(n16465), .ip2(\ANSWER/mem[2][5][11] ), .s(n16742), .op(
        n2777) );
  mux2_1 U16820 ( .ip1(n16465), .ip2(\ANSWER/mem[2][6][11] ), .s(n16743), .op(
        n2776) );
  mux2_1 U16821 ( .ip1(n16465), .ip2(\ANSWER/mem[2][7][11] ), .s(n16744), .op(
        n2775) );
  mux2_1 U16822 ( .ip1(n16465), .ip2(\ANSWER/mem[2][8][11] ), .s(n16745), .op(
        n2774) );
  mux2_1 U16823 ( .ip1(n16465), .ip2(\ANSWER/mem[2][9][11] ), .s(n16746), .op(
        n2773) );
  mux2_1 U16824 ( .ip1(n16465), .ip2(\ANSWER/mem[3][0][11] ), .s(n16747), .op(
        n2772) );
  mux2_1 U16825 ( .ip1(n16465), .ip2(\ANSWER/mem[3][1][11] ), .s(n16748), .op(
        n2771) );
  mux2_1 U16826 ( .ip1(n16465), .ip2(\ANSWER/mem[3][2][11] ), .s(n16749), .op(
        n2770) );
  mux2_1 U16827 ( .ip1(n16465), .ip2(\ANSWER/mem[3][3][11] ), .s(n16750), .op(
        n2769) );
  mux2_1 U16828 ( .ip1(n16465), .ip2(\ANSWER/mem[3][4][11] ), .s(n16751), .op(
        n2768) );
  mux2_1 U16829 ( .ip1(n16465), .ip2(\ANSWER/mem[3][5][11] ), .s(n16752), .op(
        n2767) );
  mux2_1 U16830 ( .ip1(n16467), .ip2(\ANSWER/mem[3][6][11] ), .s(n16753), .op(
        n2766) );
  mux2_1 U16831 ( .ip1(n16467), .ip2(\ANSWER/mem[3][7][11] ), .s(n16754), .op(
        n2765) );
  mux2_1 U16832 ( .ip1(n16467), .ip2(\ANSWER/mem[3][8][11] ), .s(n16755), .op(
        n2764) );
  mux2_1 U16833 ( .ip1(n16467), .ip2(\ANSWER/mem[3][9][11] ), .s(n16756), .op(
        n2763) );
  mux2_1 U16834 ( .ip1(n16466), .ip2(\ANSWER/mem[4][0][11] ), .s(n16757), .op(
        n2762) );
  mux2_1 U16835 ( .ip1(n16466), .ip2(\ANSWER/mem[4][1][11] ), .s(n16758), .op(
        n2761) );
  mux2_1 U16836 ( .ip1(n16466), .ip2(\ANSWER/mem[4][2][11] ), .s(n16759), .op(
        n2760) );
  mux2_1 U16837 ( .ip1(n16466), .ip2(\ANSWER/mem[4][3][11] ), .s(n16760), .op(
        n2759) );
  mux2_1 U16838 ( .ip1(n16467), .ip2(\ANSWER/mem[4][4][11] ), .s(n16761), .op(
        n2758) );
  mux2_1 U16839 ( .ip1(n16467), .ip2(\ANSWER/mem[4][5][11] ), .s(n16762), .op(
        n2757) );
  mux2_1 U16840 ( .ip1(n16467), .ip2(\ANSWER/mem[4][6][11] ), .s(n16763), .op(
        n2756) );
  mux2_1 U16841 ( .ip1(n16467), .ip2(\ANSWER/mem[4][7][11] ), .s(n16764), .op(
        n2755) );
  mux2_1 U16842 ( .ip1(n16467), .ip2(\ANSWER/mem[4][8][11] ), .s(n16765), .op(
        n2754) );
  mux2_1 U16843 ( .ip1(n16467), .ip2(\ANSWER/mem[4][9][11] ), .s(n16766), .op(
        n2753) );
  mux2_1 U16844 ( .ip1(n16467), .ip2(\ANSWER/mem[5][0][11] ), .s(n16767), .op(
        n2752) );
  mux2_1 U16845 ( .ip1(n16466), .ip2(\ANSWER/mem[5][1][11] ), .s(n16768), .op(
        n2751) );
  mux2_1 U16846 ( .ip1(n16467), .ip2(\ANSWER/mem[5][2][11] ), .s(n16769), .op(
        n2750) );
  mux2_1 U16847 ( .ip1(n16466), .ip2(\ANSWER/mem[5][3][11] ), .s(n16770), .op(
        n2749) );
  mux2_1 U16848 ( .ip1(n16467), .ip2(\ANSWER/mem[5][4][11] ), .s(n16771), .op(
        n2748) );
  mux2_1 U16849 ( .ip1(n16466), .ip2(\ANSWER/mem[5][5][11] ), .s(n16772), .op(
        n2747) );
  mux2_1 U16850 ( .ip1(n16466), .ip2(\ANSWER/mem[5][6][11] ), .s(n16773), .op(
        n2746) );
  mux2_1 U16851 ( .ip1(n16466), .ip2(\ANSWER/mem[5][7][11] ), .s(n16774), .op(
        n2745) );
  mux2_1 U16852 ( .ip1(n16466), .ip2(\ANSWER/mem[5][8][11] ), .s(n16775), .op(
        n2744) );
  mux2_1 U16853 ( .ip1(n16466), .ip2(\ANSWER/mem[5][9][11] ), .s(n16776), .op(
        n2743) );
  mux2_1 U16854 ( .ip1(n16466), .ip2(\ANSWER/mem[6][0][11] ), .s(n16777), .op(
        n2742) );
  mux2_1 U16855 ( .ip1(n16466), .ip2(\ANSWER/mem[6][1][11] ), .s(n16778), .op(
        n2741) );
  mux2_1 U16856 ( .ip1(n16466), .ip2(\ANSWER/mem[6][2][11] ), .s(n16779), .op(
        n2740) );
  mux2_1 U16857 ( .ip1(n16466), .ip2(\ANSWER/mem[6][3][11] ), .s(n16780), .op(
        n2739) );
  mux2_1 U16858 ( .ip1(n16466), .ip2(\ANSWER/mem[6][4][11] ), .s(n16781), .op(
        n2738) );
  mux2_1 U16859 ( .ip1(n16466), .ip2(\ANSWER/mem[6][5][11] ), .s(n16782), .op(
        n2737) );
  mux2_1 U16860 ( .ip1(n16466), .ip2(\ANSWER/mem[6][6][11] ), .s(n16783), .op(
        n2736) );
  mux2_1 U16861 ( .ip1(n16466), .ip2(\ANSWER/mem[6][7][11] ), .s(n16784), .op(
        n2735) );
  mux2_1 U16862 ( .ip1(n16466), .ip2(\ANSWER/mem[6][8][11] ), .s(n16785), .op(
        n2734) );
  mux2_1 U16863 ( .ip1(n16466), .ip2(\ANSWER/mem[6][9][11] ), .s(n16786), .op(
        n2733) );
  mux2_1 U16864 ( .ip1(n16466), .ip2(\ANSWER/mem[7][0][11] ), .s(n16787), .op(
        n2732) );
  mux2_1 U16865 ( .ip1(n16466), .ip2(\ANSWER/mem[7][1][11] ), .s(n16788), .op(
        n2731) );
  buf_1 U16866 ( .ip(n16466), .op(n16467) );
  mux2_1 U16867 ( .ip1(n16467), .ip2(\ANSWER/mem[7][2][11] ), .s(n16790), .op(
        n2730) );
  mux2_1 U16868 ( .ip1(n16467), .ip2(\ANSWER/mem[7][3][11] ), .s(n16791), .op(
        n2729) );
  mux2_1 U16869 ( .ip1(n16467), .ip2(\ANSWER/mem[7][4][11] ), .s(n16792), .op(
        n2728) );
  mux2_1 U16870 ( .ip1(n16466), .ip2(\ANSWER/mem[7][5][11] ), .s(n16793), .op(
        n2727) );
  mux2_1 U16871 ( .ip1(n16466), .ip2(\ANSWER/mem[7][6][11] ), .s(n16794), .op(
        n2726) );
  mux2_1 U16872 ( .ip1(n16467), .ip2(\ANSWER/mem[7][7][11] ), .s(n16795), .op(
        n2725) );
  mux2_1 U16873 ( .ip1(n16467), .ip2(\ANSWER/mem[7][8][11] ), .s(n16796), .op(
        n2724) );
  mux2_1 U16874 ( .ip1(n16467), .ip2(\ANSWER/mem[7][9][11] ), .s(n16797), .op(
        n2723) );
  mux2_1 U16875 ( .ip1(n16467), .ip2(\ANSWER/mem[8][0][11] ), .s(n16798), .op(
        n2722) );
  mux2_1 U16876 ( .ip1(n16467), .ip2(\ANSWER/mem[8][1][11] ), .s(n16799), .op(
        n2721) );
  mux2_1 U16877 ( .ip1(n16467), .ip2(\ANSWER/mem[8][2][11] ), .s(n16800), .op(
        n2720) );
  mux2_1 U16878 ( .ip1(n16467), .ip2(\ANSWER/mem[8][3][11] ), .s(n16801), .op(
        n2719) );
  mux2_1 U16879 ( .ip1(n16466), .ip2(\ANSWER/mem[8][4][11] ), .s(n16803), .op(
        n2718) );
  mux2_1 U16880 ( .ip1(n16466), .ip2(\ANSWER/mem[8][5][11] ), .s(n16804), .op(
        n2717) );
  mux2_1 U16881 ( .ip1(n16466), .ip2(\ANSWER/mem[8][6][11] ), .s(n16805), .op(
        n2716) );
  mux2_1 U16882 ( .ip1(n16466), .ip2(\ANSWER/mem[8][7][11] ), .s(n16806), .op(
        n2715) );
  mux2_1 U16883 ( .ip1(n16466), .ip2(\ANSWER/mem[8][8][11] ), .s(n16807), .op(
        n2714) );
  mux2_1 U16884 ( .ip1(n16466), .ip2(\ANSWER/mem[8][9][11] ), .s(n16808), .op(
        n2713) );
  mux2_1 U16885 ( .ip1(n16466), .ip2(\ANSWER/mem[9][0][11] ), .s(n16809), .op(
        n2712) );
  mux2_1 U16886 ( .ip1(n16466), .ip2(\ANSWER/mem[9][1][11] ), .s(n16810), .op(
        n2711) );
  mux2_1 U16887 ( .ip1(n16466), .ip2(\ANSWER/mem[9][2][11] ), .s(n16811), .op(
        n2710) );
  mux2_1 U16888 ( .ip1(n16466), .ip2(\ANSWER/mem[9][3][11] ), .s(n16812), .op(
        n2709) );
  mux2_1 U16889 ( .ip1(n16466), .ip2(\ANSWER/mem[9][4][11] ), .s(n16813), .op(
        n2708) );
  mux2_1 U16890 ( .ip1(n16466), .ip2(\ANSWER/mem[9][5][11] ), .s(n16814), .op(
        n2707) );
  mux2_1 U16891 ( .ip1(n16467), .ip2(\ANSWER/mem[9][6][11] ), .s(n16815), .op(
        n2706) );
  mux2_1 U16892 ( .ip1(n16467), .ip2(\ANSWER/mem[9][7][11] ), .s(n16816), .op(
        n2705) );
  mux2_1 U16893 ( .ip1(n16467), .ip2(\ANSWER/mem[9][8][11] ), .s(n16817), .op(
        n2704) );
  mux2_1 U16894 ( .ip1(n16467), .ip2(\ANSWER/mem[9][9][11] ), .s(n16818), .op(
        n2703) );
  fulladder U16895 ( .a(n16470), .b(n16469), .ci(n16468), .co(n16585), .s(
        n16524) );
  inv_1 U16896 ( .ip(rdata[12]), .op(n16565) );
  nand2_1 U16897 ( .ip1(m2DataIn[10]), .ip2(q_w2[11]), .op(n16677) );
  nor3_1 U16898 ( .ip1(n16690), .ip2(n16622), .ip3(n16677), .op(n16567) );
  or2_1 U16899 ( .ip1(q_w2[11]), .ip2(n16541), .op(n16472) );
  or2_1 U16900 ( .ip1(m2DataIn[9]), .ip2(n16541), .op(n16471) );
  nand2_1 U16901 ( .ip1(n16472), .ip2(n16471), .op(n16473) );
  or2_1 U16902 ( .ip1(n16567), .ip2(n16473), .op(n16564) );
  mux2_1 U16903 ( .ip1(rdata[12]), .ip2(n16565), .s(n16564), .op(n16571) );
  fulladder U16904 ( .a(n16476), .b(n16475), .ci(n16474), .co(n16570), .s(
        n16448) );
  or2_1 U16905 ( .ip1(rdata[11]), .ip2(n16477), .op(n16480) );
  or2_1 U16906 ( .ip1(n16478), .ip2(n16477), .op(n16479) );
  nand2_1 U16907 ( .ip1(n16480), .ip2(n16479), .op(n16569) );
  inv_1 U16908 ( .ip(n16481), .op(n16578) );
  fulladder U16909 ( .a(n16484), .b(n16483), .ci(n16482), .co(n16577), .s(
        n16451) );
  fulladder U16910 ( .a(n16487), .b(n16486), .ci(n16485), .co(n16576), .s(
        n16444) );
  inv_1 U16911 ( .ip(n16488), .op(n16582) );
  fulladder U16912 ( .a(n16491), .b(n16490), .ci(n16489), .co(n16581), .s(
        n16521) );
  fulladder U16913 ( .a(n16494), .b(n16493), .ci(n16492), .co(n16580), .s(
        n16470) );
  nor2_1 U16914 ( .ip1(n16496), .ip2(n16495), .op(n16556) );
  nand2_1 U16915 ( .ip1(m2DataIn[6]), .ip2(q_w2[14]), .op(n16555) );
  nand2_1 U16916 ( .ip1(m2DataIn[8]), .ip2(q_w2[12]), .op(n16554) );
  nor2_1 U16917 ( .ip1(n16498), .ip2(n16497), .op(n16549) );
  nand2_1 U16918 ( .ip1(m2DataIn[12]), .ip2(q_w2[8]), .op(n16548) );
  nand2_1 U16919 ( .ip1(m2DataIn[7]), .ip2(q_w2[13]), .op(n16547) );
  fulladder U16920 ( .a(n16501), .b(n16500), .ci(n16499), .co(n16557), .s(
        n16519) );
  inv_1 U16921 ( .ip(n16511), .op(n16502) );
  nor2_1 U16922 ( .ip1(n16502), .ip2(n16548), .op(n16504) );
  or2_1 U16923 ( .ip1(n16503), .ip2(n16504), .op(n16507) );
  or2_1 U16924 ( .ip1(n16505), .ip2(n16504), .op(n16506) );
  nand2_1 U16925 ( .ip1(n16507), .ip2(n16506), .op(n16574) );
  nor2_1 U16926 ( .ip1(n16597), .ip2(n16538), .op(n16513) );
  nand2_1 U16927 ( .ip1(q_w2[9]), .ip2(m2DataIn[11]), .op(n16509) );
  nand2_1 U16928 ( .ip1(m2DataIn[13]), .ip2(q_w2[7]), .op(n16508) );
  nand2_1 U16929 ( .ip1(n16509), .ip2(n16508), .op(n16512) );
  nor2_1 U16930 ( .ip1(n16510), .ip2(n16552), .op(n16654) );
  nand2_1 U16931 ( .ip1(n16511), .ip2(n16654), .op(n16536) );
  nand2_1 U16932 ( .ip1(n16512), .ip2(n16536), .op(n16537) );
  xor2_1 U16933 ( .ip1(n16513), .ip2(n16537), .op(n16573) );
  fulladder U16934 ( .a(n16516), .b(n16515), .ci(n16514), .co(n16572), .s(
        n16446) );
  fulladder U16935 ( .a(n16519), .b(n16518), .ci(n16517), .co(n16533), .s(
        n16493) );
  fulladder U16936 ( .a(n16522), .b(n16521), .ci(n16520), .co(n16530), .s(
        n16469) );
  fulladder U16937 ( .a(n16525), .b(n16524), .ci(n16523), .co(n16583), .s(
        n16464) );
  nor2_1 U16938 ( .ip1(n16714), .ip2(n16526), .op(n16527) );
  buf_1 U16939 ( .ip(n16527), .op(n16529) );
  mux2_1 U16940 ( .ip1(n16529), .ip2(\ANSWER/mem[0][0][12] ), .s(n16717), .op(
        n2702) );
  mux2_1 U16941 ( .ip1(n16529), .ip2(\ANSWER/mem[0][1][12] ), .s(n16718), .op(
        n2701) );
  mux2_1 U16942 ( .ip1(n16529), .ip2(\ANSWER/mem[0][2][12] ), .s(n16719), .op(
        n2700) );
  mux2_1 U16943 ( .ip1(n16529), .ip2(\ANSWER/mem[0][3][12] ), .s(n16720), .op(
        n2699) );
  mux2_1 U16944 ( .ip1(n16529), .ip2(\ANSWER/mem[0][4][12] ), .s(n16721), .op(
        n2698) );
  mux2_1 U16945 ( .ip1(n16529), .ip2(\ANSWER/mem[0][5][12] ), .s(n16722), .op(
        n2697) );
  mux2_1 U16946 ( .ip1(n16529), .ip2(\ANSWER/mem[0][6][12] ), .s(n16723), .op(
        n2696) );
  mux2_1 U16947 ( .ip1(n16529), .ip2(\ANSWER/mem[0][7][12] ), .s(n16724), .op(
        n2695) );
  mux2_1 U16948 ( .ip1(n16529), .ip2(\ANSWER/mem[0][8][12] ), .s(n16725), .op(
        n2694) );
  mux2_1 U16949 ( .ip1(n16529), .ip2(\ANSWER/mem[0][9][12] ), .s(n16726), .op(
        n2693) );
  mux2_1 U16950 ( .ip1(n16529), .ip2(\ANSWER/mem[1][0][12] ), .s(n16727), .op(
        n2692) );
  mux2_1 U16951 ( .ip1(n16529), .ip2(\ANSWER/mem[1][1][12] ), .s(n16728), .op(
        n2691) );
  mux2_1 U16952 ( .ip1(n16529), .ip2(\ANSWER/mem[1][2][12] ), .s(n16729), .op(
        n2690) );
  mux2_1 U16953 ( .ip1(n16527), .ip2(\ANSWER/mem[1][3][12] ), .s(n16730), .op(
        n2689) );
  mux2_1 U16954 ( .ip1(n16527), .ip2(\ANSWER/mem[1][4][12] ), .s(n16731), .op(
        n2688) );
  mux2_1 U16955 ( .ip1(n16527), .ip2(\ANSWER/mem[1][5][12] ), .s(n16732), .op(
        n2687) );
  mux2_1 U16956 ( .ip1(n16527), .ip2(\ANSWER/mem[1][6][12] ), .s(n16733), .op(
        n2686) );
  mux2_1 U16957 ( .ip1(n16527), .ip2(\ANSWER/mem[1][7][12] ), .s(n16734), .op(
        n2685) );
  mux2_1 U16958 ( .ip1(n16527), .ip2(\ANSWER/mem[1][8][12] ), .s(n16735), .op(
        n2684) );
  mux2_1 U16959 ( .ip1(n16527), .ip2(\ANSWER/mem[1][9][12] ), .s(n16736), .op(
        n2683) );
  mux2_1 U16960 ( .ip1(n16527), .ip2(\ANSWER/mem[2][0][12] ), .s(n16737), .op(
        n2682) );
  mux2_1 U16961 ( .ip1(n16527), .ip2(\ANSWER/mem[2][1][12] ), .s(n16738), .op(
        n2681) );
  mux2_1 U16962 ( .ip1(n16527), .ip2(\ANSWER/mem[2][2][12] ), .s(n16739), .op(
        n2680) );
  mux2_1 U16963 ( .ip1(n16527), .ip2(\ANSWER/mem[2][3][12] ), .s(n16740), .op(
        n2679) );
  mux2_1 U16964 ( .ip1(n16529), .ip2(\ANSWER/mem[2][4][12] ), .s(n16741), .op(
        n2678) );
  mux2_1 U16965 ( .ip1(n16527), .ip2(\ANSWER/mem[2][5][12] ), .s(n16742), .op(
        n2677) );
  mux2_1 U16966 ( .ip1(n16529), .ip2(\ANSWER/mem[2][6][12] ), .s(n16743), .op(
        n2676) );
  mux2_1 U16967 ( .ip1(n16527), .ip2(\ANSWER/mem[2][7][12] ), .s(n16744), .op(
        n2675) );
  mux2_1 U16968 ( .ip1(n16527), .ip2(\ANSWER/mem[2][8][12] ), .s(n16745), .op(
        n2674) );
  mux2_1 U16969 ( .ip1(n16527), .ip2(\ANSWER/mem[2][9][12] ), .s(n16746), .op(
        n2673) );
  mux2_1 U16970 ( .ip1(n16529), .ip2(\ANSWER/mem[3][0][12] ), .s(n16747), .op(
        n2672) );
  mux2_1 U16971 ( .ip1(n16529), .ip2(\ANSWER/mem[3][1][12] ), .s(n16748), .op(
        n2671) );
  mux2_1 U16972 ( .ip1(n16529), .ip2(\ANSWER/mem[3][2][12] ), .s(n16749), .op(
        n2670) );
  mux2_1 U16973 ( .ip1(n16529), .ip2(\ANSWER/mem[3][3][12] ), .s(n16750), .op(
        n2669) );
  mux2_1 U16974 ( .ip1(n16529), .ip2(\ANSWER/mem[3][4][12] ), .s(n16751), .op(
        n2668) );
  mux2_1 U16975 ( .ip1(n16529), .ip2(\ANSWER/mem[3][5][12] ), .s(n16752), .op(
        n2667) );
  buf_1 U16976 ( .ip(n16527), .op(n16528) );
  mux2_1 U16977 ( .ip1(n16528), .ip2(\ANSWER/mem[3][6][12] ), .s(n16753), .op(
        n2666) );
  mux2_1 U16978 ( .ip1(n16527), .ip2(\ANSWER/mem[3][7][12] ), .s(n16754), .op(
        n2665) );
  mux2_1 U16979 ( .ip1(n16527), .ip2(\ANSWER/mem[3][8][12] ), .s(n16755), .op(
        n2664) );
  mux2_1 U16980 ( .ip1(n16527), .ip2(\ANSWER/mem[3][9][12] ), .s(n16756), .op(
        n2663) );
  mux2_1 U16981 ( .ip1(n16528), .ip2(\ANSWER/mem[4][0][12] ), .s(n16757), .op(
        n2662) );
  mux2_1 U16982 ( .ip1(n16528), .ip2(\ANSWER/mem[4][1][12] ), .s(n16758), .op(
        n2661) );
  mux2_1 U16983 ( .ip1(n16528), .ip2(\ANSWER/mem[4][2][12] ), .s(n16759), .op(
        n2660) );
  mux2_1 U16984 ( .ip1(n16528), .ip2(\ANSWER/mem[4][3][12] ), .s(n16760), .op(
        n2659) );
  mux2_1 U16985 ( .ip1(n16528), .ip2(\ANSWER/mem[4][4][12] ), .s(n16761), .op(
        n2658) );
  mux2_1 U16986 ( .ip1(n16528), .ip2(\ANSWER/mem[4][5][12] ), .s(n16762), .op(
        n2657) );
  mux2_1 U16987 ( .ip1(n16528), .ip2(\ANSWER/mem[4][6][12] ), .s(n16763), .op(
        n2656) );
  mux2_1 U16988 ( .ip1(n16528), .ip2(\ANSWER/mem[4][7][12] ), .s(n16764), .op(
        n2655) );
  mux2_1 U16989 ( .ip1(n16529), .ip2(\ANSWER/mem[4][8][12] ), .s(n16765), .op(
        n2654) );
  mux2_1 U16990 ( .ip1(n16527), .ip2(\ANSWER/mem[4][9][12] ), .s(n16766), .op(
        n2653) );
  mux2_1 U16991 ( .ip1(n16527), .ip2(\ANSWER/mem[5][0][12] ), .s(n16767), .op(
        n2652) );
  mux2_1 U16992 ( .ip1(n16527), .ip2(\ANSWER/mem[5][1][12] ), .s(n16768), .op(
        n2651) );
  mux2_1 U16993 ( .ip1(n16527), .ip2(\ANSWER/mem[5][2][12] ), .s(n16769), .op(
        n2650) );
  mux2_1 U16994 ( .ip1(n16527), .ip2(\ANSWER/mem[5][3][12] ), .s(n16770), .op(
        n2649) );
  mux2_1 U16995 ( .ip1(n16527), .ip2(\ANSWER/mem[5][4][12] ), .s(n16771), .op(
        n2648) );
  mux2_1 U16996 ( .ip1(n16527), .ip2(\ANSWER/mem[5][5][12] ), .s(n16772), .op(
        n2647) );
  mux2_1 U16997 ( .ip1(n16527), .ip2(\ANSWER/mem[5][6][12] ), .s(n16773), .op(
        n2646) );
  mux2_1 U16998 ( .ip1(n16527), .ip2(\ANSWER/mem[5][7][12] ), .s(n16774), .op(
        n2645) );
  mux2_1 U16999 ( .ip1(n16527), .ip2(\ANSWER/mem[5][8][12] ), .s(n16775), .op(
        n2644) );
  mux2_1 U17000 ( .ip1(n16527), .ip2(\ANSWER/mem[5][9][12] ), .s(n16776), .op(
        n2643) );
  mux2_1 U17001 ( .ip1(n16528), .ip2(\ANSWER/mem[6][0][12] ), .s(n16777), .op(
        n2642) );
  mux2_1 U17002 ( .ip1(n16528), .ip2(\ANSWER/mem[6][1][12] ), .s(n16778), .op(
        n2641) );
  mux2_1 U17003 ( .ip1(n16528), .ip2(\ANSWER/mem[6][2][12] ), .s(n16779), .op(
        n2640) );
  mux2_1 U17004 ( .ip1(n16528), .ip2(\ANSWER/mem[6][3][12] ), .s(n16780), .op(
        n2639) );
  mux2_1 U17005 ( .ip1(n16527), .ip2(\ANSWER/mem[6][4][12] ), .s(n16781), .op(
        n2638) );
  mux2_1 U17006 ( .ip1(n16527), .ip2(\ANSWER/mem[6][5][12] ), .s(n16782), .op(
        n2637) );
  mux2_1 U17007 ( .ip1(n16527), .ip2(\ANSWER/mem[6][6][12] ), .s(n16783), .op(
        n2636) );
  mux2_1 U17008 ( .ip1(n16527), .ip2(\ANSWER/mem[6][7][12] ), .s(n16784), .op(
        n2635) );
  mux2_1 U17009 ( .ip1(n16527), .ip2(\ANSWER/mem[6][8][12] ), .s(n16785), .op(
        n2634) );
  mux2_1 U17010 ( .ip1(n16527), .ip2(\ANSWER/mem[6][9][12] ), .s(n16786), .op(
        n2633) );
  mux2_1 U17011 ( .ip1(n16527), .ip2(\ANSWER/mem[7][0][12] ), .s(n16787), .op(
        n2632) );
  mux2_1 U17012 ( .ip1(n16527), .ip2(\ANSWER/mem[7][1][12] ), .s(n16788), .op(
        n2631) );
  mux2_1 U17013 ( .ip1(n16528), .ip2(\ANSWER/mem[7][2][12] ), .s(n16790), .op(
        n2630) );
  mux2_1 U17014 ( .ip1(n16528), .ip2(\ANSWER/mem[7][3][12] ), .s(n16791), .op(
        n2629) );
  mux2_1 U17015 ( .ip1(n16528), .ip2(\ANSWER/mem[7][4][12] ), .s(n16792), .op(
        n2628) );
  mux2_1 U17016 ( .ip1(n16528), .ip2(\ANSWER/mem[7][5][12] ), .s(n16793), .op(
        n2627) );
  mux2_1 U17017 ( .ip1(n16528), .ip2(\ANSWER/mem[7][6][12] ), .s(n16794), .op(
        n2626) );
  mux2_1 U17018 ( .ip1(n16528), .ip2(\ANSWER/mem[7][7][12] ), .s(n16795), .op(
        n2625) );
  mux2_1 U17019 ( .ip1(n16528), .ip2(\ANSWER/mem[7][8][12] ), .s(n16796), .op(
        n2624) );
  mux2_1 U17020 ( .ip1(n16528), .ip2(\ANSWER/mem[7][9][12] ), .s(n16797), .op(
        n2623) );
  mux2_1 U17021 ( .ip1(n16528), .ip2(\ANSWER/mem[8][0][12] ), .s(n16798), .op(
        n2622) );
  mux2_1 U17022 ( .ip1(n16528), .ip2(\ANSWER/mem[8][1][12] ), .s(n16799), .op(
        n2621) );
  mux2_1 U17023 ( .ip1(n16528), .ip2(\ANSWER/mem[8][2][12] ), .s(n16800), .op(
        n2620) );
  mux2_1 U17024 ( .ip1(n16528), .ip2(\ANSWER/mem[8][3][12] ), .s(n16801), .op(
        n2619) );
  mux2_1 U17025 ( .ip1(n16528), .ip2(\ANSWER/mem[8][4][12] ), .s(n16803), .op(
        n2618) );
  mux2_1 U17026 ( .ip1(n16529), .ip2(\ANSWER/mem[8][5][12] ), .s(n16804), .op(
        n2617) );
  mux2_1 U17027 ( .ip1(n16528), .ip2(\ANSWER/mem[8][6][12] ), .s(n16805), .op(
        n2616) );
  mux2_1 U17028 ( .ip1(n16527), .ip2(\ANSWER/mem[8][7][12] ), .s(n16806), .op(
        n2615) );
  mux2_1 U17029 ( .ip1(n16529), .ip2(\ANSWER/mem[8][8][12] ), .s(n16807), .op(
        n2614) );
  mux2_1 U17030 ( .ip1(n16528), .ip2(\ANSWER/mem[8][9][12] ), .s(n16808), .op(
        n2613) );
  mux2_1 U17031 ( .ip1(n16529), .ip2(\ANSWER/mem[9][0][12] ), .s(n16809), .op(
        n2612) );
  mux2_1 U17032 ( .ip1(n16528), .ip2(\ANSWER/mem[9][1][12] ), .s(n16810), .op(
        n2611) );
  mux2_1 U17033 ( .ip1(n16529), .ip2(\ANSWER/mem[9][2][12] ), .s(n16811), .op(
        n2610) );
  mux2_1 U17034 ( .ip1(n16528), .ip2(\ANSWER/mem[9][3][12] ), .s(n16812), .op(
        n2609) );
  mux2_1 U17035 ( .ip1(n16529), .ip2(\ANSWER/mem[9][4][12] ), .s(n16813), .op(
        n2608) );
  mux2_1 U17036 ( .ip1(n16528), .ip2(\ANSWER/mem[9][5][12] ), .s(n16814), .op(
        n2607) );
  mux2_1 U17037 ( .ip1(n16529), .ip2(\ANSWER/mem[9][6][12] ), .s(n16815), .op(
        n2606) );
  mux2_1 U17038 ( .ip1(n16529), .ip2(\ANSWER/mem[9][7][12] ), .s(n16816), .op(
        n2605) );
  mux2_1 U17039 ( .ip1(n16529), .ip2(\ANSWER/mem[9][8][12] ), .s(n16817), .op(
        n2604) );
  mux2_1 U17040 ( .ip1(n16529), .ip2(\ANSWER/mem[9][9][12] ), .s(n16818), .op(
        n2603) );
  fulladder U17041 ( .a(n16532), .b(n16531), .ci(n16530), .co(n16641), .s(
        n16584) );
  fulladder U17042 ( .a(n16535), .b(n16534), .ci(n16533), .co(n16592), .s(
        n16531) );
  inv_1 U17043 ( .ip(n16536), .op(n16540) );
  nor3_1 U17044 ( .ip1(n16597), .ip2(n16538), .ip3(n16537), .op(n16539) );
  nor2_1 U17045 ( .ip1(n16540), .ip2(n16539), .op(n16628) );
  inv_1 U17046 ( .ip(rdata[13]), .op(n16546) );
  nand3_1 U17047 ( .ip1(m2DataIn[11]), .ip2(q_w2[11]), .ip3(n16541), .op(
        n16610) );
  inv_1 U17048 ( .ip(n16610), .op(n16542) );
  or2_1 U17049 ( .ip1(n16677), .ip2(n16542), .op(n16545) );
  nand2_1 U17050 ( .ip1(m2DataIn[11]), .ip2(q_w2[10]), .op(n16543) );
  or2_1 U17051 ( .ip1(n16543), .ip2(n16542), .op(n16544) );
  nand2_1 U17052 ( .ip1(n16545), .ip2(n16544), .op(n16608) );
  mux2_1 U17053 ( .ip1(n16546), .ip2(rdata[13]), .s(n16608), .op(n16627) );
  fulladder U17054 ( .a(n16549), .b(n16548), .ci(n16547), .co(n16626), .s(
        n16558) );
  nor2_1 U17055 ( .ip1(n16690), .ip2(n16678), .op(n16613) );
  nor2_1 U17056 ( .ip1(n16550), .ip2(n16689), .op(n16612) );
  nand2_1 U17057 ( .ip1(m2DataIn[15]), .ip2(q_w2[6]), .op(n16611) );
  inv_1 U17058 ( .ip(n16551), .op(n16617) );
  nor2_1 U17059 ( .ip1(n16623), .ip2(n16552), .op(n16595) );
  nor2_1 U17060 ( .ip1(n16624), .ip2(n16598), .op(n16594) );
  nand2_1 U17061 ( .ip1(m2DataIn[6]), .ip2(q_w2[15]), .op(n16593) );
  inv_1 U17062 ( .ip(n16553), .op(n16616) );
  fulladder U17063 ( .a(n16556), .b(n16555), .ci(n16554), .co(n16615), .s(
        n16559) );
  fulladder U17064 ( .a(n16559), .b(n16558), .ci(n16557), .co(n16636), .s(
        n16535) );
  inv_1 U17065 ( .ip(n16560), .op(n16634) );
  nor2_1 U17066 ( .ip1(n16561), .ip2(n16597), .op(n16563) );
  nand2_1 U17067 ( .ip1(q_w2[8]), .ip2(m2DataIn[13]), .op(n16562) );
  xor2_1 U17068 ( .ip1(n16563), .ip2(n16562), .op(n16618) );
  inv_1 U17069 ( .ip(n16618), .op(n16568) );
  nor2_1 U17070 ( .ip1(n16565), .ip2(n16564), .op(n16566) );
  nor2_1 U17071 ( .ip1(n16567), .ip2(n16566), .op(n16619) );
  mux2_1 U17072 ( .ip1(n16568), .ip2(n16618), .s(n16619), .op(n16631) );
  fulladder U17073 ( .a(n16571), .b(n16570), .ci(n16569), .co(n16630), .s(
        n16481) );
  fulladder U17074 ( .a(n16574), .b(n16573), .ci(n16572), .co(n16629), .s(
        n16534) );
  inv_1 U17075 ( .ip(n16575), .op(n16633) );
  fulladder U17076 ( .a(n16578), .b(n16577), .ci(n16576), .co(n16632), .s(
        n16488) );
  inv_1 U17077 ( .ip(n16579), .op(n16591) );
  fulladder U17078 ( .a(n16582), .b(n16581), .ci(n16580), .co(n16590), .s(
        n16532) );
  fulladder U17079 ( .a(n16585), .b(n16584), .ci(n16583), .co(n16639), .s(
        n16526) );
  nor2_1 U17080 ( .ip1(n16714), .ip2(n16586), .op(n16588) );
  buf_1 U17081 ( .ip(n16588), .op(n16587) );
  mux2_1 U17082 ( .ip1(n16587), .ip2(\ANSWER/mem[0][0][13] ), .s(n16717), .op(
        n2602) );
  mux2_1 U17083 ( .ip1(n16587), .ip2(\ANSWER/mem[0][1][13] ), .s(n16718), .op(
        n2601) );
  mux2_1 U17084 ( .ip1(n16587), .ip2(\ANSWER/mem[0][2][13] ), .s(n16719), .op(
        n2600) );
  mux2_1 U17085 ( .ip1(n16587), .ip2(\ANSWER/mem[0][3][13] ), .s(n16720), .op(
        n2599) );
  mux2_1 U17086 ( .ip1(n16587), .ip2(\ANSWER/mem[0][4][13] ), .s(n16721), .op(
        n2598) );
  mux2_1 U17087 ( .ip1(n16587), .ip2(\ANSWER/mem[0][5][13] ), .s(n16722), .op(
        n2597) );
  mux2_1 U17088 ( .ip1(n16587), .ip2(\ANSWER/mem[0][6][13] ), .s(n16723), .op(
        n2596) );
  mux2_1 U17089 ( .ip1(n16587), .ip2(\ANSWER/mem[0][7][13] ), .s(n16724), .op(
        n2595) );
  mux2_1 U17090 ( .ip1(n16587), .ip2(\ANSWER/mem[0][8][13] ), .s(n16725), .op(
        n2594) );
  mux2_1 U17091 ( .ip1(n16587), .ip2(\ANSWER/mem[0][9][13] ), .s(n16726), .op(
        n2593) );
  mux2_1 U17092 ( .ip1(n16587), .ip2(\ANSWER/mem[1][0][13] ), .s(n16727), .op(
        n2592) );
  mux2_1 U17093 ( .ip1(n16587), .ip2(\ANSWER/mem[1][1][13] ), .s(n16728), .op(
        n2591) );
  mux2_1 U17094 ( .ip1(n16587), .ip2(\ANSWER/mem[1][2][13] ), .s(n16729), .op(
        n2590) );
  mux2_1 U17095 ( .ip1(n16587), .ip2(\ANSWER/mem[1][3][13] ), .s(n16730), .op(
        n2589) );
  mux2_1 U17096 ( .ip1(n16587), .ip2(\ANSWER/mem[1][4][13] ), .s(n16731), .op(
        n2588) );
  mux2_1 U17097 ( .ip1(n16587), .ip2(\ANSWER/mem[1][5][13] ), .s(n16732), .op(
        n2587) );
  mux2_1 U17098 ( .ip1(n16587), .ip2(\ANSWER/mem[1][6][13] ), .s(n16733), .op(
        n2586) );
  mux2_1 U17099 ( .ip1(n16587), .ip2(\ANSWER/mem[1][7][13] ), .s(n16734), .op(
        n2585) );
  mux2_1 U17100 ( .ip1(n16587), .ip2(\ANSWER/mem[1][8][13] ), .s(n16735), .op(
        n2584) );
  mux2_1 U17101 ( .ip1(n16587), .ip2(\ANSWER/mem[1][9][13] ), .s(n16736), .op(
        n2583) );
  mux2_1 U17102 ( .ip1(n16587), .ip2(\ANSWER/mem[2][0][13] ), .s(n16737), .op(
        n2582) );
  mux2_1 U17103 ( .ip1(n16587), .ip2(\ANSWER/mem[2][1][13] ), .s(n16738), .op(
        n2581) );
  mux2_1 U17104 ( .ip1(n16587), .ip2(\ANSWER/mem[2][2][13] ), .s(n16739), .op(
        n2580) );
  mux2_1 U17105 ( .ip1(n16587), .ip2(\ANSWER/mem[2][3][13] ), .s(n16740), .op(
        n2579) );
  mux2_1 U17106 ( .ip1(n16587), .ip2(\ANSWER/mem[2][4][13] ), .s(n16741), .op(
        n2578) );
  mux2_1 U17107 ( .ip1(n16587), .ip2(\ANSWER/mem[2][5][13] ), .s(n16742), .op(
        n2577) );
  mux2_1 U17108 ( .ip1(n16587), .ip2(\ANSWER/mem[2][6][13] ), .s(n16743), .op(
        n2576) );
  mux2_1 U17109 ( .ip1(n16587), .ip2(\ANSWER/mem[2][7][13] ), .s(n16744), .op(
        n2575) );
  mux2_1 U17110 ( .ip1(n16587), .ip2(\ANSWER/mem[2][8][13] ), .s(n16745), .op(
        n2574) );
  mux2_1 U17111 ( .ip1(n16587), .ip2(\ANSWER/mem[2][9][13] ), .s(n16746), .op(
        n2573) );
  mux2_1 U17112 ( .ip1(n16587), .ip2(\ANSWER/mem[3][0][13] ), .s(n16747), .op(
        n2572) );
  mux2_1 U17113 ( .ip1(n16587), .ip2(\ANSWER/mem[3][1][13] ), .s(n16748), .op(
        n2571) );
  mux2_1 U17114 ( .ip1(n16587), .ip2(\ANSWER/mem[3][2][13] ), .s(n16749), .op(
        n2570) );
  mux2_1 U17115 ( .ip1(n16587), .ip2(\ANSWER/mem[3][3][13] ), .s(n16750), .op(
        n2569) );
  mux2_1 U17116 ( .ip1(n16587), .ip2(\ANSWER/mem[3][4][13] ), .s(n16751), .op(
        n2568) );
  mux2_1 U17117 ( .ip1(n16587), .ip2(\ANSWER/mem[3][5][13] ), .s(n16752), .op(
        n2567) );
  mux2_1 U17118 ( .ip1(n16589), .ip2(\ANSWER/mem[3][6][13] ), .s(n16753), .op(
        n2566) );
  mux2_1 U17119 ( .ip1(n16589), .ip2(\ANSWER/mem[3][7][13] ), .s(n16754), .op(
        n2565) );
  mux2_1 U17120 ( .ip1(n16589), .ip2(\ANSWER/mem[3][8][13] ), .s(n16755), .op(
        n2564) );
  mux2_1 U17121 ( .ip1(n16589), .ip2(\ANSWER/mem[3][9][13] ), .s(n16756), .op(
        n2563) );
  mux2_1 U17122 ( .ip1(n16588), .ip2(\ANSWER/mem[4][0][13] ), .s(n16757), .op(
        n2562) );
  mux2_1 U17123 ( .ip1(n16588), .ip2(\ANSWER/mem[4][1][13] ), .s(n16758), .op(
        n2561) );
  mux2_1 U17124 ( .ip1(n16588), .ip2(\ANSWER/mem[4][2][13] ), .s(n16759), .op(
        n2560) );
  mux2_1 U17125 ( .ip1(n16588), .ip2(\ANSWER/mem[4][3][13] ), .s(n16760), .op(
        n2559) );
  mux2_1 U17126 ( .ip1(n16589), .ip2(\ANSWER/mem[4][4][13] ), .s(n16761), .op(
        n2558) );
  mux2_1 U17127 ( .ip1(n16589), .ip2(\ANSWER/mem[4][5][13] ), .s(n16762), .op(
        n2557) );
  mux2_1 U17128 ( .ip1(n16589), .ip2(\ANSWER/mem[4][6][13] ), .s(n16763), .op(
        n2556) );
  mux2_1 U17129 ( .ip1(n16589), .ip2(\ANSWER/mem[4][7][13] ), .s(n16764), .op(
        n2555) );
  mux2_1 U17130 ( .ip1(n16589), .ip2(\ANSWER/mem[4][8][13] ), .s(n16765), .op(
        n2554) );
  mux2_1 U17131 ( .ip1(n16589), .ip2(\ANSWER/mem[4][9][13] ), .s(n16766), .op(
        n2553) );
  mux2_1 U17132 ( .ip1(n16589), .ip2(\ANSWER/mem[5][0][13] ), .s(n16767), .op(
        n2552) );
  mux2_1 U17133 ( .ip1(n16588), .ip2(\ANSWER/mem[5][1][13] ), .s(n16768), .op(
        n2551) );
  mux2_1 U17134 ( .ip1(n16589), .ip2(\ANSWER/mem[5][2][13] ), .s(n16769), .op(
        n2550) );
  mux2_1 U17135 ( .ip1(n16588), .ip2(\ANSWER/mem[5][3][13] ), .s(n16770), .op(
        n2549) );
  mux2_1 U17136 ( .ip1(n16589), .ip2(\ANSWER/mem[5][4][13] ), .s(n16771), .op(
        n2548) );
  mux2_1 U17137 ( .ip1(n16588), .ip2(\ANSWER/mem[5][5][13] ), .s(n16772), .op(
        n2547) );
  mux2_1 U17138 ( .ip1(n16588), .ip2(\ANSWER/mem[5][6][13] ), .s(n16773), .op(
        n2546) );
  mux2_1 U17139 ( .ip1(n16588), .ip2(\ANSWER/mem[5][7][13] ), .s(n16774), .op(
        n2545) );
  mux2_1 U17140 ( .ip1(n16588), .ip2(\ANSWER/mem[5][8][13] ), .s(n16775), .op(
        n2544) );
  mux2_1 U17141 ( .ip1(n16588), .ip2(\ANSWER/mem[5][9][13] ), .s(n16776), .op(
        n2543) );
  mux2_1 U17142 ( .ip1(n16588), .ip2(\ANSWER/mem[6][0][13] ), .s(n16777), .op(
        n2542) );
  mux2_1 U17143 ( .ip1(n16588), .ip2(\ANSWER/mem[6][1][13] ), .s(n16778), .op(
        n2541) );
  mux2_1 U17144 ( .ip1(n16588), .ip2(\ANSWER/mem[6][2][13] ), .s(n16779), .op(
        n2540) );
  mux2_1 U17145 ( .ip1(n16588), .ip2(\ANSWER/mem[6][3][13] ), .s(n16780), .op(
        n2539) );
  mux2_1 U17146 ( .ip1(n16588), .ip2(\ANSWER/mem[6][4][13] ), .s(n16781), .op(
        n2538) );
  mux2_1 U17147 ( .ip1(n16588), .ip2(\ANSWER/mem[6][5][13] ), .s(n16782), .op(
        n2537) );
  mux2_1 U17148 ( .ip1(n16588), .ip2(\ANSWER/mem[6][6][13] ), .s(n16783), .op(
        n2536) );
  mux2_1 U17149 ( .ip1(n16588), .ip2(\ANSWER/mem[6][7][13] ), .s(n16784), .op(
        n2535) );
  mux2_1 U17150 ( .ip1(n16588), .ip2(\ANSWER/mem[6][8][13] ), .s(n16785), .op(
        n2534) );
  mux2_1 U17151 ( .ip1(n16588), .ip2(\ANSWER/mem[6][9][13] ), .s(n16786), .op(
        n2533) );
  mux2_1 U17152 ( .ip1(n16588), .ip2(\ANSWER/mem[7][0][13] ), .s(n16787), .op(
        n2532) );
  mux2_1 U17153 ( .ip1(n16588), .ip2(\ANSWER/mem[7][1][13] ), .s(n16788), .op(
        n2531) );
  buf_1 U17154 ( .ip(n16588), .op(n16589) );
  mux2_1 U17155 ( .ip1(n16589), .ip2(\ANSWER/mem[7][2][13] ), .s(n16790), .op(
        n2530) );
  mux2_1 U17156 ( .ip1(n16589), .ip2(\ANSWER/mem[7][3][13] ), .s(n16791), .op(
        n2529) );
  mux2_1 U17157 ( .ip1(n16589), .ip2(\ANSWER/mem[7][4][13] ), .s(n16792), .op(
        n2528) );
  mux2_1 U17158 ( .ip1(n16588), .ip2(\ANSWER/mem[7][5][13] ), .s(n16793), .op(
        n2527) );
  mux2_1 U17159 ( .ip1(n16588), .ip2(\ANSWER/mem[7][6][13] ), .s(n16794), .op(
        n2526) );
  mux2_1 U17160 ( .ip1(n16589), .ip2(\ANSWER/mem[7][7][13] ), .s(n16795), .op(
        n2525) );
  mux2_1 U17161 ( .ip1(n16589), .ip2(\ANSWER/mem[7][8][13] ), .s(n16796), .op(
        n2524) );
  mux2_1 U17162 ( .ip1(n16589), .ip2(\ANSWER/mem[7][9][13] ), .s(n16797), .op(
        n2523) );
  mux2_1 U17163 ( .ip1(n16589), .ip2(\ANSWER/mem[8][0][13] ), .s(n16798), .op(
        n2522) );
  mux2_1 U17164 ( .ip1(n16589), .ip2(\ANSWER/mem[8][1][13] ), .s(n16799), .op(
        n2521) );
  mux2_1 U17165 ( .ip1(n16589), .ip2(\ANSWER/mem[8][2][13] ), .s(n16800), .op(
        n2520) );
  mux2_1 U17166 ( .ip1(n16589), .ip2(\ANSWER/mem[8][3][13] ), .s(n16801), .op(
        n2519) );
  mux2_1 U17167 ( .ip1(n16588), .ip2(\ANSWER/mem[8][4][13] ), .s(n16803), .op(
        n2518) );
  mux2_1 U17168 ( .ip1(n16588), .ip2(\ANSWER/mem[8][5][13] ), .s(n16804), .op(
        n2517) );
  mux2_1 U17169 ( .ip1(n16588), .ip2(\ANSWER/mem[8][6][13] ), .s(n16805), .op(
        n2516) );
  mux2_1 U17170 ( .ip1(n16588), .ip2(\ANSWER/mem[8][7][13] ), .s(n16806), .op(
        n2515) );
  mux2_1 U17171 ( .ip1(n16588), .ip2(\ANSWER/mem[8][8][13] ), .s(n16807), .op(
        n2514) );
  mux2_1 U17172 ( .ip1(n16588), .ip2(\ANSWER/mem[8][9][13] ), .s(n16808), .op(
        n2513) );
  mux2_1 U17173 ( .ip1(n16588), .ip2(\ANSWER/mem[9][0][13] ), .s(n16809), .op(
        n2512) );
  mux2_1 U17174 ( .ip1(n16588), .ip2(\ANSWER/mem[9][1][13] ), .s(n16810), .op(
        n2511) );
  mux2_1 U17175 ( .ip1(n16588), .ip2(\ANSWER/mem[9][2][13] ), .s(n16811), .op(
        n2510) );
  mux2_1 U17176 ( .ip1(n16588), .ip2(\ANSWER/mem[9][3][13] ), .s(n16812), .op(
        n2509) );
  mux2_1 U17177 ( .ip1(n16588), .ip2(\ANSWER/mem[9][4][13] ), .s(n16813), .op(
        n2508) );
  mux2_1 U17178 ( .ip1(n16588), .ip2(\ANSWER/mem[9][5][13] ), .s(n16814), .op(
        n2507) );
  mux2_1 U17179 ( .ip1(n16589), .ip2(\ANSWER/mem[9][6][13] ), .s(n16815), .op(
        n2506) );
  mux2_1 U17180 ( .ip1(n16589), .ip2(\ANSWER/mem[9][7][13] ), .s(n16816), .op(
        n2505) );
  mux2_1 U17181 ( .ip1(n16589), .ip2(\ANSWER/mem[9][8][13] ), .s(n16817), .op(
        n2504) );
  mux2_1 U17182 ( .ip1(n16589), .ip2(\ANSWER/mem[9][9][13] ), .s(n16818), .op(
        n2503) );
  fulladder U17183 ( .a(n16592), .b(n16591), .ci(n16590), .co(n16696), .s(
        n16640) );
  fulladder U17184 ( .a(n16595), .b(n16594), .ci(n16593), .co(n16693), .s(
        n16553) );
  nor2_1 U17185 ( .ip1(n16597), .ip2(n16596), .op(n16662) );
  nor2_1 U17186 ( .ip1(n16690), .ip2(n16598), .op(n16661) );
  nand2_1 U17187 ( .ip1(m2DataIn[7]), .ip2(q_w2[15]), .op(n16660) );
  inv_1 U17188 ( .ip(rdata[14]), .op(n16606) );
  nand2_1 U17189 ( .ip1(m2DataIn[11]), .ip2(q_w2[11]), .op(n16601) );
  nor4_1 U17190 ( .ip1(n16679), .ip2(n16600), .ip3(n16599), .ip4(n16678), .op(
        n16602) );
  or2_1 U17191 ( .ip1(n16601), .ip2(n16602), .op(n16605) );
  nand2_1 U17192 ( .ip1(m2DataIn[10]), .ip2(q_w2[12]), .op(n16603) );
  or2_1 U17193 ( .ip1(n16603), .ip2(n16602), .op(n16604) );
  nand2_1 U17194 ( .ip1(n16605), .ip2(n16604), .op(n16676) );
  mux2_1 U17195 ( .ip1(rdata[14]), .ip2(n16606), .s(n16676), .op(n16691) );
  inv_1 U17196 ( .ip(n16607), .op(n16657) );
  nand2_1 U17197 ( .ip1(rdata[13]), .ip2(n16608), .op(n16609) );
  nand2_1 U17198 ( .ip1(n16610), .ip2(n16609), .op(n16653) );
  fulladder U17199 ( .a(n16613), .b(n16612), .ci(n16611), .co(n16652), .s(
        n16551) );
  inv_1 U17200 ( .ip(n16614), .op(n16656) );
  fulladder U17201 ( .a(n16617), .b(n16616), .ci(n16615), .co(n16655), .s(
        n16637) );
  and3_1 U17202 ( .ip1(m2DataIn[13]), .ip2(q_w2[7]), .ip3(n16662), .op(n16621)
         );
  nor2_1 U17203 ( .ip1(n16619), .ip2(n16618), .op(n16620) );
  nor2_1 U17204 ( .ip1(n16621), .ip2(n16620), .op(n16668) );
  nor2_1 U17205 ( .ip1(n16623), .ip2(n16622), .op(n16671) );
  nor2_1 U17206 ( .ip1(n16624), .ip2(n16689), .op(n16670) );
  nand2_1 U17207 ( .ip1(m2DataIn[15]), .ip2(q_w2[7]), .op(n16669) );
  inv_1 U17208 ( .ip(n16625), .op(n16667) );
  fulladder U17209 ( .a(n16628), .b(n16627), .ci(n16626), .co(n16666), .s(
        n16638) );
  fulladder U17210 ( .a(n16631), .b(n16630), .ci(n16629), .co(n16699), .s(
        n16575) );
  fulladder U17211 ( .a(n16634), .b(n16633), .ci(n16632), .co(n16635), .s(
        n16579) );
  inv_1 U17212 ( .ip(n16635), .op(n16703) );
  fulladder U17213 ( .a(n16638), .b(n16637), .ci(n16636), .co(n16702), .s(
        n16560) );
  fulladder U17214 ( .a(n16641), .b(n16640), .ci(n16639), .co(n16694), .s(
        n16586) );
  nor2_1 U17215 ( .ip1(n16714), .ip2(n16642), .op(n16644) );
  buf_1 U17216 ( .ip(n16644), .op(n16643) );
  mux2_1 U17217 ( .ip1(n16643), .ip2(\ANSWER/mem[0][0][14] ), .s(n16717), .op(
        n2502) );
  mux2_1 U17218 ( .ip1(n16643), .ip2(\ANSWER/mem[0][1][14] ), .s(n16718), .op(
        n2501) );
  mux2_1 U17219 ( .ip1(n16643), .ip2(\ANSWER/mem[0][2][14] ), .s(n16719), .op(
        n2500) );
  mux2_1 U17220 ( .ip1(n16643), .ip2(\ANSWER/mem[0][3][14] ), .s(n16720), .op(
        n2499) );
  mux2_1 U17221 ( .ip1(n16643), .ip2(\ANSWER/mem[0][4][14] ), .s(n16721), .op(
        n2498) );
  mux2_1 U17222 ( .ip1(n16643), .ip2(\ANSWER/mem[0][5][14] ), .s(n16722), .op(
        n2497) );
  mux2_1 U17223 ( .ip1(n16643), .ip2(\ANSWER/mem[0][6][14] ), .s(n16723), .op(
        n2496) );
  mux2_1 U17224 ( .ip1(n16643), .ip2(\ANSWER/mem[0][7][14] ), .s(n16724), .op(
        n2495) );
  mux2_1 U17225 ( .ip1(n16643), .ip2(\ANSWER/mem[0][8][14] ), .s(n16725), .op(
        n2494) );
  mux2_1 U17226 ( .ip1(n16643), .ip2(\ANSWER/mem[0][9][14] ), .s(n16726), .op(
        n2493) );
  mux2_1 U17227 ( .ip1(n16643), .ip2(\ANSWER/mem[1][0][14] ), .s(n16727), .op(
        n2492) );
  mux2_1 U17228 ( .ip1(n16643), .ip2(\ANSWER/mem[1][1][14] ), .s(n16728), .op(
        n2491) );
  mux2_1 U17229 ( .ip1(n16643), .ip2(\ANSWER/mem[1][2][14] ), .s(n16729), .op(
        n2490) );
  mux2_1 U17230 ( .ip1(n16643), .ip2(\ANSWER/mem[1][3][14] ), .s(n16730), .op(
        n2489) );
  mux2_1 U17231 ( .ip1(n16643), .ip2(\ANSWER/mem[1][4][14] ), .s(n16731), .op(
        n2488) );
  mux2_1 U17232 ( .ip1(n16643), .ip2(\ANSWER/mem[1][5][14] ), .s(n16732), .op(
        n2487) );
  mux2_1 U17233 ( .ip1(n16643), .ip2(\ANSWER/mem[1][6][14] ), .s(n16733), .op(
        n2486) );
  mux2_1 U17234 ( .ip1(n16643), .ip2(\ANSWER/mem[1][7][14] ), .s(n16734), .op(
        n2485) );
  mux2_1 U17235 ( .ip1(n16643), .ip2(\ANSWER/mem[1][8][14] ), .s(n16735), .op(
        n2484) );
  mux2_1 U17236 ( .ip1(n16643), .ip2(\ANSWER/mem[1][9][14] ), .s(n16736), .op(
        n2483) );
  mux2_1 U17237 ( .ip1(n16643), .ip2(\ANSWER/mem[2][0][14] ), .s(n16737), .op(
        n2482) );
  mux2_1 U17238 ( .ip1(n16643), .ip2(\ANSWER/mem[2][1][14] ), .s(n16738), .op(
        n2481) );
  mux2_1 U17239 ( .ip1(n16643), .ip2(\ANSWER/mem[2][2][14] ), .s(n16739), .op(
        n2480) );
  mux2_1 U17240 ( .ip1(n16643), .ip2(\ANSWER/mem[2][3][14] ), .s(n16740), .op(
        n2479) );
  mux2_1 U17241 ( .ip1(n16643), .ip2(\ANSWER/mem[2][4][14] ), .s(n16741), .op(
        n2478) );
  mux2_1 U17242 ( .ip1(n16643), .ip2(\ANSWER/mem[2][5][14] ), .s(n16742), .op(
        n2477) );
  mux2_1 U17243 ( .ip1(n16643), .ip2(\ANSWER/mem[2][6][14] ), .s(n16743), .op(
        n2476) );
  mux2_1 U17244 ( .ip1(n16643), .ip2(\ANSWER/mem[2][7][14] ), .s(n16744), .op(
        n2475) );
  mux2_1 U17245 ( .ip1(n16643), .ip2(\ANSWER/mem[2][8][14] ), .s(n16745), .op(
        n2474) );
  mux2_1 U17246 ( .ip1(n16643), .ip2(\ANSWER/mem[2][9][14] ), .s(n16746), .op(
        n2473) );
  mux2_1 U17247 ( .ip1(n16643), .ip2(\ANSWER/mem[3][0][14] ), .s(n16747), .op(
        n2472) );
  mux2_1 U17248 ( .ip1(n16643), .ip2(\ANSWER/mem[3][1][14] ), .s(n16748), .op(
        n2471) );
  mux2_1 U17249 ( .ip1(n16643), .ip2(\ANSWER/mem[3][2][14] ), .s(n16749), .op(
        n2470) );
  mux2_1 U17250 ( .ip1(n16643), .ip2(\ANSWER/mem[3][3][14] ), .s(n16750), .op(
        n2469) );
  mux2_1 U17251 ( .ip1(n16643), .ip2(\ANSWER/mem[3][4][14] ), .s(n16751), .op(
        n2468) );
  mux2_1 U17252 ( .ip1(n16643), .ip2(\ANSWER/mem[3][5][14] ), .s(n16752), .op(
        n2467) );
  mux2_1 U17253 ( .ip1(n16645), .ip2(\ANSWER/mem[3][6][14] ), .s(n16753), .op(
        n2466) );
  mux2_1 U17254 ( .ip1(n16645), .ip2(\ANSWER/mem[3][7][14] ), .s(n16754), .op(
        n2465) );
  mux2_1 U17255 ( .ip1(n16645), .ip2(\ANSWER/mem[3][8][14] ), .s(n16755), .op(
        n2464) );
  mux2_1 U17256 ( .ip1(n16645), .ip2(\ANSWER/mem[3][9][14] ), .s(n16756), .op(
        n2463) );
  mux2_1 U17257 ( .ip1(n16644), .ip2(\ANSWER/mem[4][0][14] ), .s(n16757), .op(
        n2462) );
  mux2_1 U17258 ( .ip1(n16644), .ip2(\ANSWER/mem[4][1][14] ), .s(n16758), .op(
        n2461) );
  mux2_1 U17259 ( .ip1(n16644), .ip2(\ANSWER/mem[4][2][14] ), .s(n16759), .op(
        n2460) );
  mux2_1 U17260 ( .ip1(n16644), .ip2(\ANSWER/mem[4][3][14] ), .s(n16760), .op(
        n2459) );
  mux2_1 U17261 ( .ip1(n16645), .ip2(\ANSWER/mem[4][4][14] ), .s(n16761), .op(
        n2458) );
  mux2_1 U17262 ( .ip1(n16645), .ip2(\ANSWER/mem[4][5][14] ), .s(n16762), .op(
        n2457) );
  mux2_1 U17263 ( .ip1(n16645), .ip2(\ANSWER/mem[4][6][14] ), .s(n16763), .op(
        n2456) );
  mux2_1 U17264 ( .ip1(n16645), .ip2(\ANSWER/mem[4][7][14] ), .s(n16764), .op(
        n2455) );
  mux2_1 U17265 ( .ip1(n16645), .ip2(\ANSWER/mem[4][8][14] ), .s(n16765), .op(
        n2454) );
  mux2_1 U17266 ( .ip1(n16645), .ip2(\ANSWER/mem[4][9][14] ), .s(n16766), .op(
        n2453) );
  mux2_1 U17267 ( .ip1(n16645), .ip2(\ANSWER/mem[5][0][14] ), .s(n16767), .op(
        n2452) );
  mux2_1 U17268 ( .ip1(n16644), .ip2(\ANSWER/mem[5][1][14] ), .s(n16768), .op(
        n2451) );
  mux2_1 U17269 ( .ip1(n16645), .ip2(\ANSWER/mem[5][2][14] ), .s(n16769), .op(
        n2450) );
  mux2_1 U17270 ( .ip1(n16644), .ip2(\ANSWER/mem[5][3][14] ), .s(n16770), .op(
        n2449) );
  mux2_1 U17271 ( .ip1(n16645), .ip2(\ANSWER/mem[5][4][14] ), .s(n16771), .op(
        n2448) );
  mux2_1 U17272 ( .ip1(n16644), .ip2(\ANSWER/mem[5][5][14] ), .s(n16772), .op(
        n2447) );
  mux2_1 U17273 ( .ip1(n16644), .ip2(\ANSWER/mem[5][6][14] ), .s(n16773), .op(
        n2446) );
  mux2_1 U17274 ( .ip1(n16644), .ip2(\ANSWER/mem[5][7][14] ), .s(n16774), .op(
        n2445) );
  mux2_1 U17275 ( .ip1(n16644), .ip2(\ANSWER/mem[5][8][14] ), .s(n16775), .op(
        n2444) );
  mux2_1 U17276 ( .ip1(n16644), .ip2(\ANSWER/mem[5][9][14] ), .s(n16776), .op(
        n2443) );
  mux2_1 U17277 ( .ip1(n16644), .ip2(\ANSWER/mem[6][0][14] ), .s(n16777), .op(
        n2442) );
  mux2_1 U17278 ( .ip1(n16644), .ip2(\ANSWER/mem[6][1][14] ), .s(n16778), .op(
        n2441) );
  mux2_1 U17279 ( .ip1(n16644), .ip2(\ANSWER/mem[6][2][14] ), .s(n16779), .op(
        n2440) );
  mux2_1 U17280 ( .ip1(n16644), .ip2(\ANSWER/mem[6][3][14] ), .s(n16780), .op(
        n2439) );
  mux2_1 U17281 ( .ip1(n16644), .ip2(\ANSWER/mem[6][4][14] ), .s(n16781), .op(
        n2438) );
  mux2_1 U17282 ( .ip1(n16644), .ip2(\ANSWER/mem[6][5][14] ), .s(n16782), .op(
        n2437) );
  mux2_1 U17283 ( .ip1(n16644), .ip2(\ANSWER/mem[6][6][14] ), .s(n16783), .op(
        n2436) );
  mux2_1 U17284 ( .ip1(n16644), .ip2(\ANSWER/mem[6][7][14] ), .s(n16784), .op(
        n2435) );
  mux2_1 U17285 ( .ip1(n16644), .ip2(\ANSWER/mem[6][8][14] ), .s(n16785), .op(
        n2434) );
  mux2_1 U17286 ( .ip1(n16644), .ip2(\ANSWER/mem[6][9][14] ), .s(n16786), .op(
        n2433) );
  mux2_1 U17287 ( .ip1(n16644), .ip2(\ANSWER/mem[7][0][14] ), .s(n16787), .op(
        n2432) );
  mux2_1 U17288 ( .ip1(n16644), .ip2(\ANSWER/mem[7][1][14] ), .s(n16788), .op(
        n2431) );
  buf_1 U17289 ( .ip(n16644), .op(n16645) );
  mux2_1 U17290 ( .ip1(n16645), .ip2(\ANSWER/mem[7][2][14] ), .s(n16790), .op(
        n2430) );
  mux2_1 U17291 ( .ip1(n16645), .ip2(\ANSWER/mem[7][3][14] ), .s(n16791), .op(
        n2429) );
  mux2_1 U17292 ( .ip1(n16645), .ip2(\ANSWER/mem[7][4][14] ), .s(n16792), .op(
        n2428) );
  mux2_1 U17293 ( .ip1(n16644), .ip2(\ANSWER/mem[7][5][14] ), .s(n16793), .op(
        n2427) );
  mux2_1 U17294 ( .ip1(n16644), .ip2(\ANSWER/mem[7][6][14] ), .s(n16794), .op(
        n2426) );
  mux2_1 U17295 ( .ip1(n16645), .ip2(\ANSWER/mem[7][7][14] ), .s(n16795), .op(
        n2425) );
  mux2_1 U17296 ( .ip1(n16645), .ip2(\ANSWER/mem[7][8][14] ), .s(n16796), .op(
        n2424) );
  mux2_1 U17297 ( .ip1(n16645), .ip2(\ANSWER/mem[7][9][14] ), .s(n16797), .op(
        n2423) );
  mux2_1 U17298 ( .ip1(n16645), .ip2(\ANSWER/mem[8][0][14] ), .s(n16798), .op(
        n2422) );
  mux2_1 U17299 ( .ip1(n16645), .ip2(\ANSWER/mem[8][1][14] ), .s(n16799), .op(
        n2421) );
  mux2_1 U17300 ( .ip1(n16645), .ip2(\ANSWER/mem[8][2][14] ), .s(n16800), .op(
        n2420) );
  mux2_1 U17301 ( .ip1(n16645), .ip2(\ANSWER/mem[8][3][14] ), .s(n16801), .op(
        n2419) );
  mux2_1 U17302 ( .ip1(n16644), .ip2(\ANSWER/mem[8][4][14] ), .s(n16803), .op(
        n2418) );
  mux2_1 U17303 ( .ip1(n16644), .ip2(\ANSWER/mem[8][5][14] ), .s(n16804), .op(
        n2417) );
  mux2_1 U17304 ( .ip1(n16644), .ip2(\ANSWER/mem[8][6][14] ), .s(n16805), .op(
        n2416) );
  mux2_1 U17305 ( .ip1(n16644), .ip2(\ANSWER/mem[8][7][14] ), .s(n16806), .op(
        n2415) );
  mux2_1 U17306 ( .ip1(n16644), .ip2(\ANSWER/mem[8][8][14] ), .s(n16807), .op(
        n2414) );
  mux2_1 U17307 ( .ip1(n16644), .ip2(\ANSWER/mem[8][9][14] ), .s(n16808), .op(
        n2413) );
  mux2_1 U17308 ( .ip1(n16644), .ip2(\ANSWER/mem[9][0][14] ), .s(n16809), .op(
        n2412) );
  mux2_1 U17309 ( .ip1(n16644), .ip2(\ANSWER/mem[9][1][14] ), .s(n16810), .op(
        n2411) );
  mux2_1 U17310 ( .ip1(n16644), .ip2(\ANSWER/mem[9][2][14] ), .s(n16811), .op(
        n2410) );
  mux2_1 U17311 ( .ip1(n16644), .ip2(\ANSWER/mem[9][3][14] ), .s(n16812), .op(
        n2409) );
  mux2_1 U17312 ( .ip1(n16644), .ip2(\ANSWER/mem[9][4][14] ), .s(n16813), .op(
        n2408) );
  mux2_1 U17313 ( .ip1(n16644), .ip2(\ANSWER/mem[9][5][14] ), .s(n16814), .op(
        n2407) );
  mux2_1 U17314 ( .ip1(n16645), .ip2(\ANSWER/mem[9][6][14] ), .s(n16815), .op(
        n2406) );
  mux2_1 U17315 ( .ip1(n16645), .ip2(\ANSWER/mem[9][7][14] ), .s(n16816), .op(
        n2405) );
  mux2_1 U17316 ( .ip1(n16645), .ip2(\ANSWER/mem[9][8][14] ), .s(n16817), .op(
        n2404) );
  mux2_1 U17317 ( .ip1(n16645), .ip2(\ANSWER/mem[9][9][14] ), .s(n16818), .op(
        n2403) );
  nand2_1 U17318 ( .ip1(q_w2[15]), .ip2(m2DataIn[8]), .op(n16647) );
  nand2_1 U17319 ( .ip1(q_w2[10]), .ip2(m2DataIn[13]), .op(n16646) );
  xor2_1 U17320 ( .ip1(n16647), .ip2(n16646), .op(n16651) );
  nand2_1 U17321 ( .ip1(q_w2[11]), .ip2(m2DataIn[12]), .op(n16649) );
  nand2_1 U17322 ( .ip1(q_w2[9]), .ip2(m2DataIn[14]), .op(n16648) );
  xor2_1 U17323 ( .ip1(n16649), .ip2(n16648), .op(n16650) );
  xor2_1 U17324 ( .ip1(n16651), .ip2(n16650), .op(n16716) );
  fulladder U17325 ( .a(n16654), .b(n16653), .ci(n16652), .co(n16659), .s(
        n16614) );
  fulladder U17326 ( .a(n16657), .b(n16656), .ci(n16655), .co(n16658), .s(
        n16701) );
  xor2_1 U17327 ( .ip1(n16659), .ip2(n16658), .op(n16665) );
  fulladder U17328 ( .a(n16662), .b(n16661), .ci(n16660), .co(n16663), .s(
        n16692) );
  xor2_1 U17329 ( .ip1(rdata[15]), .ip2(n16663), .op(n16664) );
  xor2_1 U17330 ( .ip1(n16665), .ip2(n16664), .op(n16675) );
  fulladder U17331 ( .a(n16668), .b(n16667), .ci(n16666), .co(n16673), .s(
        n16700) );
  fulladder U17332 ( .a(n16671), .b(n16670), .ci(n16669), .co(n16672), .s(
        n16625) );
  xor2_1 U17333 ( .ip1(n16673), .ip2(n16672), .op(n16674) );
  xor2_1 U17334 ( .ip1(n16675), .ip2(n16674), .op(n16684) );
  nand2_1 U17335 ( .ip1(rdata[14]), .ip2(n16676), .op(n16682) );
  nand2_1 U17336 ( .ip1(n16677), .ip2(n16682), .op(n16681) );
  nor2_1 U17337 ( .ip1(n16679), .ip2(n16678), .op(n16680) );
  mux2_1 U17338 ( .ip1(n16682), .ip2(n16681), .s(n16680), .op(n16683) );
  xor2_1 U17339 ( .ip1(n16684), .ip2(n16683), .op(n16688) );
  nand2_1 U17340 ( .ip1(q_w2[13]), .ip2(m2DataIn[10]), .op(n16686) );
  nand2_1 U17341 ( .ip1(q_w2[8]), .ip2(m2DataIn[15]), .op(n16685) );
  xor2_1 U17342 ( .ip1(n16686), .ip2(n16685), .op(n16687) );
  xor2_1 U17343 ( .ip1(n16688), .ip2(n16687), .op(n16712) );
  nor2_1 U17344 ( .ip1(n16690), .ip2(n16689), .op(n16710) );
  fulladder U17345 ( .a(n16693), .b(n16692), .ci(n16691), .co(n16698), .s(
        n16607) );
  fulladder U17346 ( .a(n16696), .b(n16695), .ci(n16694), .co(n16697), .s(
        n16642) );
  xor2_1 U17347 ( .ip1(n16698), .ip2(n16697), .op(n16708) );
  fulladder U17348 ( .a(n16701), .b(n16700), .ci(n16699), .co(n16706), .s(
        n16704) );
  fulladder U17349 ( .a(n16704), .b(n16703), .ci(n16702), .co(n16705), .s(
        n16695) );
  xor2_1 U17350 ( .ip1(n16706), .ip2(n16705), .op(n16707) );
  xor2_1 U17351 ( .ip1(n16708), .ip2(n16707), .op(n16709) );
  xor2_1 U17352 ( .ip1(n16710), .ip2(n16709), .op(n16711) );
  xor2_1 U17353 ( .ip1(n16712), .ip2(n16711), .op(n16715) );
  nor2_1 U17354 ( .ip1(n16716), .ip2(n16715), .op(n16713) );
  not_ab_or_c_or_d U17355 ( .ip1(n16716), .ip2(n16715), .ip3(n16714), .ip4(
        n16713), .op(n16789) );
  buf_1 U17356 ( .ip(n16789), .op(n16819) );
  mux2_1 U17357 ( .ip1(n16819), .ip2(\ANSWER/mem[0][0][15] ), .s(n16717), .op(
        n2402) );
  mux2_1 U17358 ( .ip1(n16819), .ip2(\ANSWER/mem[0][1][15] ), .s(n16718), .op(
        n2401) );
  mux2_1 U17359 ( .ip1(n16819), .ip2(\ANSWER/mem[0][2][15] ), .s(n16719), .op(
        n2400) );
  mux2_1 U17360 ( .ip1(n16819), .ip2(\ANSWER/mem[0][3][15] ), .s(n16720), .op(
        n2399) );
  mux2_1 U17361 ( .ip1(n16819), .ip2(\ANSWER/mem[0][4][15] ), .s(n16721), .op(
        n2398) );
  mux2_1 U17362 ( .ip1(n16819), .ip2(\ANSWER/mem[0][5][15] ), .s(n16722), .op(
        n2397) );
  mux2_1 U17363 ( .ip1(n16819), .ip2(\ANSWER/mem[0][6][15] ), .s(n16723), .op(
        n2396) );
  mux2_1 U17364 ( .ip1(n16819), .ip2(\ANSWER/mem[0][7][15] ), .s(n16724), .op(
        n2395) );
  mux2_1 U17365 ( .ip1(n16819), .ip2(\ANSWER/mem[0][8][15] ), .s(n16725), .op(
        n2394) );
  mux2_1 U17366 ( .ip1(n16819), .ip2(\ANSWER/mem[0][9][15] ), .s(n16726), .op(
        n2393) );
  mux2_1 U17367 ( .ip1(n16819), .ip2(\ANSWER/mem[1][0][15] ), .s(n16727), .op(
        n2392) );
  mux2_1 U17368 ( .ip1(n16819), .ip2(\ANSWER/mem[1][1][15] ), .s(n16728), .op(
        n2391) );
  mux2_1 U17369 ( .ip1(n16819), .ip2(\ANSWER/mem[1][2][15] ), .s(n16729), .op(
        n2390) );
  mux2_1 U17370 ( .ip1(n16789), .ip2(\ANSWER/mem[1][3][15] ), .s(n16730), .op(
        n2389) );
  mux2_1 U17371 ( .ip1(n16789), .ip2(\ANSWER/mem[1][4][15] ), .s(n16731), .op(
        n2388) );
  mux2_1 U17372 ( .ip1(n16789), .ip2(\ANSWER/mem[1][5][15] ), .s(n16732), .op(
        n2387) );
  mux2_1 U17373 ( .ip1(n16789), .ip2(\ANSWER/mem[1][6][15] ), .s(n16733), .op(
        n2386) );
  mux2_1 U17374 ( .ip1(n16789), .ip2(\ANSWER/mem[1][7][15] ), .s(n16734), .op(
        n2385) );
  mux2_1 U17375 ( .ip1(n16789), .ip2(\ANSWER/mem[1][8][15] ), .s(n16735), .op(
        n2384) );
  mux2_1 U17376 ( .ip1(n16789), .ip2(\ANSWER/mem[1][9][15] ), .s(n16736), .op(
        n2383) );
  mux2_1 U17377 ( .ip1(n16789), .ip2(\ANSWER/mem[2][0][15] ), .s(n16737), .op(
        n2382) );
  mux2_1 U17378 ( .ip1(n16789), .ip2(\ANSWER/mem[2][1][15] ), .s(n16738), .op(
        n2381) );
  mux2_1 U17379 ( .ip1(n16789), .ip2(\ANSWER/mem[2][2][15] ), .s(n16739), .op(
        n2380) );
  mux2_1 U17380 ( .ip1(n16789), .ip2(\ANSWER/mem[2][3][15] ), .s(n16740), .op(
        n2379) );
  mux2_1 U17381 ( .ip1(n16819), .ip2(\ANSWER/mem[2][4][15] ), .s(n16741), .op(
        n2378) );
  mux2_1 U17382 ( .ip1(n16789), .ip2(\ANSWER/mem[2][5][15] ), .s(n16742), .op(
        n2377) );
  mux2_1 U17383 ( .ip1(n16819), .ip2(\ANSWER/mem[2][6][15] ), .s(n16743), .op(
        n2376) );
  mux2_1 U17384 ( .ip1(n16789), .ip2(\ANSWER/mem[2][7][15] ), .s(n16744), .op(
        n2375) );
  mux2_1 U17385 ( .ip1(n16789), .ip2(\ANSWER/mem[2][8][15] ), .s(n16745), .op(
        n2374) );
  mux2_1 U17386 ( .ip1(n16789), .ip2(\ANSWER/mem[2][9][15] ), .s(n16746), .op(
        n2373) );
  mux2_1 U17387 ( .ip1(n16819), .ip2(\ANSWER/mem[3][0][15] ), .s(n16747), .op(
        n2372) );
  mux2_1 U17388 ( .ip1(n16819), .ip2(\ANSWER/mem[3][1][15] ), .s(n16748), .op(
        n2371) );
  mux2_1 U17389 ( .ip1(n16819), .ip2(\ANSWER/mem[3][2][15] ), .s(n16749), .op(
        n2370) );
  mux2_1 U17390 ( .ip1(n16819), .ip2(\ANSWER/mem[3][3][15] ), .s(n16750), .op(
        n2369) );
  mux2_1 U17391 ( .ip1(n16819), .ip2(\ANSWER/mem[3][4][15] ), .s(n16751), .op(
        n2368) );
  mux2_1 U17392 ( .ip1(n16819), .ip2(\ANSWER/mem[3][5][15] ), .s(n16752), .op(
        n2367) );
  buf_1 U17393 ( .ip(n16789), .op(n16802) );
  mux2_1 U17394 ( .ip1(n16802), .ip2(\ANSWER/mem[3][6][15] ), .s(n16753), .op(
        n2366) );
  mux2_1 U17395 ( .ip1(n16789), .ip2(\ANSWER/mem[3][7][15] ), .s(n16754), .op(
        n2365) );
  mux2_1 U17396 ( .ip1(n16789), .ip2(\ANSWER/mem[3][8][15] ), .s(n16755), .op(
        n2364) );
  mux2_1 U17397 ( .ip1(n16789), .ip2(\ANSWER/mem[3][9][15] ), .s(n16756), .op(
        n2363) );
  mux2_1 U17398 ( .ip1(n16802), .ip2(\ANSWER/mem[4][0][15] ), .s(n16757), .op(
        n2362) );
  mux2_1 U17399 ( .ip1(n16802), .ip2(\ANSWER/mem[4][1][15] ), .s(n16758), .op(
        n2361) );
  mux2_1 U17400 ( .ip1(n16802), .ip2(\ANSWER/mem[4][2][15] ), .s(n16759), .op(
        n2360) );
  mux2_1 U17401 ( .ip1(n16802), .ip2(\ANSWER/mem[4][3][15] ), .s(n16760), .op(
        n2359) );
  mux2_1 U17402 ( .ip1(n16802), .ip2(\ANSWER/mem[4][4][15] ), .s(n16761), .op(
        n2358) );
  mux2_1 U17403 ( .ip1(n16802), .ip2(\ANSWER/mem[4][5][15] ), .s(n16762), .op(
        n2357) );
  mux2_1 U17404 ( .ip1(n16802), .ip2(\ANSWER/mem[4][6][15] ), .s(n16763), .op(
        n2356) );
  mux2_1 U17405 ( .ip1(n16802), .ip2(\ANSWER/mem[4][7][15] ), .s(n16764), .op(
        n2355) );
  mux2_1 U17406 ( .ip1(n16819), .ip2(\ANSWER/mem[4][8][15] ), .s(n16765), .op(
        n2354) );
  mux2_1 U17407 ( .ip1(n16789), .ip2(\ANSWER/mem[4][9][15] ), .s(n16766), .op(
        n2353) );
  mux2_1 U17408 ( .ip1(n16789), .ip2(\ANSWER/mem[5][0][15] ), .s(n16767), .op(
        n2352) );
  mux2_1 U17409 ( .ip1(n16789), .ip2(\ANSWER/mem[5][1][15] ), .s(n16768), .op(
        n2351) );
  mux2_1 U17410 ( .ip1(n16789), .ip2(\ANSWER/mem[5][2][15] ), .s(n16769), .op(
        n2350) );
  mux2_1 U17411 ( .ip1(n16789), .ip2(\ANSWER/mem[5][3][15] ), .s(n16770), .op(
        n2349) );
  mux2_1 U17412 ( .ip1(n16789), .ip2(\ANSWER/mem[5][4][15] ), .s(n16771), .op(
        n2348) );
  mux2_1 U17413 ( .ip1(n16789), .ip2(\ANSWER/mem[5][5][15] ), .s(n16772), .op(
        n2347) );
  mux2_1 U17414 ( .ip1(n16789), .ip2(\ANSWER/mem[5][6][15] ), .s(n16773), .op(
        n2346) );
  mux2_1 U17415 ( .ip1(n16789), .ip2(\ANSWER/mem[5][7][15] ), .s(n16774), .op(
        n2345) );
  mux2_1 U17416 ( .ip1(n16789), .ip2(\ANSWER/mem[5][8][15] ), .s(n16775), .op(
        n2344) );
  mux2_1 U17417 ( .ip1(n16789), .ip2(\ANSWER/mem[5][9][15] ), .s(n16776), .op(
        n2343) );
  mux2_1 U17418 ( .ip1(n16802), .ip2(\ANSWER/mem[6][0][15] ), .s(n16777), .op(
        n2342) );
  mux2_1 U17419 ( .ip1(n16802), .ip2(\ANSWER/mem[6][1][15] ), .s(n16778), .op(
        n2341) );
  mux2_1 U17420 ( .ip1(n16802), .ip2(\ANSWER/mem[6][2][15] ), .s(n16779), .op(
        n2340) );
  mux2_1 U17421 ( .ip1(n16802), .ip2(\ANSWER/mem[6][3][15] ), .s(n16780), .op(
        n2339) );
  mux2_1 U17422 ( .ip1(n16789), .ip2(\ANSWER/mem[6][4][15] ), .s(n16781), .op(
        n2338) );
  mux2_1 U17423 ( .ip1(n16789), .ip2(\ANSWER/mem[6][5][15] ), .s(n16782), .op(
        n2337) );
  mux2_1 U17424 ( .ip1(n16789), .ip2(\ANSWER/mem[6][6][15] ), .s(n16783), .op(
        n2336) );
  mux2_1 U17425 ( .ip1(n16789), .ip2(\ANSWER/mem[6][7][15] ), .s(n16784), .op(
        n2335) );
  mux2_1 U17426 ( .ip1(n16789), .ip2(\ANSWER/mem[6][8][15] ), .s(n16785), .op(
        n2334) );
  mux2_1 U17427 ( .ip1(n16789), .ip2(\ANSWER/mem[6][9][15] ), .s(n16786), .op(
        n2333) );
  mux2_1 U17428 ( .ip1(n16789), .ip2(\ANSWER/mem[7][0][15] ), .s(n16787), .op(
        n2332) );
  mux2_1 U17429 ( .ip1(n16789), .ip2(\ANSWER/mem[7][1][15] ), .s(n16788), .op(
        n2331) );
  mux2_1 U17430 ( .ip1(n16802), .ip2(\ANSWER/mem[7][2][15] ), .s(n16790), .op(
        n2330) );
  mux2_1 U17431 ( .ip1(n16802), .ip2(\ANSWER/mem[7][3][15] ), .s(n16791), .op(
        n2329) );
  mux2_1 U17432 ( .ip1(n16802), .ip2(\ANSWER/mem[7][4][15] ), .s(n16792), .op(
        n2328) );
  mux2_1 U17433 ( .ip1(n16802), .ip2(\ANSWER/mem[7][5][15] ), .s(n16793), .op(
        n2327) );
  mux2_1 U17434 ( .ip1(n16802), .ip2(\ANSWER/mem[7][6][15] ), .s(n16794), .op(
        n2326) );
  mux2_1 U17435 ( .ip1(n16802), .ip2(\ANSWER/mem[7][7][15] ), .s(n16795), .op(
        n2325) );
  mux2_1 U17436 ( .ip1(n16802), .ip2(\ANSWER/mem[7][8][15] ), .s(n16796), .op(
        n2324) );
  mux2_1 U17437 ( .ip1(n16802), .ip2(\ANSWER/mem[7][9][15] ), .s(n16797), .op(
        n2323) );
  mux2_1 U17438 ( .ip1(n16802), .ip2(\ANSWER/mem[8][0][15] ), .s(n16798), .op(
        n2322) );
  mux2_1 U17439 ( .ip1(n16802), .ip2(\ANSWER/mem[8][1][15] ), .s(n16799), .op(
        n2321) );
  mux2_1 U17440 ( .ip1(n16802), .ip2(\ANSWER/mem[8][2][15] ), .s(n16800), .op(
        n2320) );
  mux2_1 U17441 ( .ip1(n16802), .ip2(\ANSWER/mem[8][3][15] ), .s(n16801), .op(
        n2319) );
  mux2_1 U17442 ( .ip1(n16802), .ip2(\ANSWER/mem[8][4][15] ), .s(n16803), .op(
        n2318) );
  mux2_1 U17443 ( .ip1(n16819), .ip2(\ANSWER/mem[8][5][15] ), .s(n16804), .op(
        n2317) );
  mux2_1 U17444 ( .ip1(n16802), .ip2(\ANSWER/mem[8][6][15] ), .s(n16805), .op(
        n2316) );
  mux2_1 U17445 ( .ip1(n16819), .ip2(\ANSWER/mem[8][7][15] ), .s(n16806), .op(
        n2315) );
  mux2_1 U17446 ( .ip1(n16802), .ip2(\ANSWER/mem[8][8][15] ), .s(n16807), .op(
        n2314) );
  mux2_1 U17447 ( .ip1(n16789), .ip2(\ANSWER/mem[8][9][15] ), .s(n16808), .op(
        n2313) );
  mux2_1 U17448 ( .ip1(n16819), .ip2(\ANSWER/mem[9][0][15] ), .s(n16809), .op(
        n2312) );
  mux2_1 U17449 ( .ip1(n16802), .ip2(\ANSWER/mem[9][1][15] ), .s(n16810), .op(
        n2311) );
  mux2_1 U17450 ( .ip1(n16819), .ip2(\ANSWER/mem[9][2][15] ), .s(n16811), .op(
        n2310) );
  mux2_1 U17451 ( .ip1(n16802), .ip2(\ANSWER/mem[9][3][15] ), .s(n16812), .op(
        n2309) );
  mux2_1 U17452 ( .ip1(n16819), .ip2(\ANSWER/mem[9][4][15] ), .s(n16813), .op(
        n2308) );
  mux2_1 U17453 ( .ip1(n16802), .ip2(\ANSWER/mem[9][5][15] ), .s(n16814), .op(
        n2307) );
  mux2_1 U17454 ( .ip1(n16819), .ip2(\ANSWER/mem[9][6][15] ), .s(n16815), .op(
        n2306) );
  mux2_1 U17455 ( .ip1(n16819), .ip2(\ANSWER/mem[9][7][15] ), .s(n16816), .op(
        n2305) );
  mux2_1 U17456 ( .ip1(n16819), .ip2(\ANSWER/mem[9][8][15] ), .s(n16817), .op(
        n2304) );
  mux2_1 U17457 ( .ip1(n16819), .ip2(\ANSWER/mem[9][9][15] ), .s(n16818), .op(
        n2303) );
  buf_1 U17458 ( .ip(inputSramWe), .op(n16821) );
  buf_1 U17459 ( .ip(n16821), .op(n16820) );
  mux2_1 U17460 ( .ip1(\INPUTSRAM/mem_i[0][0] ), .ip2(pixels[0]), .s(n16820), 
        .op(n2302) );
  mux2_1 U17461 ( .ip1(\INPUTSRAM/mem_i[0][1] ), .ip2(pixels[1]), .s(n16820), 
        .op(n2301) );
  mux2_1 U17462 ( .ip1(\INPUTSRAM/mem_i[0][2] ), .ip2(pixels[2]), .s(n16820), 
        .op(n2300) );
  mux2_1 U17463 ( .ip1(\INPUTSRAM/mem_i[0][3] ), .ip2(pixels[3]), .s(n16820), 
        .op(n2299) );
  mux2_1 U17464 ( .ip1(\INPUTSRAM/mem_i[0][4] ), .ip2(pixels[4]), .s(n16820), 
        .op(n2298) );
  mux2_1 U17465 ( .ip1(\INPUTSRAM/mem_i[0][5] ), .ip2(pixels[5]), .s(n16820), 
        .op(n2297) );
  mux2_1 U17466 ( .ip1(\INPUTSRAM/mem_i[0][6] ), .ip2(pixels[6]), .s(n16820), 
        .op(n2296) );
  mux2_1 U17467 ( .ip1(\INPUTSRAM/mem_i[0][7] ), .ip2(pixels[7]), .s(n16820), 
        .op(n2295) );
  mux2_1 U17468 ( .ip1(\INPUTSRAM/mem_i[0][8] ), .ip2(pixels[8]), .s(n16820), 
        .op(n2294) );
  mux2_1 U17469 ( .ip1(\INPUTSRAM/mem_i[0][9] ), .ip2(pixels[9]), .s(n16820), 
        .op(n2293) );
  mux2_1 U17470 ( .ip1(\INPUTSRAM/mem_i[0][10] ), .ip2(pixels[10]), .s(n16820), 
        .op(n2292) );
  mux2_1 U17471 ( .ip1(\INPUTSRAM/mem_i[0][11] ), .ip2(pixels[11]), .s(n16820), 
        .op(n2291) );
  mux2_1 U17472 ( .ip1(\INPUTSRAM/mem_i[0][12] ), .ip2(pixels[12]), .s(n16820), 
        .op(n2290) );
  buf_1 U17473 ( .ip(inputSramWe), .op(n16822) );
  buf_1 U17474 ( .ip(n16822), .op(n16823) );
  mux2_1 U17475 ( .ip1(\INPUTSRAM/mem_i[0][13] ), .ip2(pixels[13]), .s(n16823), 
        .op(n2289) );
  mux2_1 U17476 ( .ip1(\INPUTSRAM/mem_i[0][14] ), .ip2(pixels[14]), .s(n16823), 
        .op(n2288) );
  mux2_1 U17477 ( .ip1(\INPUTSRAM/mem_i[1][0] ), .ip2(pixels[15]), .s(n16823), 
        .op(n2287) );
  mux2_1 U17478 ( .ip1(\INPUTSRAM/mem_i[1][1] ), .ip2(pixels[16]), .s(n16823), 
        .op(n2286) );
  mux2_1 U17479 ( .ip1(\INPUTSRAM/mem_i[1][2] ), .ip2(pixels[17]), .s(n16823), 
        .op(n2285) );
  mux2_1 U17480 ( .ip1(\INPUTSRAM/mem_i[1][3] ), .ip2(pixels[18]), .s(n16823), 
        .op(n2284) );
  mux2_1 U17481 ( .ip1(\INPUTSRAM/mem_i[1][4] ), .ip2(pixels[19]), .s(n16823), 
        .op(n2283) );
  mux2_1 U17482 ( .ip1(\INPUTSRAM/mem_i[1][5] ), .ip2(pixels[20]), .s(n16823), 
        .op(n2282) );
  mux2_1 U17483 ( .ip1(\INPUTSRAM/mem_i[1][6] ), .ip2(pixels[21]), .s(n16823), 
        .op(n2281) );
  mux2_1 U17484 ( .ip1(\INPUTSRAM/mem_i[1][7] ), .ip2(pixels[22]), .s(n16823), 
        .op(n2280) );
  mux2_1 U17485 ( .ip1(\INPUTSRAM/mem_i[1][8] ), .ip2(pixels[23]), .s(n16823), 
        .op(n2279) );
  mux2_1 U17486 ( .ip1(\INPUTSRAM/mem_i[1][9] ), .ip2(pixels[24]), .s(n16823), 
        .op(n2278) );
  mux2_1 U17487 ( .ip1(\INPUTSRAM/mem_i[1][10] ), .ip2(pixels[25]), .s(n16823), 
        .op(n2277) );
  mux2_1 U17488 ( .ip1(\INPUTSRAM/mem_i[1][11] ), .ip2(pixels[26]), .s(n16820), 
        .op(n2276) );
  mux2_1 U17489 ( .ip1(\INPUTSRAM/mem_i[1][12] ), .ip2(pixels[27]), .s(
        inputSramWe), .op(n2275) );
  mux2_1 U17490 ( .ip1(\INPUTSRAM/mem_i[1][13] ), .ip2(pixels[28]), .s(n16821), 
        .op(n2274) );
  buf_1 U17491 ( .ip(n16821), .op(n16826) );
  mux2_1 U17492 ( .ip1(\INPUTSRAM/mem_i[1][14] ), .ip2(pixels[29]), .s(n16826), 
        .op(n2273) );
  mux2_1 U17493 ( .ip1(\INPUTSRAM/mem_i[1][15] ), .ip2(pixels[30]), .s(n16820), 
        .op(n2272) );
  mux2_1 U17494 ( .ip1(\INPUTSRAM/mem_i[2][0] ), .ip2(pixels[32]), .s(
        inputSramWe), .op(n2271) );
  mux2_1 U17495 ( .ip1(\INPUTSRAM/mem_i[2][1] ), .ip2(pixels[33]), .s(n16821), 
        .op(n2270) );
  mux2_1 U17496 ( .ip1(\INPUTSRAM/mem_i[2][2] ), .ip2(pixels[34]), .s(n16826), 
        .op(n2269) );
  mux2_1 U17497 ( .ip1(\INPUTSRAM/mem_i[2][3] ), .ip2(pixels[35]), .s(n16820), 
        .op(n2268) );
  mux2_1 U17498 ( .ip1(\INPUTSRAM/mem_i[2][4] ), .ip2(pixels[36]), .s(
        inputSramWe), .op(n2267) );
  mux2_1 U17499 ( .ip1(\INPUTSRAM/mem_i[2][5] ), .ip2(pixels[37]), .s(n16821), 
        .op(n2266) );
  mux2_1 U17500 ( .ip1(\INPUTSRAM/mem_i[2][6] ), .ip2(pixels[38]), .s(n16826), 
        .op(n2265) );
  mux2_1 U17501 ( .ip1(\INPUTSRAM/mem_i[2][7] ), .ip2(pixels[39]), .s(n16820), 
        .op(n2264) );
  buf_1 U17502 ( .ip(n16822), .op(n16824) );
  mux2_1 U17503 ( .ip1(\INPUTSRAM/mem_i[2][8] ), .ip2(pixels[40]), .s(n16824), 
        .op(n2263) );
  mux2_1 U17504 ( .ip1(\INPUTSRAM/mem_i[2][9] ), .ip2(pixels[41]), .s(n16824), 
        .op(n2262) );
  mux2_1 U17505 ( .ip1(\INPUTSRAM/mem_i[2][10] ), .ip2(pixels[42]), .s(n16824), 
        .op(n2261) );
  mux2_1 U17506 ( .ip1(\INPUTSRAM/mem_i[2][11] ), .ip2(pixels[43]), .s(n16824), 
        .op(n2260) );
  mux2_1 U17507 ( .ip1(\INPUTSRAM/mem_i[2][12] ), .ip2(pixels[44]), .s(n16824), 
        .op(n2259) );
  mux2_1 U17508 ( .ip1(\INPUTSRAM/mem_i[2][13] ), .ip2(pixels[45]), .s(n16824), 
        .op(n2258) );
  mux2_1 U17509 ( .ip1(\INPUTSRAM/mem_i[2][14] ), .ip2(pixels[46]), .s(n16824), 
        .op(n2257) );
  mux2_1 U17510 ( .ip1(\INPUTSRAM/mem_i[3][0] ), .ip2(pixels[47]), .s(n16824), 
        .op(n2256) );
  mux2_1 U17511 ( .ip1(\INPUTSRAM/mem_i[3][1] ), .ip2(pixels[48]), .s(n16824), 
        .op(n2255) );
  mux2_1 U17512 ( .ip1(\INPUTSRAM/mem_i[3][2] ), .ip2(pixels[49]), .s(n16824), 
        .op(n2254) );
  mux2_1 U17513 ( .ip1(\INPUTSRAM/mem_i[3][3] ), .ip2(pixels[50]), .s(n16824), 
        .op(n2253) );
  mux2_1 U17514 ( .ip1(\INPUTSRAM/mem_i[3][4] ), .ip2(pixels[51]), .s(n16824), 
        .op(n2252) );
  mux2_1 U17515 ( .ip1(\INPUTSRAM/mem_i[3][5] ), .ip2(pixels[52]), .s(n16824), 
        .op(n2251) );
  mux2_1 U17516 ( .ip1(\INPUTSRAM/mem_i[3][6] ), .ip2(pixels[53]), .s(n16821), 
        .op(n2250) );
  mux2_1 U17517 ( .ip1(\INPUTSRAM/mem_i[3][7] ), .ip2(pixels[54]), .s(n16821), 
        .op(n2249) );
  mux2_1 U17518 ( .ip1(\INPUTSRAM/mem_i[3][8] ), .ip2(pixels[55]), .s(n16821), 
        .op(n2248) );
  mux2_1 U17519 ( .ip1(\INPUTSRAM/mem_i[3][9] ), .ip2(pixels[56]), .s(n16821), 
        .op(n2247) );
  mux2_1 U17520 ( .ip1(\INPUTSRAM/mem_i[3][10] ), .ip2(pixels[57]), .s(
        inputSramWe), .op(n2246) );
  mux2_1 U17521 ( .ip1(\INPUTSRAM/mem_i[3][11] ), .ip2(pixels[58]), .s(n16826), 
        .op(n2245) );
  mux2_1 U17522 ( .ip1(\INPUTSRAM/mem_i[3][12] ), .ip2(pixels[59]), .s(n16820), 
        .op(n2244) );
  mux2_1 U17523 ( .ip1(\INPUTSRAM/mem_i[3][13] ), .ip2(pixels[60]), .s(n16821), 
        .op(n2243) );
  mux2_1 U17524 ( .ip1(\INPUTSRAM/mem_i[3][14] ), .ip2(pixels[61]), .s(n16821), 
        .op(n2242) );
  mux2_1 U17525 ( .ip1(\INPUTSRAM/mem_i[3][15] ), .ip2(pixels[62]), .s(
        inputSramWe), .op(n2241) );
  mux2_1 U17526 ( .ip1(\INPUTSRAM/mem_i[4][0] ), .ip2(pixels[64]), .s(n16826), 
        .op(n2240) );
  mux2_1 U17527 ( .ip1(\INPUTSRAM/mem_i[4][1] ), .ip2(pixels[65]), .s(n16820), 
        .op(n2239) );
  mux2_1 U17528 ( .ip1(\INPUTSRAM/mem_i[4][2] ), .ip2(pixels[66]), .s(n16826), 
        .op(n2238) );
  mux2_1 U17529 ( .ip1(\INPUTSRAM/mem_i[4][3] ), .ip2(pixels[67]), .s(n16824), 
        .op(n2237) );
  mux2_1 U17530 ( .ip1(\INPUTSRAM/mem_i[4][4] ), .ip2(pixels[68]), .s(n16822), 
        .op(n2236) );
  buf_1 U17531 ( .ip(n16822), .op(n16825) );
  mux2_1 U17532 ( .ip1(\INPUTSRAM/mem_i[4][5] ), .ip2(pixels[69]), .s(n16825), 
        .op(n2235) );
  mux2_1 U17533 ( .ip1(\INPUTSRAM/mem_i[4][6] ), .ip2(pixels[70]), .s(n16823), 
        .op(n2234) );
  mux2_1 U17534 ( .ip1(\INPUTSRAM/mem_i[4][7] ), .ip2(pixels[71]), .s(n16824), 
        .op(n2233) );
  mux2_1 U17535 ( .ip1(\INPUTSRAM/mem_i[4][8] ), .ip2(pixels[72]), .s(n16822), 
        .op(n2232) );
  mux2_1 U17536 ( .ip1(\INPUTSRAM/mem_i[4][9] ), .ip2(pixels[73]), .s(n16825), 
        .op(n2231) );
  mux2_1 U17537 ( .ip1(\INPUTSRAM/mem_i[4][10] ), .ip2(pixels[74]), .s(n16823), 
        .op(n2230) );
  mux2_1 U17538 ( .ip1(\INPUTSRAM/mem_i[4][11] ), .ip2(pixels[75]), .s(n16824), 
        .op(n2229) );
  mux2_1 U17539 ( .ip1(\INPUTSRAM/mem_i[4][12] ), .ip2(pixels[76]), .s(n16822), 
        .op(n2228) );
  mux2_1 U17540 ( .ip1(\INPUTSRAM/mem_i[4][13] ), .ip2(pixels[77]), .s(
        inputSramWe), .op(n2227) );
  mux2_1 U17541 ( .ip1(\INPUTSRAM/mem_i[4][14] ), .ip2(pixels[78]), .s(n16825), 
        .op(n2226) );
  mux2_1 U17542 ( .ip1(\INPUTSRAM/mem_i[4][15] ), .ip2(pixels[79]), .s(n16823), 
        .op(n2225) );
  mux2_1 U17543 ( .ip1(\INPUTSRAM/mem_i[5][0] ), .ip2(pixels[80]), .s(n16821), 
        .op(n2224) );
  mux2_1 U17544 ( .ip1(\INPUTSRAM/mem_i[5][1] ), .ip2(pixels[81]), .s(n16821), 
        .op(n2223) );
  mux2_1 U17545 ( .ip1(\INPUTSRAM/mem_i[5][2] ), .ip2(pixels[82]), .s(
        inputSramWe), .op(n2222) );
  mux2_1 U17546 ( .ip1(\INPUTSRAM/mem_i[5][3] ), .ip2(pixels[83]), .s(n16826), 
        .op(n2221) );
  mux2_1 U17547 ( .ip1(\INPUTSRAM/mem_i[5][4] ), .ip2(pixels[84]), .s(n16820), 
        .op(n2220) );
  mux2_1 U17548 ( .ip1(\INPUTSRAM/mem_i[5][5] ), .ip2(pixels[85]), .s(n16821), 
        .op(n2219) );
  mux2_1 U17549 ( .ip1(\INPUTSRAM/mem_i[5][6] ), .ip2(pixels[86]), .s(n16821), 
        .op(n2218) );
  mux2_1 U17550 ( .ip1(\INPUTSRAM/mem_i[5][7] ), .ip2(pixels[87]), .s(n16821), 
        .op(n2217) );
  mux2_1 U17551 ( .ip1(\INPUTSRAM/mem_i[5][8] ), .ip2(pixels[88]), .s(
        inputSramWe), .op(n2216) );
  mux2_1 U17552 ( .ip1(\INPUTSRAM/mem_i[5][9] ), .ip2(pixels[89]), .s(n16826), 
        .op(n2215) );
  mux2_1 U17553 ( .ip1(\INPUTSRAM/mem_i[5][10] ), .ip2(pixels[90]), .s(n16820), 
        .op(n2214) );
  mux2_1 U17554 ( .ip1(\INPUTSRAM/mem_i[5][11] ), .ip2(pixels[91]), .s(
        inputSramWe), .op(n2213) );
  mux2_1 U17555 ( .ip1(\INPUTSRAM/mem_i[5][12] ), .ip2(pixels[92]), .s(n16821), 
        .op(n2212) );
  mux2_1 U17556 ( .ip1(\INPUTSRAM/mem_i[5][13] ), .ip2(pixels[93]), .s(n16822), 
        .op(n2211) );
  mux2_1 U17557 ( .ip1(\INPUTSRAM/mem_i[5][14] ), .ip2(pixels[94]), .s(n16822), 
        .op(n2210) );
  mux2_1 U17558 ( .ip1(\INPUTSRAM/mem_i[5][15] ), .ip2(pixels[95]), .s(n16822), 
        .op(n2209) );
  mux2_1 U17559 ( .ip1(\INPUTSRAM/mem_i[6][0] ), .ip2(pixels[96]), .s(n16822), 
        .op(n2208) );
  mux2_1 U17560 ( .ip1(\INPUTSRAM/mem_i[6][1] ), .ip2(pixels[97]), .s(n16822), 
        .op(n2207) );
  mux2_1 U17561 ( .ip1(\INPUTSRAM/mem_i[6][2] ), .ip2(pixels[98]), .s(n16822), 
        .op(n2206) );
  mux2_1 U17562 ( .ip1(\INPUTSRAM/mem_i[6][3] ), .ip2(pixels[99]), .s(n16822), 
        .op(n2205) );
  mux2_1 U17563 ( .ip1(\INPUTSRAM/mem_i[6][4] ), .ip2(pixels[100]), .s(n16825), 
        .op(n2204) );
  mux2_1 U17564 ( .ip1(\INPUTSRAM/mem_i[6][5] ), .ip2(pixels[101]), .s(n16823), 
        .op(n2203) );
  mux2_1 U17565 ( .ip1(\INPUTSRAM/mem_i[6][6] ), .ip2(pixels[102]), .s(n16824), 
        .op(n2202) );
  mux2_1 U17566 ( .ip1(\INPUTSRAM/mem_i[6][7] ), .ip2(pixels[103]), .s(n16823), 
        .op(n2201) );
  mux2_1 U17567 ( .ip1(\INPUTSRAM/mem_i[6][8] ), .ip2(pixels[104]), .s(n16822), 
        .op(n2200) );
  mux2_1 U17568 ( .ip1(\INPUTSRAM/mem_i[6][9] ), .ip2(pixels[105]), .s(n16825), 
        .op(n2199) );
  mux2_1 U17569 ( .ip1(\INPUTSRAM/mem_i[6][10] ), .ip2(pixels[106]), .s(n16821), .op(n2198) );
  mux2_1 U17570 ( .ip1(\INPUTSRAM/mem_i[6][11] ), .ip2(pixels[107]), .s(
        inputSramWe), .op(n2197) );
  mux2_1 U17571 ( .ip1(\INPUTSRAM/mem_i[6][12] ), .ip2(pixels[108]), .s(n16826), .op(n2196) );
  mux2_1 U17572 ( .ip1(\INPUTSRAM/mem_i[6][13] ), .ip2(pixels[109]), .s(n16821), .op(n2195) );
  mux2_1 U17573 ( .ip1(\INPUTSRAM/mem_i[6][14] ), .ip2(pixels[110]), .s(
        inputSramWe), .op(n2194) );
  mux2_1 U17574 ( .ip1(\INPUTSRAM/mem_i[6][15] ), .ip2(pixels[111]), .s(n16826), .op(n2193) );
  mux2_1 U17575 ( .ip1(\INPUTSRAM/mem_i[7][0] ), .ip2(pixels[112]), .s(n16821), 
        .op(n2192) );
  mux2_1 U17576 ( .ip1(\INPUTSRAM/mem_i[7][1] ), .ip2(pixels[113]), .s(
        inputSramWe), .op(n2191) );
  mux2_1 U17577 ( .ip1(\INPUTSRAM/mem_i[7][2] ), .ip2(pixels[114]), .s(n16826), 
        .op(n2190) );
  mux2_1 U17578 ( .ip1(\INPUTSRAM/mem_i[7][3] ), .ip2(pixels[115]), .s(n16821), 
        .op(n2189) );
  mux2_1 U17579 ( .ip1(\INPUTSRAM/mem_i[7][4] ), .ip2(pixels[116]), .s(
        inputSramWe), .op(n2188) );
  mux2_1 U17580 ( .ip1(\INPUTSRAM/mem_i[7][5] ), .ip2(pixels[117]), .s(n16826), 
        .op(n2187) );
  mux2_1 U17581 ( .ip1(\INPUTSRAM/mem_i[7][6] ), .ip2(pixels[118]), .s(n16821), 
        .op(n2186) );
  mux2_1 U17582 ( .ip1(\INPUTSRAM/mem_i[7][7] ), .ip2(pixels[119]), .s(n16822), 
        .op(n2185) );
  mux2_1 U17583 ( .ip1(\INPUTSRAM/mem_i[7][8] ), .ip2(pixels[120]), .s(n16822), 
        .op(n2184) );
  mux2_1 U17584 ( .ip1(\INPUTSRAM/mem_i[7][9] ), .ip2(pixels[121]), .s(n16822), 
        .op(n2183) );
  mux2_1 U17585 ( .ip1(\INPUTSRAM/mem_i[7][10] ), .ip2(pixels[122]), .s(n16822), .op(n2182) );
  mux2_1 U17586 ( .ip1(\INPUTSRAM/mem_i[7][11] ), .ip2(pixels[123]), .s(n16825), .op(n2181) );
  mux2_1 U17587 ( .ip1(\INPUTSRAM/mem_i[7][12] ), .ip2(pixels[124]), .s(n16823), .op(n2180) );
  mux2_1 U17588 ( .ip1(\INPUTSRAM/mem_i[7][13] ), .ip2(pixels[125]), .s(n16824), .op(n2179) );
  mux2_1 U17589 ( .ip1(\INPUTSRAM/mem_i[7][14] ), .ip2(pixels[126]), .s(n16822), .op(n2178) );
  mux2_1 U17590 ( .ip1(\INPUTSRAM/mem_i[7][15] ), .ip2(pixels[127]), .s(n16822), .op(n2177) );
  mux2_1 U17591 ( .ip1(\INPUTSRAM/mem_i[8][0] ), .ip2(pixels[128]), .s(n16822), 
        .op(n2176) );
  mux2_1 U17592 ( .ip1(\INPUTSRAM/mem_i[8][1] ), .ip2(pixels[129]), .s(n16825), 
        .op(n2175) );
  mux2_1 U17593 ( .ip1(\INPUTSRAM/mem_i[8][2] ), .ip2(pixels[130]), .s(n16823), 
        .op(n2174) );
  mux2_1 U17594 ( .ip1(\INPUTSRAM/mem_i[8][3] ), .ip2(pixels[131]), .s(n16824), 
        .op(n2173) );
  mux2_1 U17595 ( .ip1(\INPUTSRAM/mem_i[8][4] ), .ip2(pixels[132]), .s(n16826), 
        .op(n2172) );
  mux2_1 U17596 ( .ip1(\INPUTSRAM/mem_i[8][5] ), .ip2(pixels[133]), .s(n16826), 
        .op(n2171) );
  mux2_1 U17597 ( .ip1(\INPUTSRAM/mem_i[8][6] ), .ip2(pixels[134]), .s(
        inputSramWe), .op(n2170) );
  mux2_1 U17598 ( .ip1(\INPUTSRAM/mem_i[8][7] ), .ip2(pixels[135]), .s(n16826), 
        .op(n2169) );
  mux2_1 U17599 ( .ip1(\INPUTSRAM/mem_i[8][8] ), .ip2(pixels[136]), .s(
        inputSramWe), .op(n2168) );
  mux2_1 U17600 ( .ip1(\INPUTSRAM/mem_i[8][9] ), .ip2(pixels[137]), .s(n16826), 
        .op(n2167) );
  mux2_1 U17601 ( .ip1(\INPUTSRAM/mem_i[8][10] ), .ip2(pixels[138]), .s(
        inputSramWe), .op(n2166) );
  mux2_1 U17602 ( .ip1(\INPUTSRAM/mem_i[8][11] ), .ip2(pixels[139]), .s(n16826), .op(n2165) );
  mux2_1 U17603 ( .ip1(\INPUTSRAM/mem_i[8][12] ), .ip2(pixels[140]), .s(
        inputSramWe), .op(n2164) );
  mux2_1 U17604 ( .ip1(\INPUTSRAM/mem_i[8][13] ), .ip2(pixels[141]), .s(n16826), .op(n2163) );
  mux2_1 U17605 ( .ip1(\INPUTSRAM/mem_i[8][14] ), .ip2(pixels[142]), .s(
        inputSramWe), .op(n2162) );
  mux2_1 U17606 ( .ip1(\INPUTSRAM/mem_i[8][15] ), .ip2(pixels[143]), .s(n16826), .op(n2161) );
  mux2_1 U17607 ( .ip1(\INPUTSRAM/mem_i[9][0] ), .ip2(pixels[144]), .s(
        inputSramWe), .op(n2160) );
  mux2_1 U17608 ( .ip1(\INPUTSRAM/mem_i[9][1] ), .ip2(pixels[145]), .s(n16825), 
        .op(n2159) );
  mux2_1 U17609 ( .ip1(\INPUTSRAM/mem_i[9][2] ), .ip2(pixels[146]), .s(n16825), 
        .op(n2158) );
  mux2_1 U17610 ( .ip1(\INPUTSRAM/mem_i[9][3] ), .ip2(pixels[147]), .s(n16825), 
        .op(n2157) );
  mux2_1 U17611 ( .ip1(\INPUTSRAM/mem_i[9][4] ), .ip2(pixels[148]), .s(n16825), 
        .op(n2156) );
  mux2_1 U17612 ( .ip1(\INPUTSRAM/mem_i[9][5] ), .ip2(pixels[149]), .s(n16825), 
        .op(n2155) );
  mux2_1 U17613 ( .ip1(\INPUTSRAM/mem_i[9][6] ), .ip2(pixels[150]), .s(n16825), 
        .op(n2154) );
  mux2_1 U17614 ( .ip1(\INPUTSRAM/mem_i[9][7] ), .ip2(pixels[151]), .s(n16825), 
        .op(n2153) );
  mux2_1 U17615 ( .ip1(\INPUTSRAM/mem_i[9][8] ), .ip2(pixels[152]), .s(n16825), 
        .op(n2152) );
  mux2_1 U17616 ( .ip1(\INPUTSRAM/mem_i[9][9] ), .ip2(pixels[153]), .s(n16825), 
        .op(n2151) );
  mux2_1 U17617 ( .ip1(\INPUTSRAM/mem_i[9][10] ), .ip2(pixels[154]), .s(n16825), .op(n2150) );
  mux2_1 U17618 ( .ip1(\INPUTSRAM/mem_i[9][11] ), .ip2(pixels[155]), .s(n16825), .op(n2149) );
  mux2_1 U17619 ( .ip1(\INPUTSRAM/mem_i[9][12] ), .ip2(pixels[156]), .s(n16825), .op(n2148) );
  mux2_1 U17620 ( .ip1(\INPUTSRAM/mem_i[9][13] ), .ip2(pixels[157]), .s(n16825), .op(n2147) );
  mux2_1 U17621 ( .ip1(\INPUTSRAM/mem_i[9][14] ), .ip2(pixels[158]), .s(n16826), .op(n2146) );
  mux2_1 U17622 ( .ip1(\INPUTSRAM/mem_i[9][15] ), .ip2(pixels[159]), .s(n16826), .op(n2145) );
  buf_1 U17623 ( .ip(n17289), .op(n17282) );
  nand2_1 U17624 ( .ip1(column[8]), .ip2(n17282), .op(n16830) );
  nand2_1 U17625 ( .ip1(n17243), .ip2(n16860), .op(n17244) );
  nand2_1 U17626 ( .ip1(\ROUTEDATA/regData [8]), .ip2(n17244), .op(n16829) );
  nand2_1 U17627 ( .ip1(n16827), .ip2(n17241), .op(n16865) );
  inv_1 U17628 ( .ip(n16865), .op(n16861) );
  nand2_1 U17629 ( .ip1(n17243), .ip2(n16861), .op(n16828) );
  nand3_1 U17630 ( .ip1(n16830), .ip2(n16829), .ip3(n16828), .op(n2128) );
  nand2_1 U17631 ( .ip1(column[24]), .ip2(n17282), .op(n16834) );
  or2_1 U17632 ( .ip1(n17229), .ip2(n16831), .op(n17249) );
  nand2_1 U17633 ( .ip1(n16860), .ip2(n17249), .op(n17250) );
  nand2_1 U17634 ( .ip1(\ROUTEDATA/regData [24]), .ip2(n17250), .op(n16833) );
  nand2_1 U17635 ( .ip1(n16861), .ip2(n17249), .op(n16832) );
  nand3_1 U17636 ( .ip1(n16834), .ip2(n16833), .ip3(n16832), .op(n2127) );
  nand2_1 U17637 ( .ip1(column[40]), .ip2(n17282), .op(n16838) );
  or2_1 U17638 ( .ip1(n17229), .ip2(n16835), .op(n17210) );
  nand2_1 U17639 ( .ip1(n16861), .ip2(n17210), .op(n16837) );
  nand2_1 U17640 ( .ip1(n16860), .ip2(n17210), .op(n17255) );
  nand2_1 U17641 ( .ip1(\ROUTEDATA/regData [40]), .ip2(n17255), .op(n16836) );
  nand3_1 U17642 ( .ip1(n16838), .ip2(n16837), .ip3(n16836), .op(n2126) );
  nand2_1 U17643 ( .ip1(column[56]), .ip2(n17282), .op(n16842) );
  or2_1 U17644 ( .ip1(n17229), .ip2(n16839), .op(n17257) );
  nand2_1 U17645 ( .ip1(n16861), .ip2(n17257), .op(n16841) );
  nand2_1 U17646 ( .ip1(n16860), .ip2(n17257), .op(n17258) );
  nand2_1 U17647 ( .ip1(\ROUTEDATA/regData [56]), .ip2(n17258), .op(n16840) );
  nand3_1 U17648 ( .ip1(n16842), .ip2(n16841), .ip3(n16840), .op(n2125) );
  nand2_1 U17649 ( .ip1(column[72]), .ip2(n17282), .op(n16846) );
  or2_1 U17650 ( .ip1(n17229), .ip2(n16843), .op(n17262) );
  nand2_1 U17651 ( .ip1(n16860), .ip2(n17262), .op(n17263) );
  nand2_1 U17652 ( .ip1(\ROUTEDATA/regData [72]), .ip2(n17263), .op(n16845) );
  nand2_1 U17653 ( .ip1(n16861), .ip2(n17262), .op(n16844) );
  nand3_1 U17654 ( .ip1(n16846), .ip2(n16845), .ip3(n16844), .op(n2124) );
  nand2_1 U17655 ( .ip1(column[88]), .ip2(n17282), .op(n16850) );
  or2_1 U17656 ( .ip1(n17229), .ip2(n16847), .op(n17267) );
  nand2_1 U17657 ( .ip1(n16861), .ip2(n17267), .op(n16849) );
  nand2_1 U17658 ( .ip1(n16860), .ip2(n17267), .op(n17268) );
  nand2_1 U17659 ( .ip1(\ROUTEDATA/regData [88]), .ip2(n17268), .op(n16848) );
  nand3_1 U17660 ( .ip1(n16850), .ip2(n16849), .ip3(n16848), .op(n2123) );
  buf_1 U17661 ( .ip(n17282), .op(n17248) );
  nand2_1 U17662 ( .ip1(column[104]), .ip2(n17248), .op(n16854) );
  or2_1 U17663 ( .ip1(n17229), .ip2(n16851), .op(n17272) );
  nand2_1 U17664 ( .ip1(n16861), .ip2(n17272), .op(n16853) );
  nand2_1 U17665 ( .ip1(n16860), .ip2(n17272), .op(n17273) );
  nand2_1 U17666 ( .ip1(\ROUTEDATA/regData [104]), .ip2(n17273), .op(n16852)
         );
  nand3_1 U17667 ( .ip1(n16854), .ip2(n16853), .ip3(n16852), .op(n2122) );
  nand2_1 U17668 ( .ip1(column[120]), .ip2(n17248), .op(n16858) );
  or2_1 U17669 ( .ip1(n17229), .ip2(n16855), .op(n17277) );
  nand2_1 U17670 ( .ip1(n16861), .ip2(n17277), .op(n16857) );
  nand2_1 U17671 ( .ip1(n16860), .ip2(n17277), .op(n17278) );
  nand2_1 U17672 ( .ip1(\ROUTEDATA/regData [120]), .ip2(n17278), .op(n16856)
         );
  nand3_1 U17673 ( .ip1(n16858), .ip2(n16857), .ip3(n16856), .op(n2121) );
  nand2_1 U17674 ( .ip1(column[136]), .ip2(n17248), .op(n16864) );
  nor2_1 U17675 ( .ip1(n17229), .ip2(n16859), .op(n17233) );
  inv_1 U17676 ( .ip(n17233), .op(n17283) );
  nand2_1 U17677 ( .ip1(n16860), .ip2(n17283), .op(n17285) );
  nand2_1 U17678 ( .ip1(\ROUTEDATA/regData [136]), .ip2(n17285), .op(n16863)
         );
  nand2_1 U17679 ( .ip1(n16861), .ip2(n17283), .op(n16862) );
  nand3_1 U17680 ( .ip1(n16864), .ip2(n16863), .ip3(n16862), .op(n2120) );
  nand2_1 U17681 ( .ip1(n17289), .ip2(column[152]), .op(n16866) );
  nand2_1 U17682 ( .ip1(n16866), .ip2(n16865), .op(n16867) );
  nor2_1 U17683 ( .ip1(n17229), .ip2(weight2_loadNextRow), .op(n17292) );
  mux2_1 U17684 ( .ip1(n16867), .ip2(\ROUTEDATA/regData [152]), .s(n17292), 
        .op(n2119) );
  nand2_1 U17685 ( .ip1(n17289), .ip2(column[9]), .op(n16869) );
  nand2_1 U17686 ( .ip1(\ROUTEDATA/regData [9]), .ip2(n17244), .op(n16868) );
  nand2_1 U17687 ( .ip1(n16869), .ip2(n16868), .op(n2118) );
  nand2_1 U17688 ( .ip1(n17289), .ip2(column[25]), .op(n16871) );
  nand2_1 U17689 ( .ip1(\ROUTEDATA/regData [25]), .ip2(n17250), .op(n16870) );
  nand2_1 U17690 ( .ip1(n16871), .ip2(n16870), .op(n2117) );
  nand2_1 U17691 ( .ip1(n17289), .ip2(column[41]), .op(n16873) );
  nand2_1 U17692 ( .ip1(\ROUTEDATA/regData [41]), .ip2(n17255), .op(n16872) );
  nand2_1 U17693 ( .ip1(n16873), .ip2(n16872), .op(n2116) );
  nand2_1 U17694 ( .ip1(n17289), .ip2(column[57]), .op(n16875) );
  nand2_1 U17695 ( .ip1(\ROUTEDATA/regData [57]), .ip2(n17258), .op(n16874) );
  nand2_1 U17696 ( .ip1(n16875), .ip2(n16874), .op(n2115) );
  nand2_1 U17697 ( .ip1(n17229), .ip2(column[73]), .op(n16877) );
  nand2_1 U17698 ( .ip1(\ROUTEDATA/regData [73]), .ip2(n17263), .op(n16876) );
  nand2_1 U17699 ( .ip1(n16877), .ip2(n16876), .op(n2114) );
  nand2_1 U17700 ( .ip1(n17229), .ip2(column[89]), .op(n16879) );
  nand2_1 U17701 ( .ip1(\ROUTEDATA/regData [89]), .ip2(n17268), .op(n16878) );
  nand2_1 U17702 ( .ip1(n16879), .ip2(n16878), .op(n2113) );
  nand2_1 U17703 ( .ip1(n17289), .ip2(column[105]), .op(n16881) );
  nand2_1 U17704 ( .ip1(\ROUTEDATA/regData [105]), .ip2(n17273), .op(n16880)
         );
  nand2_1 U17705 ( .ip1(n16881), .ip2(n16880), .op(n2112) );
  nand2_1 U17706 ( .ip1(n17289), .ip2(column[121]), .op(n16883) );
  nand2_1 U17707 ( .ip1(\ROUTEDATA/regData [121]), .ip2(n17278), .op(n16882)
         );
  nand2_1 U17708 ( .ip1(n16883), .ip2(n16882), .op(n2111) );
  nand2_1 U17709 ( .ip1(n17289), .ip2(column[137]), .op(n16885) );
  nand2_1 U17710 ( .ip1(\ROUTEDATA/regData [137]), .ip2(n17285), .op(n16884)
         );
  nand2_1 U17711 ( .ip1(n16885), .ip2(n16884), .op(n2110) );
  nand2_1 U17712 ( .ip1(n17292), .ip2(\ROUTEDATA/regData [153]), .op(n16887)
         );
  nand2_1 U17713 ( .ip1(column[153]), .ip2(n17248), .op(n16886) );
  nand2_1 U17714 ( .ip1(n16887), .ip2(n16886), .op(n2109) );
  nand2_1 U17715 ( .ip1(n17229), .ip2(column[10]), .op(n16889) );
  nand2_1 U17716 ( .ip1(\ROUTEDATA/regData [10]), .ip2(n17244), .op(n16888) );
  nand2_1 U17717 ( .ip1(n16889), .ip2(n16888), .op(n2108) );
  nand2_1 U17718 ( .ip1(n17229), .ip2(column[26]), .op(n16891) );
  nand2_1 U17719 ( .ip1(\ROUTEDATA/regData [26]), .ip2(n17250), .op(n16890) );
  nand2_1 U17720 ( .ip1(n16891), .ip2(n16890), .op(n2107) );
  nand2_1 U17721 ( .ip1(n17289), .ip2(column[42]), .op(n16893) );
  nand2_1 U17722 ( .ip1(\ROUTEDATA/regData [42]), .ip2(n17255), .op(n16892) );
  nand2_1 U17723 ( .ip1(n16893), .ip2(n16892), .op(n2106) );
  nand2_1 U17724 ( .ip1(n17289), .ip2(column[58]), .op(n16895) );
  nand2_1 U17725 ( .ip1(\ROUTEDATA/regData [58]), .ip2(n17258), .op(n16894) );
  nand2_1 U17726 ( .ip1(n16895), .ip2(n16894), .op(n2105) );
  nand2_1 U17727 ( .ip1(n17289), .ip2(column[74]), .op(n16897) );
  nand2_1 U17728 ( .ip1(\ROUTEDATA/regData [74]), .ip2(n17263), .op(n16896) );
  nand2_1 U17729 ( .ip1(n16897), .ip2(n16896), .op(n2104) );
  nand2_1 U17730 ( .ip1(n17289), .ip2(column[90]), .op(n16899) );
  nand2_1 U17731 ( .ip1(\ROUTEDATA/regData [90]), .ip2(n17268), .op(n16898) );
  nand2_1 U17732 ( .ip1(n16899), .ip2(n16898), .op(n2103) );
  nand2_1 U17733 ( .ip1(n17289), .ip2(column[106]), .op(n16901) );
  nand2_1 U17734 ( .ip1(\ROUTEDATA/regData [106]), .ip2(n17273), .op(n16900)
         );
  nand2_1 U17735 ( .ip1(n16901), .ip2(n16900), .op(n2102) );
  nand2_1 U17736 ( .ip1(n17289), .ip2(column[122]), .op(n16903) );
  nand2_1 U17737 ( .ip1(\ROUTEDATA/regData [122]), .ip2(n17278), .op(n16902)
         );
  nand2_1 U17738 ( .ip1(n16903), .ip2(n16902), .op(n2101) );
  nand2_1 U17739 ( .ip1(n17289), .ip2(column[138]), .op(n16905) );
  nand2_1 U17740 ( .ip1(\ROUTEDATA/regData [138]), .ip2(n17285), .op(n16904)
         );
  nand2_1 U17741 ( .ip1(n16905), .ip2(n16904), .op(n2100) );
  nand2_1 U17742 ( .ip1(n17292), .ip2(\ROUTEDATA/regData [154]), .op(n16907)
         );
  nand2_1 U17743 ( .ip1(column[154]), .ip2(n17248), .op(n16906) );
  nand2_1 U17744 ( .ip1(n16907), .ip2(n16906), .op(n2099) );
  nand2_1 U17745 ( .ip1(n17289), .ip2(column[11]), .op(n16909) );
  nand2_1 U17746 ( .ip1(\ROUTEDATA/regData [11]), .ip2(n17244), .op(n16908) );
  nand2_1 U17747 ( .ip1(n16909), .ip2(n16908), .op(n2098) );
  nand2_1 U17748 ( .ip1(n17289), .ip2(column[27]), .op(n16911) );
  nand2_1 U17749 ( .ip1(\ROUTEDATA/regData [27]), .ip2(n17250), .op(n16910) );
  nand2_1 U17750 ( .ip1(n16911), .ip2(n16910), .op(n2097) );
  nand2_1 U17751 ( .ip1(n17289), .ip2(column[43]), .op(n16913) );
  nand2_1 U17752 ( .ip1(\ROUTEDATA/regData [43]), .ip2(n17255), .op(n16912) );
  nand2_1 U17753 ( .ip1(n16913), .ip2(n16912), .op(n2096) );
  nand2_1 U17754 ( .ip1(n17289), .ip2(column[59]), .op(n16915) );
  nand2_1 U17755 ( .ip1(\ROUTEDATA/regData [59]), .ip2(n17258), .op(n16914) );
  nand2_1 U17756 ( .ip1(n16915), .ip2(n16914), .op(n2095) );
  nand2_1 U17757 ( .ip1(n17289), .ip2(column[75]), .op(n16917) );
  nand2_1 U17758 ( .ip1(\ROUTEDATA/regData [75]), .ip2(n17263), .op(n16916) );
  nand2_1 U17759 ( .ip1(n16917), .ip2(n16916), .op(n2094) );
  nand2_1 U17760 ( .ip1(n17289), .ip2(column[91]), .op(n16919) );
  nand2_1 U17761 ( .ip1(\ROUTEDATA/regData [91]), .ip2(n17268), .op(n16918) );
  nand2_1 U17762 ( .ip1(n16919), .ip2(n16918), .op(n2093) );
  nand2_1 U17763 ( .ip1(n17289), .ip2(column[107]), .op(n16921) );
  nand2_1 U17764 ( .ip1(\ROUTEDATA/regData [107]), .ip2(n17273), .op(n16920)
         );
  nand2_1 U17765 ( .ip1(n16921), .ip2(n16920), .op(n2092) );
  nand2_1 U17766 ( .ip1(n17248), .ip2(column[123]), .op(n16923) );
  nand2_1 U17767 ( .ip1(\ROUTEDATA/regData [123]), .ip2(n17278), .op(n16922)
         );
  nand2_1 U17768 ( .ip1(n16923), .ip2(n16922), .op(n2091) );
  nand2_1 U17769 ( .ip1(n17248), .ip2(column[139]), .op(n16925) );
  nand2_1 U17770 ( .ip1(\ROUTEDATA/regData [139]), .ip2(n17285), .op(n16924)
         );
  nand2_1 U17771 ( .ip1(n16925), .ip2(n16924), .op(n2090) );
  nand2_1 U17772 ( .ip1(n17292), .ip2(\ROUTEDATA/regData [155]), .op(n16927)
         );
  nand2_1 U17773 ( .ip1(column[155]), .ip2(n17282), .op(n16926) );
  nand2_1 U17774 ( .ip1(n16927), .ip2(n16926), .op(n2089) );
  nand2_1 U17775 ( .ip1(n17248), .ip2(column[12]), .op(n16929) );
  nand2_1 U17776 ( .ip1(\ROUTEDATA/regData [12]), .ip2(n17244), .op(n16928) );
  nand2_1 U17777 ( .ip1(n16929), .ip2(n16928), .op(n2088) );
  nand2_1 U17778 ( .ip1(n17248), .ip2(column[28]), .op(n16931) );
  nand2_1 U17779 ( .ip1(\ROUTEDATA/regData [28]), .ip2(n17250), .op(n16930) );
  nand2_1 U17780 ( .ip1(n16931), .ip2(n16930), .op(n2087) );
  nand2_1 U17781 ( .ip1(n17248), .ip2(column[44]), .op(n16933) );
  nand2_1 U17782 ( .ip1(\ROUTEDATA/regData [44]), .ip2(n17255), .op(n16932) );
  nand2_1 U17783 ( .ip1(n16933), .ip2(n16932), .op(n2086) );
  nand2_1 U17784 ( .ip1(n17229), .ip2(column[60]), .op(n16935) );
  nand2_1 U17785 ( .ip1(\ROUTEDATA/regData [60]), .ip2(n17258), .op(n16934) );
  nand2_1 U17786 ( .ip1(n16935), .ip2(n16934), .op(n2085) );
  nand2_1 U17787 ( .ip1(n17229), .ip2(column[76]), .op(n16937) );
  nand2_1 U17788 ( .ip1(\ROUTEDATA/regData [76]), .ip2(n17263), .op(n16936) );
  nand2_1 U17789 ( .ip1(n16937), .ip2(n16936), .op(n2084) );
  nand2_1 U17790 ( .ip1(n17229), .ip2(column[92]), .op(n16939) );
  nand2_1 U17791 ( .ip1(\ROUTEDATA/regData [92]), .ip2(n17268), .op(n16938) );
  nand2_1 U17792 ( .ip1(n16939), .ip2(n16938), .op(n2083) );
  nand2_1 U17793 ( .ip1(n17289), .ip2(column[108]), .op(n16941) );
  nand2_1 U17794 ( .ip1(\ROUTEDATA/regData [108]), .ip2(n17273), .op(n16940)
         );
  nand2_1 U17795 ( .ip1(n16941), .ip2(n16940), .op(n2082) );
  nand2_1 U17796 ( .ip1(n17229), .ip2(column[124]), .op(n16943) );
  nand2_1 U17797 ( .ip1(\ROUTEDATA/regData [124]), .ip2(n17278), .op(n16942)
         );
  nand2_1 U17798 ( .ip1(n16943), .ip2(n16942), .op(n2081) );
  nand2_1 U17799 ( .ip1(n17229), .ip2(column[140]), .op(n16945) );
  nand2_1 U17800 ( .ip1(\ROUTEDATA/regData [140]), .ip2(n17285), .op(n16944)
         );
  nand2_1 U17801 ( .ip1(n16945), .ip2(n16944), .op(n2080) );
  nand2_1 U17802 ( .ip1(n17292), .ip2(\ROUTEDATA/regData [156]), .op(n16947)
         );
  nand2_1 U17803 ( .ip1(column[156]), .ip2(n17282), .op(n16946) );
  nand2_1 U17804 ( .ip1(n16947), .ip2(n16946), .op(n2079) );
  nand2_1 U17805 ( .ip1(n17229), .ip2(column[13]), .op(n16949) );
  nand2_1 U17806 ( .ip1(\ROUTEDATA/regData [13]), .ip2(n17244), .op(n16948) );
  nand2_1 U17807 ( .ip1(n16949), .ip2(n16948), .op(n2078) );
  nand2_1 U17808 ( .ip1(n17229), .ip2(column[29]), .op(n16951) );
  nand2_1 U17809 ( .ip1(\ROUTEDATA/regData [29]), .ip2(n17250), .op(n16950) );
  nand2_1 U17810 ( .ip1(n16951), .ip2(n16950), .op(n2077) );
  nand2_1 U17811 ( .ip1(n17229), .ip2(column[45]), .op(n16953) );
  nand2_1 U17812 ( .ip1(\ROUTEDATA/regData [45]), .ip2(n17255), .op(n16952) );
  nand2_1 U17813 ( .ip1(n16953), .ip2(n16952), .op(n2076) );
  nand2_1 U17814 ( .ip1(n17229), .ip2(column[61]), .op(n16955) );
  nand2_1 U17815 ( .ip1(\ROUTEDATA/regData [61]), .ip2(n17258), .op(n16954) );
  nand2_1 U17816 ( .ip1(n16955), .ip2(n16954), .op(n2075) );
  nand2_1 U17817 ( .ip1(n17229), .ip2(column[77]), .op(n16957) );
  nand2_1 U17818 ( .ip1(\ROUTEDATA/regData [77]), .ip2(n17263), .op(n16956) );
  nand2_1 U17819 ( .ip1(n16957), .ip2(n16956), .op(n2074) );
  nand2_1 U17820 ( .ip1(n17229), .ip2(column[93]), .op(n16959) );
  nand2_1 U17821 ( .ip1(\ROUTEDATA/regData [93]), .ip2(n17268), .op(n16958) );
  nand2_1 U17822 ( .ip1(n16959), .ip2(n16958), .op(n2073) );
  nand2_1 U17823 ( .ip1(n17229), .ip2(column[109]), .op(n16961) );
  nand2_1 U17824 ( .ip1(\ROUTEDATA/regData [109]), .ip2(n17273), .op(n16960)
         );
  nand2_1 U17825 ( .ip1(n16961), .ip2(n16960), .op(n2072) );
  nand2_1 U17826 ( .ip1(n17229), .ip2(column[125]), .op(n16963) );
  nand2_1 U17827 ( .ip1(\ROUTEDATA/regData [125]), .ip2(n17278), .op(n16962)
         );
  nand2_1 U17828 ( .ip1(n16963), .ip2(n16962), .op(n2071) );
  nand2_1 U17829 ( .ip1(n17229), .ip2(column[141]), .op(n16965) );
  nand2_1 U17830 ( .ip1(\ROUTEDATA/regData [141]), .ip2(n17285), .op(n16964)
         );
  nand2_1 U17831 ( .ip1(n16965), .ip2(n16964), .op(n2070) );
  nand2_1 U17832 ( .ip1(n17292), .ip2(\ROUTEDATA/regData [157]), .op(n16967)
         );
  nand2_1 U17833 ( .ip1(column[157]), .ip2(n17229), .op(n16966) );
  nand2_1 U17834 ( .ip1(n16967), .ip2(n16966), .op(n2069) );
  nand2_1 U17835 ( .ip1(n17229), .ip2(column[14]), .op(n16969) );
  nand2_1 U17836 ( .ip1(\ROUTEDATA/regData [14]), .ip2(n17244), .op(n16968) );
  nand2_1 U17837 ( .ip1(n16969), .ip2(n16968), .op(n2068) );
  nand2_1 U17838 ( .ip1(n17229), .ip2(column[30]), .op(n16971) );
  nand2_1 U17839 ( .ip1(\ROUTEDATA/regData [30]), .ip2(n17250), .op(n16970) );
  nand2_1 U17840 ( .ip1(n16971), .ip2(n16970), .op(n2067) );
  nand2_1 U17841 ( .ip1(n17229), .ip2(column[46]), .op(n16973) );
  nand2_1 U17842 ( .ip1(\ROUTEDATA/regData [46]), .ip2(n17255), .op(n16972) );
  nand2_1 U17843 ( .ip1(n16973), .ip2(n16972), .op(n2066) );
  nand2_1 U17844 ( .ip1(n17229), .ip2(column[62]), .op(n16975) );
  nand2_1 U17845 ( .ip1(\ROUTEDATA/regData [62]), .ip2(n17258), .op(n16974) );
  nand2_1 U17846 ( .ip1(n16975), .ip2(n16974), .op(n2065) );
  nand2_1 U17847 ( .ip1(n17229), .ip2(column[78]), .op(n16977) );
  nand2_1 U17848 ( .ip1(\ROUTEDATA/regData [78]), .ip2(n17263), .op(n16976) );
  nand2_1 U17849 ( .ip1(n16977), .ip2(n16976), .op(n2064) );
  nand2_1 U17850 ( .ip1(n17229), .ip2(column[94]), .op(n16979) );
  nand2_1 U17851 ( .ip1(\ROUTEDATA/regData [94]), .ip2(n17268), .op(n16978) );
  nand2_1 U17852 ( .ip1(n16979), .ip2(n16978), .op(n2063) );
  nand2_1 U17853 ( .ip1(n17229), .ip2(column[110]), .op(n16981) );
  nand2_1 U17854 ( .ip1(\ROUTEDATA/regData [110]), .ip2(n17273), .op(n16980)
         );
  nand2_1 U17855 ( .ip1(n16981), .ip2(n16980), .op(n2062) );
  nand2_1 U17856 ( .ip1(n17229), .ip2(column[126]), .op(n16983) );
  nand2_1 U17857 ( .ip1(\ROUTEDATA/regData [126]), .ip2(n17278), .op(n16982)
         );
  nand2_1 U17858 ( .ip1(n16983), .ip2(n16982), .op(n2061) );
  nand2_1 U17859 ( .ip1(n17289), .ip2(column[142]), .op(n16985) );
  nand2_1 U17860 ( .ip1(\ROUTEDATA/regData [142]), .ip2(n17285), .op(n16984)
         );
  nand2_1 U17861 ( .ip1(n16985), .ip2(n16984), .op(n2060) );
  nand2_1 U17862 ( .ip1(n17292), .ip2(\ROUTEDATA/regData [158]), .op(n16987)
         );
  nand2_1 U17863 ( .ip1(column[158]), .ip2(n17229), .op(n16986) );
  nand2_1 U17864 ( .ip1(n16987), .ip2(n16986), .op(n2059) );
  nand2_1 U17865 ( .ip1(n17289), .ip2(column[15]), .op(n16989) );
  nand2_1 U17866 ( .ip1(\ROUTEDATA/regData [15]), .ip2(n17244), .op(n16988) );
  nand2_1 U17867 ( .ip1(n16989), .ip2(n16988), .op(n2058) );
  nand2_1 U17868 ( .ip1(n17289), .ip2(column[31]), .op(n16991) );
  nand2_1 U17869 ( .ip1(\ROUTEDATA/regData [31]), .ip2(n17250), .op(n16990) );
  nand2_1 U17870 ( .ip1(n16991), .ip2(n16990), .op(n2057) );
  nand2_1 U17871 ( .ip1(n17289), .ip2(column[47]), .op(n16993) );
  nand2_1 U17872 ( .ip1(\ROUTEDATA/regData [47]), .ip2(n17255), .op(n16992) );
  nand2_1 U17873 ( .ip1(n16993), .ip2(n16992), .op(n2056) );
  nand2_1 U17874 ( .ip1(n17289), .ip2(column[63]), .op(n16995) );
  nand2_1 U17875 ( .ip1(\ROUTEDATA/regData [63]), .ip2(n17258), .op(n16994) );
  nand2_1 U17876 ( .ip1(n16995), .ip2(n16994), .op(n2055) );
  nand2_1 U17877 ( .ip1(n17289), .ip2(column[79]), .op(n16997) );
  nand2_1 U17878 ( .ip1(\ROUTEDATA/regData [79]), .ip2(n17263), .op(n16996) );
  nand2_1 U17879 ( .ip1(n16997), .ip2(n16996), .op(n2054) );
  nand2_1 U17880 ( .ip1(n17289), .ip2(column[95]), .op(n16999) );
  nand2_1 U17881 ( .ip1(\ROUTEDATA/regData [95]), .ip2(n17268), .op(n16998) );
  nand2_1 U17882 ( .ip1(n16999), .ip2(n16998), .op(n2053) );
  nand2_1 U17883 ( .ip1(n17289), .ip2(column[111]), .op(n17001) );
  nand2_1 U17884 ( .ip1(\ROUTEDATA/regData [111]), .ip2(n17273), .op(n17000)
         );
  nand2_1 U17885 ( .ip1(n17001), .ip2(n17000), .op(n2052) );
  nand2_1 U17886 ( .ip1(n17289), .ip2(column[127]), .op(n17003) );
  nand2_1 U17887 ( .ip1(\ROUTEDATA/regData [127]), .ip2(n17278), .op(n17002)
         );
  nand2_1 U17888 ( .ip1(n17003), .ip2(n17002), .op(n2051) );
  nand2_1 U17889 ( .ip1(n17289), .ip2(column[143]), .op(n17005) );
  nand2_1 U17890 ( .ip1(\ROUTEDATA/regData [143]), .ip2(n17285), .op(n17004)
         );
  nand2_1 U17891 ( .ip1(n17005), .ip2(n17004), .op(n2050) );
  nand2_1 U17892 ( .ip1(n17292), .ip2(\ROUTEDATA/regData [159]), .op(n17007)
         );
  nand2_1 U17893 ( .ip1(column[159]), .ip2(n17289), .op(n17006) );
  nand2_1 U17894 ( .ip1(n17007), .ip2(n17006), .op(n2049) );
  nand2_1 U17895 ( .ip1(column[0]), .ip2(n17289), .op(n17010) );
  nand2_1 U17896 ( .ip1(\SIGMOID/N64 ), .ip2(n17241), .op(n17014) );
  inv_1 U17897 ( .ip(n17014), .op(n17035) );
  nand2_1 U17898 ( .ip1(n17243), .ip2(n17035), .op(n17009) );
  nand2_1 U17899 ( .ip1(\ROUTEDATA/regData [0]), .ip2(n17244), .op(n17008) );
  nand3_1 U17900 ( .ip1(n17010), .ip2(n17009), .ip3(n17008), .op(n2048) );
  nand2_1 U17901 ( .ip1(column[16]), .ip2(n17248), .op(n17013) );
  nand2_1 U17902 ( .ip1(n17035), .ip2(n17249), .op(n17012) );
  nand2_1 U17903 ( .ip1(\ROUTEDATA/regData [16]), .ip2(n17250), .op(n17011) );
  nand3_1 U17904 ( .ip1(n17013), .ip2(n17012), .ip3(n17011), .op(n2047) );
  nand2_1 U17905 ( .ip1(n17248), .ip2(column[32]), .op(n17015) );
  nand2_1 U17906 ( .ip1(n17015), .ip2(n17014), .op(n17016) );
  mux2_1 U17907 ( .ip1(n17016), .ip2(\ROUTEDATA/regData [32]), .s(n17255), 
        .op(n2046) );
  nand2_1 U17908 ( .ip1(column[48]), .ip2(n17248), .op(n17019) );
  nand2_1 U17909 ( .ip1(\ROUTEDATA/regData [48]), .ip2(n17258), .op(n17018) );
  nand2_1 U17910 ( .ip1(n17035), .ip2(n17257), .op(n17017) );
  nand3_1 U17911 ( .ip1(n17019), .ip2(n17018), .ip3(n17017), .op(n2045) );
  nand2_1 U17912 ( .ip1(column[64]), .ip2(n17289), .op(n17022) );
  nand2_1 U17913 ( .ip1(n17035), .ip2(n17262), .op(n17021) );
  nand2_1 U17914 ( .ip1(\ROUTEDATA/regData [64]), .ip2(n17263), .op(n17020) );
  nand3_1 U17915 ( .ip1(n17022), .ip2(n17021), .ip3(n17020), .op(n2044) );
  nand2_1 U17916 ( .ip1(column[80]), .ip2(n17289), .op(n17025) );
  nand2_1 U17917 ( .ip1(n17035), .ip2(n17267), .op(n17024) );
  nand2_1 U17918 ( .ip1(\ROUTEDATA/regData [80]), .ip2(n17268), .op(n17023) );
  nand3_1 U17919 ( .ip1(n17025), .ip2(n17024), .ip3(n17023), .op(n2043) );
  nand2_1 U17920 ( .ip1(column[96]), .ip2(n17248), .op(n17028) );
  nand2_1 U17921 ( .ip1(n17035), .ip2(n17272), .op(n17027) );
  nand2_1 U17922 ( .ip1(\ROUTEDATA/regData [96]), .ip2(n17273), .op(n17026) );
  nand3_1 U17923 ( .ip1(n17028), .ip2(n17027), .ip3(n17026), .op(n2042) );
  nand2_1 U17924 ( .ip1(column[112]), .ip2(n17289), .op(n17031) );
  nand2_1 U17925 ( .ip1(n17035), .ip2(n17277), .op(n17030) );
  nand2_1 U17926 ( .ip1(\ROUTEDATA/regData [112]), .ip2(n17278), .op(n17029)
         );
  nand3_1 U17927 ( .ip1(n17031), .ip2(n17030), .ip3(n17029), .op(n2041) );
  nand2_1 U17928 ( .ip1(column[128]), .ip2(n17248), .op(n17034) );
  nand2_1 U17929 ( .ip1(\ROUTEDATA/regData [128]), .ip2(n17285), .op(n17033)
         );
  nand2_1 U17930 ( .ip1(n17035), .ip2(n17283), .op(n17032) );
  nand3_1 U17931 ( .ip1(n17034), .ip2(n17033), .ip3(n17032), .op(n2040) );
  inv_1 U17932 ( .ip(n17292), .op(n17237) );
  nand2_1 U17933 ( .ip1(n17237), .ip2(n17035), .op(n17038) );
  nand2_1 U17934 ( .ip1(n17289), .ip2(column[144]), .op(n17037) );
  nand2_1 U17935 ( .ip1(n17292), .ip2(\ROUTEDATA/regData [144]), .op(n17036)
         );
  nand3_1 U17936 ( .ip1(n17038), .ip2(n17037), .ip3(n17036), .op(n2039) );
  nand2_1 U17937 ( .ip1(column[1]), .ip2(n17248), .op(n17042) );
  and2_1 U17938 ( .ip1(n17241), .ip2(n17039), .op(n17067) );
  nand2_1 U17939 ( .ip1(n17243), .ip2(n17067), .op(n17041) );
  nand2_1 U17940 ( .ip1(\ROUTEDATA/regData [1]), .ip2(n17244), .op(n17040) );
  nand3_1 U17941 ( .ip1(n17042), .ip2(n17041), .ip3(n17040), .op(n2038) );
  nand2_1 U17942 ( .ip1(column[17]), .ip2(n17289), .op(n17045) );
  nand2_1 U17943 ( .ip1(n17067), .ip2(n17249), .op(n17044) );
  nand2_1 U17944 ( .ip1(\ROUTEDATA/regData [17]), .ip2(n17250), .op(n17043) );
  nand3_1 U17945 ( .ip1(n17045), .ip2(n17044), .ip3(n17043), .op(n2037) );
  nand2_1 U17946 ( .ip1(column[33]), .ip2(n17248), .op(n17048) );
  nand2_1 U17947 ( .ip1(n17067), .ip2(n17210), .op(n17047) );
  nand2_1 U17948 ( .ip1(\ROUTEDATA/regData [33]), .ip2(n17255), .op(n17046) );
  nand3_1 U17949 ( .ip1(n17048), .ip2(n17047), .ip3(n17046), .op(n2036) );
  nand2_1 U17950 ( .ip1(column[49]), .ip2(n17289), .op(n17051) );
  nand2_1 U17951 ( .ip1(n17067), .ip2(n17257), .op(n17050) );
  nand2_1 U17952 ( .ip1(\ROUTEDATA/regData [49]), .ip2(n17258), .op(n17049) );
  nand3_1 U17953 ( .ip1(n17051), .ip2(n17050), .ip3(n17049), .op(n2035) );
  nand2_1 U17954 ( .ip1(column[65]), .ip2(n17289), .op(n17054) );
  nand2_1 U17955 ( .ip1(\ROUTEDATA/regData [65]), .ip2(n17263), .op(n17053) );
  nand2_1 U17956 ( .ip1(n17067), .ip2(n17262), .op(n17052) );
  nand3_1 U17957 ( .ip1(n17054), .ip2(n17053), .ip3(n17052), .op(n2034) );
  nand2_1 U17958 ( .ip1(column[81]), .ip2(n17282), .op(n17057) );
  nand2_1 U17959 ( .ip1(\ROUTEDATA/regData [81]), .ip2(n17268), .op(n17056) );
  nand2_1 U17960 ( .ip1(n17067), .ip2(n17267), .op(n17055) );
  nand3_1 U17961 ( .ip1(n17057), .ip2(n17056), .ip3(n17055), .op(n2033) );
  nand2_1 U17962 ( .ip1(column[97]), .ip2(n17248), .op(n17060) );
  nand2_1 U17963 ( .ip1(n17067), .ip2(n17272), .op(n17059) );
  nand2_1 U17964 ( .ip1(\ROUTEDATA/regData [97]), .ip2(n17273), .op(n17058) );
  nand3_1 U17965 ( .ip1(n17060), .ip2(n17059), .ip3(n17058), .op(n2032) );
  nand2_1 U17966 ( .ip1(column[113]), .ip2(n17282), .op(n17063) );
  nand2_1 U17967 ( .ip1(\ROUTEDATA/regData [113]), .ip2(n17278), .op(n17062)
         );
  nand2_1 U17968 ( .ip1(n17067), .ip2(n17277), .op(n17061) );
  nand3_1 U17969 ( .ip1(n17063), .ip2(n17062), .ip3(n17061), .op(n2031) );
  nand2_1 U17970 ( .ip1(column[129]), .ip2(n17248), .op(n17066) );
  nand2_1 U17971 ( .ip1(n17067), .ip2(n17283), .op(n17065) );
  nand2_1 U17972 ( .ip1(\ROUTEDATA/regData [129]), .ip2(n17285), .op(n17064)
         );
  nand3_1 U17973 ( .ip1(n17066), .ip2(n17065), .ip3(n17064), .op(n2030) );
  nand2_1 U17974 ( .ip1(n17237), .ip2(n17067), .op(n17070) );
  nand2_1 U17975 ( .ip1(n17248), .ip2(column[145]), .op(n17069) );
  nand2_1 U17976 ( .ip1(n17292), .ip2(\ROUTEDATA/regData [145]), .op(n17068)
         );
  nand3_1 U17977 ( .ip1(n17070), .ip2(n17069), .ip3(n17068), .op(n2029) );
  nand2_1 U17978 ( .ip1(column[2]), .ip2(n17248), .op(n17075) );
  nand2_1 U17979 ( .ip1(n17241), .ip2(n17071), .op(n17072) );
  inv_1 U17980 ( .ip(n17072), .op(n17100) );
  nand2_1 U17981 ( .ip1(n17243), .ip2(n17100), .op(n17074) );
  nand2_1 U17982 ( .ip1(\ROUTEDATA/regData [2]), .ip2(n17244), .op(n17073) );
  nand3_1 U17983 ( .ip1(n17075), .ip2(n17074), .ip3(n17073), .op(n2028) );
  nand2_1 U17984 ( .ip1(column[18]), .ip2(n17282), .op(n17078) );
  nand2_1 U17985 ( .ip1(n17100), .ip2(n17249), .op(n17077) );
  nand2_1 U17986 ( .ip1(\ROUTEDATA/regData [18]), .ip2(n17250), .op(n17076) );
  nand3_1 U17987 ( .ip1(n17078), .ip2(n17077), .ip3(n17076), .op(n2027) );
  nand2_1 U17988 ( .ip1(column[34]), .ip2(n17282), .op(n17081) );
  nand2_1 U17989 ( .ip1(n17100), .ip2(n17210), .op(n17080) );
  nand2_1 U17990 ( .ip1(\ROUTEDATA/regData [34]), .ip2(n17255), .op(n17079) );
  nand3_1 U17991 ( .ip1(n17081), .ip2(n17080), .ip3(n17079), .op(n2026) );
  nand2_1 U17992 ( .ip1(column[50]), .ip2(n17282), .op(n17084) );
  nand2_1 U17993 ( .ip1(n17100), .ip2(n17257), .op(n17083) );
  nand2_1 U17994 ( .ip1(\ROUTEDATA/regData [50]), .ip2(n17258), .op(n17082) );
  nand3_1 U17995 ( .ip1(n17084), .ip2(n17083), .ip3(n17082), .op(n2025) );
  nand2_1 U17996 ( .ip1(column[66]), .ip2(n17282), .op(n17087) );
  nand2_1 U17997 ( .ip1(n17100), .ip2(n17262), .op(n17086) );
  nand2_1 U17998 ( .ip1(\ROUTEDATA/regData [66]), .ip2(n17263), .op(n17085) );
  nand3_1 U17999 ( .ip1(n17087), .ip2(n17086), .ip3(n17085), .op(n2024) );
  nand2_1 U18000 ( .ip1(column[82]), .ip2(n17282), .op(n17090) );
  nand2_1 U18001 ( .ip1(n17100), .ip2(n17267), .op(n17089) );
  nand2_1 U18002 ( .ip1(\ROUTEDATA/regData [82]), .ip2(n17268), .op(n17088) );
  nand3_1 U18003 ( .ip1(n17090), .ip2(n17089), .ip3(n17088), .op(n2023) );
  nand2_1 U18004 ( .ip1(column[98]), .ip2(n17282), .op(n17093) );
  nand2_1 U18005 ( .ip1(\ROUTEDATA/regData [98]), .ip2(n17273), .op(n17092) );
  nand2_1 U18006 ( .ip1(n17100), .ip2(n17272), .op(n17091) );
  nand3_1 U18007 ( .ip1(n17093), .ip2(n17092), .ip3(n17091), .op(n2022) );
  nand2_1 U18008 ( .ip1(column[114]), .ip2(n17282), .op(n17096) );
  nand2_1 U18009 ( .ip1(n17100), .ip2(n17277), .op(n17095) );
  nand2_1 U18010 ( .ip1(\ROUTEDATA/regData [114]), .ip2(n17278), .op(n17094)
         );
  nand3_1 U18011 ( .ip1(n17096), .ip2(n17095), .ip3(n17094), .op(n2021) );
  nand2_1 U18012 ( .ip1(column[130]), .ip2(n17282), .op(n17099) );
  nand2_1 U18013 ( .ip1(n17100), .ip2(n17283), .op(n17098) );
  nand2_1 U18014 ( .ip1(\ROUTEDATA/regData [130]), .ip2(n17285), .op(n17097)
         );
  nand3_1 U18015 ( .ip1(n17099), .ip2(n17098), .ip3(n17097), .op(n2020) );
  nand2_1 U18016 ( .ip1(n17237), .ip2(n17100), .op(n17103) );
  nand2_1 U18017 ( .ip1(n17248), .ip2(column[146]), .op(n17102) );
  nand2_1 U18018 ( .ip1(n17292), .ip2(\ROUTEDATA/regData [146]), .op(n17101)
         );
  nand3_1 U18019 ( .ip1(n17103), .ip2(n17102), .ip3(n17101), .op(n2019) );
  nand2_1 U18020 ( .ip1(column[3]), .ip2(n17282), .op(n17108) );
  nand2_1 U18021 ( .ip1(n17241), .ip2(n17104), .op(n17105) );
  inv_1 U18022 ( .ip(n17105), .op(n17133) );
  nand2_1 U18023 ( .ip1(n17243), .ip2(n17133), .op(n17107) );
  nand2_1 U18024 ( .ip1(\ROUTEDATA/regData [3]), .ip2(n17244), .op(n17106) );
  nand3_1 U18025 ( .ip1(n17108), .ip2(n17107), .ip3(n17106), .op(n2018) );
  nand2_1 U18026 ( .ip1(column[19]), .ip2(n17282), .op(n17111) );
  nand2_1 U18027 ( .ip1(n17133), .ip2(n17249), .op(n17110) );
  nand2_1 U18028 ( .ip1(\ROUTEDATA/regData [19]), .ip2(n17250), .op(n17109) );
  nand3_1 U18029 ( .ip1(n17111), .ip2(n17110), .ip3(n17109), .op(n2017) );
  nand2_1 U18030 ( .ip1(column[35]), .ip2(n17282), .op(n17114) );
  nand2_1 U18031 ( .ip1(\ROUTEDATA/regData [35]), .ip2(n17255), .op(n17113) );
  nand2_1 U18032 ( .ip1(n17133), .ip2(n17210), .op(n17112) );
  nand3_1 U18033 ( .ip1(n17114), .ip2(n17113), .ip3(n17112), .op(n2016) );
  nand2_1 U18034 ( .ip1(column[51]), .ip2(n17248), .op(n17117) );
  nand2_1 U18035 ( .ip1(n17133), .ip2(n17257), .op(n17116) );
  nand2_1 U18036 ( .ip1(\ROUTEDATA/regData [51]), .ip2(n17258), .op(n17115) );
  nand3_1 U18037 ( .ip1(n17117), .ip2(n17116), .ip3(n17115), .op(n2015) );
  nand2_1 U18038 ( .ip1(column[67]), .ip2(n17282), .op(n17120) );
  nand2_1 U18039 ( .ip1(\ROUTEDATA/regData [67]), .ip2(n17263), .op(n17119) );
  nand2_1 U18040 ( .ip1(n17133), .ip2(n17262), .op(n17118) );
  nand3_1 U18041 ( .ip1(n17120), .ip2(n17119), .ip3(n17118), .op(n2014) );
  nand2_1 U18042 ( .ip1(column[83]), .ip2(n17282), .op(n17123) );
  nand2_1 U18043 ( .ip1(n17133), .ip2(n17267), .op(n17122) );
  nand2_1 U18044 ( .ip1(\ROUTEDATA/regData [83]), .ip2(n17268), .op(n17121) );
  nand3_1 U18045 ( .ip1(n17123), .ip2(n17122), .ip3(n17121), .op(n2013) );
  nand2_1 U18046 ( .ip1(column[99]), .ip2(n17282), .op(n17126) );
  nand2_1 U18047 ( .ip1(n17133), .ip2(n17272), .op(n17125) );
  nand2_1 U18048 ( .ip1(\ROUTEDATA/regData [99]), .ip2(n17273), .op(n17124) );
  nand3_1 U18049 ( .ip1(n17126), .ip2(n17125), .ip3(n17124), .op(n2012) );
  nand2_1 U18050 ( .ip1(column[115]), .ip2(n17282), .op(n17129) );
  nand2_1 U18051 ( .ip1(n17133), .ip2(n17277), .op(n17128) );
  nand2_1 U18052 ( .ip1(\ROUTEDATA/regData [115]), .ip2(n17278), .op(n17127)
         );
  nand3_1 U18053 ( .ip1(n17129), .ip2(n17128), .ip3(n17127), .op(n2011) );
  nand2_1 U18054 ( .ip1(column[131]), .ip2(n17282), .op(n17132) );
  nand2_1 U18055 ( .ip1(\ROUTEDATA/regData [131]), .ip2(n17285), .op(n17131)
         );
  nand2_1 U18056 ( .ip1(n17133), .ip2(n17283), .op(n17130) );
  nand3_1 U18057 ( .ip1(n17132), .ip2(n17131), .ip3(n17130), .op(n2010) );
  nand2_1 U18058 ( .ip1(n17237), .ip2(n17133), .op(n17136) );
  nand2_1 U18059 ( .ip1(n17248), .ip2(column[147]), .op(n17135) );
  nand2_1 U18060 ( .ip1(n17292), .ip2(\ROUTEDATA/regData [147]), .op(n17134)
         );
  nand3_1 U18061 ( .ip1(n17136), .ip2(n17135), .ip3(n17134), .op(n2009) );
  nand2_1 U18062 ( .ip1(column[4]), .ip2(n17282), .op(n17140) );
  nand2_1 U18063 ( .ip1(\ROUTEDATA/regData [4]), .ip2(n17244), .op(n17139) );
  nand2_1 U18064 ( .ip1(n17137), .ip2(n17241), .op(n17166) );
  inv_1 U18065 ( .ip(n17166), .op(n17162) );
  nand2_1 U18066 ( .ip1(n17243), .ip2(n17162), .op(n17138) );
  nand3_1 U18067 ( .ip1(n17140), .ip2(n17139), .ip3(n17138), .op(n2008) );
  nand2_1 U18068 ( .ip1(column[20]), .ip2(n17248), .op(n17143) );
  nand2_1 U18069 ( .ip1(n17162), .ip2(n17249), .op(n17142) );
  nand2_1 U18070 ( .ip1(\ROUTEDATA/regData [20]), .ip2(n17250), .op(n17141) );
  nand3_1 U18071 ( .ip1(n17143), .ip2(n17142), .ip3(n17141), .op(n2007) );
  nand2_1 U18072 ( .ip1(column[36]), .ip2(n17248), .op(n17146) );
  nand2_1 U18073 ( .ip1(n17162), .ip2(n17210), .op(n17145) );
  nand2_1 U18074 ( .ip1(\ROUTEDATA/regData [36]), .ip2(n17255), .op(n17144) );
  nand3_1 U18075 ( .ip1(n17146), .ip2(n17145), .ip3(n17144), .op(n2006) );
  nand2_1 U18076 ( .ip1(column[52]), .ip2(n17282), .op(n17149) );
  nand2_1 U18077 ( .ip1(n17162), .ip2(n17257), .op(n17148) );
  nand2_1 U18078 ( .ip1(\ROUTEDATA/regData [52]), .ip2(n17258), .op(n17147) );
  nand3_1 U18079 ( .ip1(n17149), .ip2(n17148), .ip3(n17147), .op(n2005) );
  nand2_1 U18080 ( .ip1(column[68]), .ip2(n17282), .op(n17152) );
  nand2_1 U18081 ( .ip1(\ROUTEDATA/regData [68]), .ip2(n17263), .op(n17151) );
  nand2_1 U18082 ( .ip1(n17162), .ip2(n17262), .op(n17150) );
  nand3_1 U18083 ( .ip1(n17152), .ip2(n17151), .ip3(n17150), .op(n2004) );
  nand2_1 U18084 ( .ip1(column[84]), .ip2(n17282), .op(n17155) );
  nand2_1 U18085 ( .ip1(\ROUTEDATA/regData [84]), .ip2(n17268), .op(n17154) );
  nand2_1 U18086 ( .ip1(n17162), .ip2(n17267), .op(n17153) );
  nand3_1 U18087 ( .ip1(n17155), .ip2(n17154), .ip3(n17153), .op(n2003) );
  nand2_1 U18088 ( .ip1(column[100]), .ip2(n17248), .op(n17158) );
  nand2_1 U18089 ( .ip1(\ROUTEDATA/regData [100]), .ip2(n17273), .op(n17157)
         );
  nand2_1 U18090 ( .ip1(n17162), .ip2(n17272), .op(n17156) );
  nand3_1 U18091 ( .ip1(n17158), .ip2(n17157), .ip3(n17156), .op(n2002) );
  nand2_1 U18092 ( .ip1(column[116]), .ip2(n17248), .op(n17161) );
  nand2_1 U18093 ( .ip1(n17162), .ip2(n17277), .op(n17160) );
  nand2_1 U18094 ( .ip1(\ROUTEDATA/regData [116]), .ip2(n17278), .op(n17159)
         );
  nand3_1 U18095 ( .ip1(n17161), .ip2(n17160), .ip3(n17159), .op(n2001) );
  nand2_1 U18096 ( .ip1(column[132]), .ip2(n17282), .op(n17165) );
  nand2_1 U18097 ( .ip1(\ROUTEDATA/regData [132]), .ip2(n17285), .op(n17164)
         );
  nand2_1 U18098 ( .ip1(n17162), .ip2(n17283), .op(n17163) );
  nand3_1 U18099 ( .ip1(n17165), .ip2(n17164), .ip3(n17163), .op(n2000) );
  nand2_1 U18100 ( .ip1(n17289), .ip2(column[148]), .op(n17167) );
  nand2_1 U18101 ( .ip1(n17167), .ip2(n17166), .op(n17168) );
  mux2_1 U18102 ( .ip1(n17168), .ip2(\ROUTEDATA/regData [148]), .s(n17292), 
        .op(n1999) );
  nand2_1 U18103 ( .ip1(column[5]), .ip2(n17248), .op(n17172) );
  and2_1 U18104 ( .ip1(n17169), .ip2(n17241), .op(n17197) );
  nand2_1 U18105 ( .ip1(n17243), .ip2(n17197), .op(n17171) );
  nand2_1 U18106 ( .ip1(\ROUTEDATA/regData [5]), .ip2(n17244), .op(n17170) );
  nand3_1 U18107 ( .ip1(n17172), .ip2(n17171), .ip3(n17170), .op(n1998) );
  nand2_1 U18108 ( .ip1(column[21]), .ip2(n17248), .op(n17175) );
  nand2_1 U18109 ( .ip1(n17197), .ip2(n17249), .op(n17174) );
  nand2_1 U18110 ( .ip1(\ROUTEDATA/regData [21]), .ip2(n17250), .op(n17173) );
  nand3_1 U18111 ( .ip1(n17175), .ip2(n17174), .ip3(n17173), .op(n1997) );
  nand2_1 U18112 ( .ip1(column[37]), .ip2(n17248), .op(n17178) );
  nand2_1 U18113 ( .ip1(\ROUTEDATA/regData [37]), .ip2(n17255), .op(n17177) );
  nand2_1 U18114 ( .ip1(n17197), .ip2(n17210), .op(n17176) );
  nand3_1 U18115 ( .ip1(n17178), .ip2(n17177), .ip3(n17176), .op(n1996) );
  nand2_1 U18116 ( .ip1(column[53]), .ip2(n17282), .op(n17181) );
  nand2_1 U18117 ( .ip1(\ROUTEDATA/regData [53]), .ip2(n17258), .op(n17180) );
  nand2_1 U18118 ( .ip1(n17197), .ip2(n17257), .op(n17179) );
  nand3_1 U18119 ( .ip1(n17181), .ip2(n17180), .ip3(n17179), .op(n1995) );
  nand2_1 U18120 ( .ip1(column[69]), .ip2(n17282), .op(n17184) );
  nand2_1 U18121 ( .ip1(\ROUTEDATA/regData [69]), .ip2(n17263), .op(n17183) );
  nand2_1 U18122 ( .ip1(n17197), .ip2(n17262), .op(n17182) );
  nand3_1 U18123 ( .ip1(n17184), .ip2(n17183), .ip3(n17182), .op(n1994) );
  nand2_1 U18124 ( .ip1(column[85]), .ip2(n17248), .op(n17187) );
  nand2_1 U18125 ( .ip1(n17197), .ip2(n17267), .op(n17186) );
  nand2_1 U18126 ( .ip1(\ROUTEDATA/regData [85]), .ip2(n17268), .op(n17185) );
  nand3_1 U18127 ( .ip1(n17187), .ip2(n17186), .ip3(n17185), .op(n1993) );
  nand2_1 U18128 ( .ip1(column[101]), .ip2(n17282), .op(n17190) );
  nand2_1 U18129 ( .ip1(\ROUTEDATA/regData [101]), .ip2(n17273), .op(n17189)
         );
  nand2_1 U18130 ( .ip1(n17197), .ip2(n17272), .op(n17188) );
  nand3_1 U18131 ( .ip1(n17190), .ip2(n17189), .ip3(n17188), .op(n1992) );
  nand2_1 U18132 ( .ip1(column[117]), .ip2(n17282), .op(n17193) );
  nand2_1 U18133 ( .ip1(\ROUTEDATA/regData [117]), .ip2(n17278), .op(n17192)
         );
  nand2_1 U18134 ( .ip1(n17197), .ip2(n17277), .op(n17191) );
  nand3_1 U18135 ( .ip1(n17193), .ip2(n17192), .ip3(n17191), .op(n1991) );
  nand2_1 U18136 ( .ip1(column[133]), .ip2(n17248), .op(n17196) );
  nand2_1 U18137 ( .ip1(\ROUTEDATA/regData [133]), .ip2(n17285), .op(n17195)
         );
  nand2_1 U18138 ( .ip1(n17197), .ip2(n17283), .op(n17194) );
  nand3_1 U18139 ( .ip1(n17196), .ip2(n17195), .ip3(n17194), .op(n1990) );
  nand2_1 U18140 ( .ip1(n17237), .ip2(n17197), .op(n17200) );
  nand2_1 U18141 ( .ip1(n17248), .ip2(column[149]), .op(n17199) );
  nand2_1 U18142 ( .ip1(n17292), .ip2(\ROUTEDATA/regData [149]), .op(n17198)
         );
  nand3_1 U18143 ( .ip1(n17200), .ip2(n17199), .ip3(n17198), .op(n1989) );
  nand2_1 U18144 ( .ip1(column[6]), .ip2(n17248), .op(n17204) );
  nand2_1 U18145 ( .ip1(n17201), .ip2(n17241), .op(n17208) );
  inv_1 U18146 ( .ip(n17208), .op(n17236) );
  nand2_1 U18147 ( .ip1(n17243), .ip2(n17236), .op(n17203) );
  nand2_1 U18148 ( .ip1(\ROUTEDATA/regData [6]), .ip2(n17244), .op(n17202) );
  nand3_1 U18149 ( .ip1(n17204), .ip2(n17203), .ip3(n17202), .op(n1988) );
  nand2_1 U18150 ( .ip1(column[22]), .ip2(n17248), .op(n17207) );
  nand2_1 U18151 ( .ip1(n17236), .ip2(n17249), .op(n17206) );
  nand2_1 U18152 ( .ip1(\ROUTEDATA/regData [22]), .ip2(n17250), .op(n17205) );
  nand3_1 U18153 ( .ip1(n17207), .ip2(n17206), .ip3(n17205), .op(n1987) );
  nand2_1 U18154 ( .ip1(\ROUTEDATA/regData [38]), .ip2(n17255), .op(n17213) );
  nand2_1 U18155 ( .ip1(n17248), .ip2(column[38]), .op(n17209) );
  nand2_1 U18156 ( .ip1(n17209), .ip2(n17208), .op(n17211) );
  nand2_1 U18157 ( .ip1(n17211), .ip2(n17210), .op(n17212) );
  nand2_1 U18158 ( .ip1(n17213), .ip2(n17212), .op(n1986) );
  nand2_1 U18159 ( .ip1(column[54]), .ip2(n17248), .op(n17216) );
  nand2_1 U18160 ( .ip1(n17236), .ip2(n17257), .op(n17215) );
  nand2_1 U18161 ( .ip1(\ROUTEDATA/regData [54]), .ip2(n17258), .op(n17214) );
  nand3_1 U18162 ( .ip1(n17216), .ip2(n17215), .ip3(n17214), .op(n1985) );
  nand2_1 U18163 ( .ip1(column[70]), .ip2(n17248), .op(n17219) );
  nand2_1 U18164 ( .ip1(n17236), .ip2(n17262), .op(n17218) );
  nand2_1 U18165 ( .ip1(\ROUTEDATA/regData [70]), .ip2(n17263), .op(n17217) );
  nand3_1 U18166 ( .ip1(n17219), .ip2(n17218), .ip3(n17217), .op(n1984) );
  nand2_1 U18167 ( .ip1(column[86]), .ip2(n17248), .op(n17222) );
  nand2_1 U18168 ( .ip1(n17236), .ip2(n17267), .op(n17221) );
  nand2_1 U18169 ( .ip1(\ROUTEDATA/regData [86]), .ip2(n17268), .op(n17220) );
  nand3_1 U18170 ( .ip1(n17222), .ip2(n17221), .ip3(n17220), .op(n1983) );
  nand2_1 U18171 ( .ip1(column[102]), .ip2(n17282), .op(n17225) );
  nand2_1 U18172 ( .ip1(n17236), .ip2(n17272), .op(n17224) );
  nand2_1 U18173 ( .ip1(\ROUTEDATA/regData [102]), .ip2(n17273), .op(n17223)
         );
  nand3_1 U18174 ( .ip1(n17225), .ip2(n17224), .ip3(n17223), .op(n1982) );
  nand2_1 U18175 ( .ip1(column[118]), .ip2(n17248), .op(n17228) );
  nand2_1 U18176 ( .ip1(n17236), .ip2(n17277), .op(n17227) );
  nand2_1 U18177 ( .ip1(\ROUTEDATA/regData [118]), .ip2(n17278), .op(n17226)
         );
  nand3_1 U18178 ( .ip1(n17228), .ip2(n17227), .ip3(n17226), .op(n1981) );
  nand2_1 U18179 ( .ip1(\ROUTEDATA/regData [134]), .ip2(n17285), .op(n17235)
         );
  or2_1 U18180 ( .ip1(n17229), .ip2(n17236), .op(n17231) );
  or2_1 U18181 ( .ip1(column[134]), .ip2(n17236), .op(n17230) );
  nand2_1 U18182 ( .ip1(n17231), .ip2(n17230), .op(n17232) );
  or2_1 U18183 ( .ip1(n17233), .ip2(n17232), .op(n17234) );
  nand2_1 U18184 ( .ip1(n17235), .ip2(n17234), .op(n1980) );
  nand2_1 U18185 ( .ip1(n17237), .ip2(n17236), .op(n17240) );
  nand2_1 U18186 ( .ip1(n17248), .ip2(column[150]), .op(n17239) );
  nand2_1 U18187 ( .ip1(n17292), .ip2(\ROUTEDATA/regData [150]), .op(n17238)
         );
  nand3_1 U18188 ( .ip1(n17240), .ip2(n17239), .ip3(n17238), .op(n1979) );
  nand2_1 U18189 ( .ip1(column[7]), .ip2(n17248), .op(n17247) );
  nand2_1 U18190 ( .ip1(n17242), .ip2(n17241), .op(n17290) );
  inv_1 U18191 ( .ip(n17290), .op(n17284) );
  nand2_1 U18192 ( .ip1(n17243), .ip2(n17284), .op(n17246) );
  nand2_1 U18193 ( .ip1(\ROUTEDATA/regData [7]), .ip2(n17244), .op(n17245) );
  nand3_1 U18194 ( .ip1(n17247), .ip2(n17246), .ip3(n17245), .op(n1978) );
  nand2_1 U18195 ( .ip1(column[23]), .ip2(n17248), .op(n17253) );
  nand2_1 U18196 ( .ip1(n17284), .ip2(n17249), .op(n17252) );
  nand2_1 U18197 ( .ip1(\ROUTEDATA/regData [23]), .ip2(n17250), .op(n17251) );
  nand3_1 U18198 ( .ip1(n17253), .ip2(n17252), .ip3(n17251), .op(n1977) );
  nand2_1 U18199 ( .ip1(n17289), .ip2(column[39]), .op(n17254) );
  nand2_1 U18200 ( .ip1(n17254), .ip2(n17290), .op(n17256) );
  mux2_1 U18201 ( .ip1(n17256), .ip2(\ROUTEDATA/regData [39]), .s(n17255), 
        .op(n1976) );
  nand2_1 U18202 ( .ip1(column[55]), .ip2(n17282), .op(n17261) );
  nand2_1 U18203 ( .ip1(n17284), .ip2(n17257), .op(n17260) );
  nand2_1 U18204 ( .ip1(\ROUTEDATA/regData [55]), .ip2(n17258), .op(n17259) );
  nand3_1 U18205 ( .ip1(n17261), .ip2(n17260), .ip3(n17259), .op(n1975) );
  nand2_1 U18206 ( .ip1(column[71]), .ip2(n17282), .op(n17266) );
  nand2_1 U18207 ( .ip1(n17284), .ip2(n17262), .op(n17265) );
  nand2_1 U18208 ( .ip1(\ROUTEDATA/regData [71]), .ip2(n17263), .op(n17264) );
  nand3_1 U18209 ( .ip1(n17266), .ip2(n17265), .ip3(n17264), .op(n1974) );
  nand2_1 U18210 ( .ip1(column[87]), .ip2(n17282), .op(n17271) );
  nand2_1 U18211 ( .ip1(n17284), .ip2(n17267), .op(n17270) );
  nand2_1 U18212 ( .ip1(\ROUTEDATA/regData [87]), .ip2(n17268), .op(n17269) );
  nand3_1 U18213 ( .ip1(n17271), .ip2(n17270), .ip3(n17269), .op(n1973) );
  nand2_1 U18214 ( .ip1(column[103]), .ip2(n17282), .op(n17276) );
  nand2_1 U18215 ( .ip1(n17284), .ip2(n17272), .op(n17275) );
  nand2_1 U18216 ( .ip1(\ROUTEDATA/regData [103]), .ip2(n17273), .op(n17274)
         );
  nand3_1 U18217 ( .ip1(n17276), .ip2(n17275), .ip3(n17274), .op(n1972) );
  nand2_1 U18218 ( .ip1(column[119]), .ip2(n17282), .op(n17281) );
  nand2_1 U18219 ( .ip1(n17284), .ip2(n17277), .op(n17280) );
  nand2_1 U18220 ( .ip1(\ROUTEDATA/regData [119]), .ip2(n17278), .op(n17279)
         );
  nand3_1 U18221 ( .ip1(n17281), .ip2(n17280), .ip3(n17279), .op(n1971) );
  nand2_1 U18222 ( .ip1(column[135]), .ip2(n17282), .op(n17288) );
  nand2_1 U18223 ( .ip1(n17284), .ip2(n17283), .op(n17287) );
  nand2_1 U18224 ( .ip1(\ROUTEDATA/regData [135]), .ip2(n17285), .op(n17286)
         );
  nand3_1 U18225 ( .ip1(n17288), .ip2(n17287), .ip3(n17286), .op(n1970) );
  nand2_1 U18226 ( .ip1(n17289), .ip2(column[151]), .op(n17291) );
  nand2_1 U18227 ( .ip1(n17291), .ip2(n17290), .op(n17293) );
  mux2_1 U18228 ( .ip1(n17293), .ip2(\ROUTEDATA/regData [151]), .s(n17292), 
        .op(n1969) );
  inv_1 U18229 ( .ip(n4362), .op(n17394) );
  mux2_1 U18230 ( .ip1(\ANSWER/mem[0][3][0] ), .ip2(\ANSWER/mem[1][3][0] ), 
        .s(n17394), .op(n17295) );
  mux2_1 U18231 ( .ip1(\ANSWER/mem[2][3][0] ), .ip2(\ANSWER/mem[3][3][0] ), 
        .s(n17394), .op(n17294) );
  inv_1 U18232 ( .ip(n4366), .op(n17366) );
  mux2_1 U18233 ( .ip1(n17295), .ip2(n17294), .s(n17366), .op(n17299) );
  mux2_1 U18234 ( .ip1(\ANSWER/mem[4][3][0] ), .ip2(\ANSWER/mem[5][3][0] ), 
        .s(n17394), .op(n17297) );
  mux2_1 U18235 ( .ip1(\ANSWER/mem[6][3][0] ), .ip2(\ANSWER/mem[7][3][0] ), 
        .s(n17394), .op(n17296) );
  mux2_1 U18236 ( .ip1(n17297), .ip2(n17296), .s(n17366), .op(n17298) );
  mux2_1 U18237 ( .ip1(n17299), .ip2(n17298), .s(n18815), .op(n17301) );
  mux2_1 U18238 ( .ip1(\ANSWER/mem[8][3][0] ), .ip2(\ANSWER/mem[9][3][0] ), 
        .s(n17394), .op(n17300) );
  mux2_1 U18239 ( .ip1(n17301), .ip2(n17300), .s(n18227), .op(n17302) );
  nand2_1 U18240 ( .ip1(n18854), .ip2(n17302), .op(n17376) );
  inv_1 U18241 ( .ip(n4362), .op(n17344) );
  mux2_1 U18242 ( .ip1(\ANSWER/mem[0][0][0] ), .ip2(\ANSWER/mem[1][0][0] ), 
        .s(n17344), .op(n17304) );
  mux2_1 U18243 ( .ip1(\ANSWER/mem[2][0][0] ), .ip2(\ANSWER/mem[3][0][0] ), 
        .s(n17344), .op(n17303) );
  mux2_1 U18244 ( .ip1(n17304), .ip2(n17303), .s(n17366), .op(n17308) );
  mux2_1 U18245 ( .ip1(\ANSWER/mem[4][0][0] ), .ip2(\ANSWER/mem[5][0][0] ), 
        .s(n17344), .op(n17306) );
  mux2_1 U18246 ( .ip1(\ANSWER/mem[6][0][0] ), .ip2(\ANSWER/mem[7][0][0] ), 
        .s(n17344), .op(n17305) );
  mux2_1 U18247 ( .ip1(n17306), .ip2(n17305), .s(n17366), .op(n17307) );
  mux2_1 U18248 ( .ip1(n17308), .ip2(n17307), .s(n18815), .op(n17310) );
  mux2_1 U18249 ( .ip1(\ANSWER/mem[8][0][0] ), .ip2(\ANSWER/mem[9][0][0] ), 
        .s(n17344), .op(n17309) );
  mux2_1 U18250 ( .ip1(n17310), .ip2(n17309), .s(n18227), .op(n17363) );
  buf_1 U18251 ( .ip(n17394), .op(n17387) );
  mux2_1 U18252 ( .ip1(\ANSWER/mem[0][7][0] ), .ip2(\ANSWER/mem[1][7][0] ), 
        .s(n17387), .op(n17312) );
  mux2_1 U18253 ( .ip1(\ANSWER/mem[2][7][0] ), .ip2(\ANSWER/mem[3][7][0] ), 
        .s(n17387), .op(n17311) );
  mux2_1 U18254 ( .ip1(n17312), .ip2(n17311), .s(n18112), .op(n17316) );
  mux2_1 U18255 ( .ip1(\ANSWER/mem[4][7][0] ), .ip2(\ANSWER/mem[5][7][0] ), 
        .s(n17387), .op(n17314) );
  mux2_1 U18256 ( .ip1(\ANSWER/mem[6][7][0] ), .ip2(\ANSWER/mem[7][7][0] ), 
        .s(n17387), .op(n17313) );
  mux2_1 U18257 ( .ip1(n17314), .ip2(n17313), .s(n17794), .op(n17315) );
  mux2_1 U18258 ( .ip1(n17316), .ip2(n17315), .s(n18815), .op(n17318) );
  mux2_1 U18259 ( .ip1(\ANSWER/mem[8][7][0] ), .ip2(\ANSWER/mem[9][7][0] ), 
        .s(n17394), .op(n17317) );
  mux2_1 U18260 ( .ip1(n17318), .ip2(n17317), .s(n18227), .op(n17319) );
  and2_1 U18261 ( .ip1(n18865), .ip2(n17319), .op(n17362) );
  mux2_1 U18262 ( .ip1(\ANSWER/mem[0][4][0] ), .ip2(\ANSWER/mem[1][4][0] ), 
        .s(n17394), .op(n17321) );
  mux2_1 U18263 ( .ip1(\ANSWER/mem[2][4][0] ), .ip2(\ANSWER/mem[3][4][0] ), 
        .s(n17394), .op(n17320) );
  mux2_1 U18264 ( .ip1(n17321), .ip2(n17320), .s(n17366), .op(n17325) );
  mux2_1 U18265 ( .ip1(\ANSWER/mem[4][4][0] ), .ip2(\ANSWER/mem[5][4][0] ), 
        .s(n17394), .op(n17323) );
  mux2_1 U18266 ( .ip1(\ANSWER/mem[6][4][0] ), .ip2(\ANSWER/mem[7][4][0] ), 
        .s(n17394), .op(n17322) );
  mux2_1 U18267 ( .ip1(n17323), .ip2(n17322), .s(n17366), .op(n17324) );
  mux2_1 U18268 ( .ip1(n17325), .ip2(n17324), .s(n18815), .op(n17327) );
  mux2_1 U18269 ( .ip1(\ANSWER/mem[8][4][0] ), .ip2(\ANSWER/mem[9][4][0] ), 
        .s(n17394), .op(n17326) );
  mux2_1 U18270 ( .ip1(n17327), .ip2(n17326), .s(n18227), .op(n17328) );
  nand2_1 U18271 ( .ip1(n18843), .ip2(n17328), .op(n17360) );
  mux2_1 U18272 ( .ip1(\ANSWER/mem[0][2][0] ), .ip2(\ANSWER/mem[1][2][0] ), 
        .s(n17344), .op(n17330) );
  mux2_1 U18273 ( .ip1(\ANSWER/mem[2][2][0] ), .ip2(\ANSWER/mem[3][2][0] ), 
        .s(n17344), .op(n17329) );
  mux2_1 U18274 ( .ip1(n17330), .ip2(n17329), .s(n17366), .op(n17334) );
  mux2_1 U18275 ( .ip1(\ANSWER/mem[4][2][0] ), .ip2(\ANSWER/mem[5][2][0] ), 
        .s(n17344), .op(n17332) );
  mux2_1 U18276 ( .ip1(\ANSWER/mem[6][2][0] ), .ip2(\ANSWER/mem[7][2][0] ), 
        .s(n17394), .op(n17331) );
  mux2_1 U18277 ( .ip1(n17332), .ip2(n17331), .s(n17366), .op(n17333) );
  mux2_1 U18278 ( .ip1(n17334), .ip2(n17333), .s(n18815), .op(n17336) );
  mux2_1 U18279 ( .ip1(\ANSWER/mem[8][2][0] ), .ip2(\ANSWER/mem[9][2][0] ), 
        .s(n17394), .op(n17335) );
  mux2_1 U18280 ( .ip1(n17336), .ip2(n17335), .s(n18227), .op(n17337) );
  nand2_1 U18281 ( .ip1(n18884), .ip2(n17337), .op(n17359) );
  mux2_1 U18282 ( .ip1(\ANSWER/mem[0][1][0] ), .ip2(\ANSWER/mem[1][1][0] ), 
        .s(n17344), .op(n17339) );
  mux2_1 U18283 ( .ip1(\ANSWER/mem[2][1][0] ), .ip2(\ANSWER/mem[3][1][0] ), 
        .s(n17344), .op(n17338) );
  mux2_1 U18284 ( .ip1(n17339), .ip2(n17338), .s(n17366), .op(n17343) );
  mux2_1 U18285 ( .ip1(\ANSWER/mem[4][1][0] ), .ip2(\ANSWER/mem[5][1][0] ), 
        .s(n17344), .op(n17341) );
  mux2_1 U18286 ( .ip1(\ANSWER/mem[6][1][0] ), .ip2(\ANSWER/mem[7][1][0] ), 
        .s(n17344), .op(n17340) );
  mux2_1 U18287 ( .ip1(n17341), .ip2(n17340), .s(n17366), .op(n17342) );
  mux2_1 U18288 ( .ip1(n17343), .ip2(n17342), .s(n18815), .op(n17346) );
  mux2_1 U18289 ( .ip1(\ANSWER/mem[8][1][0] ), .ip2(\ANSWER/mem[9][1][0] ), 
        .s(n17344), .op(n17345) );
  mux2_1 U18290 ( .ip1(n17346), .ip2(n17345), .s(n18227), .op(n17347) );
  nand2_1 U18291 ( .ip1(n18872), .ip2(n17347), .op(n17358) );
  mux2_1 U18292 ( .ip1(\ANSWER/mem[0][6][0] ), .ip2(\ANSWER/mem[1][6][0] ), 
        .s(n17387), .op(n17349) );
  mux2_1 U18293 ( .ip1(\ANSWER/mem[2][6][0] ), .ip2(\ANSWER/mem[3][6][0] ), 
        .s(n17387), .op(n17348) );
  mux2_1 U18294 ( .ip1(n17349), .ip2(n17348), .s(n17366), .op(n17353) );
  mux2_1 U18295 ( .ip1(\ANSWER/mem[4][6][0] ), .ip2(\ANSWER/mem[5][6][0] ), 
        .s(n17387), .op(n17351) );
  mux2_1 U18296 ( .ip1(\ANSWER/mem[6][6][0] ), .ip2(\ANSWER/mem[7][6][0] ), 
        .s(n17387), .op(n17350) );
  mux2_1 U18297 ( .ip1(n17351), .ip2(n17350), .s(n17794), .op(n17352) );
  mux2_1 U18298 ( .ip1(n17353), .ip2(n17352), .s(n18815), .op(n17355) );
  mux2_1 U18299 ( .ip1(\ANSWER/mem[8][6][0] ), .ip2(\ANSWER/mem[9][6][0] ), 
        .s(n17387), .op(n17354) );
  mux2_1 U18300 ( .ip1(n17355), .ip2(n17354), .s(n18227), .op(n17356) );
  nand2_1 U18301 ( .ip1(n18821), .ip2(n17356), .op(n17357) );
  nand4_1 U18302 ( .ip1(n17360), .ip2(n17359), .ip3(n17358), .ip4(n17357), 
        .op(n17361) );
  not_ab_or_c_or_d U18303 ( .ip1(n18800), .ip2(n17363), .ip3(n17362), .ip4(
        n17361), .op(n17375) );
  mux2_1 U18304 ( .ip1(\ANSWER/mem[0][5][0] ), .ip2(\ANSWER/mem[1][5][0] ), 
        .s(n17394), .op(n17365) );
  mux2_1 U18305 ( .ip1(\ANSWER/mem[2][5][0] ), .ip2(\ANSWER/mem[3][5][0] ), 
        .s(n17387), .op(n17364) );
  mux2_1 U18306 ( .ip1(n17365), .ip2(n17364), .s(n17366), .op(n17370) );
  mux2_1 U18307 ( .ip1(\ANSWER/mem[4][5][0] ), .ip2(\ANSWER/mem[5][5][0] ), 
        .s(n17387), .op(n17368) );
  mux2_1 U18308 ( .ip1(\ANSWER/mem[6][5][0] ), .ip2(\ANSWER/mem[7][5][0] ), 
        .s(n17387), .op(n17367) );
  mux2_1 U18309 ( .ip1(n17368), .ip2(n17367), .s(n17366), .op(n17369) );
  mux2_1 U18310 ( .ip1(n17370), .ip2(n17369), .s(n18815), .op(n17372) );
  mux2_1 U18311 ( .ip1(\ANSWER/mem[8][5][0] ), .ip2(\ANSWER/mem[9][5][0] ), 
        .s(n17387), .op(n17371) );
  mux2_1 U18312 ( .ip1(n17372), .ip2(n17371), .s(n18227), .op(n17373) );
  nand2_1 U18313 ( .ip1(n18832), .ip2(n17373), .op(n17374) );
  nand3_1 U18314 ( .ip1(n17376), .ip2(n17375), .ip3(n17374), .op(n17377) );
  nand2_1 U18315 ( .ip1(n17377), .ip2(n18888), .op(n17400) );
  mux2_1 U18316 ( .ip1(\ANSWER/mem[0][8][0] ), .ip2(\ANSWER/mem[1][8][0] ), 
        .s(n17394), .op(n17379) );
  mux2_1 U18317 ( .ip1(\ANSWER/mem[2][8][0] ), .ip2(\ANSWER/mem[3][8][0] ), 
        .s(n17387), .op(n17378) );
  mux2_1 U18318 ( .ip1(n17379), .ip2(n17378), .s(n18138), .op(n17383) );
  mux2_1 U18319 ( .ip1(\ANSWER/mem[4][8][0] ), .ip2(\ANSWER/mem[5][8][0] ), 
        .s(n17394), .op(n17381) );
  mux2_1 U18320 ( .ip1(\ANSWER/mem[6][8][0] ), .ip2(\ANSWER/mem[7][8][0] ), 
        .s(n17394), .op(n17380) );
  mux2_1 U18321 ( .ip1(n17381), .ip2(n17380), .s(n17794), .op(n17382) );
  mux2_1 U18322 ( .ip1(n17383), .ip2(n17382), .s(n18815), .op(n17385) );
  mux2_1 U18323 ( .ip1(\ANSWER/mem[8][8][0] ), .ip2(\ANSWER/mem[9][8][0] ), 
        .s(n17394), .op(n17384) );
  mux2_1 U18324 ( .ip1(n17385), .ip2(n17384), .s(n18227), .op(n17386) );
  nand2_1 U18325 ( .ip1(n18914), .ip2(n17386), .op(n17399) );
  mux2_1 U18326 ( .ip1(\ANSWER/mem[0][9][0] ), .ip2(\ANSWER/mem[1][9][0] ), 
        .s(n17387), .op(n17389) );
  mux2_1 U18327 ( .ip1(\ANSWER/mem[2][9][0] ), .ip2(\ANSWER/mem[3][9][0] ), 
        .s(n17387), .op(n17388) );
  mux2_1 U18328 ( .ip1(n17389), .ip2(n17388), .s(n17688), .op(n17393) );
  mux2_1 U18329 ( .ip1(\ANSWER/mem[4][9][0] ), .ip2(\ANSWER/mem[5][9][0] ), 
        .s(n17394), .op(n17391) );
  mux2_1 U18330 ( .ip1(\ANSWER/mem[6][9][0] ), .ip2(\ANSWER/mem[7][9][0] ), 
        .s(n17394), .op(n17390) );
  mux2_1 U18331 ( .ip1(n17391), .ip2(n17390), .s(n4456), .op(n17392) );
  mux2_1 U18332 ( .ip1(n17393), .ip2(n17392), .s(n18815), .op(n17396) );
  mux2_1 U18333 ( .ip1(\ANSWER/mem[8][9][0] ), .ip2(\ANSWER/mem[9][9][0] ), 
        .s(n17394), .op(n17395) );
  mux2_1 U18334 ( .ip1(n17396), .ip2(n17395), .s(n18227), .op(n17397) );
  nand2_1 U18335 ( .ip1(n18899), .ip2(n17397), .op(n17398) );
  nand3_1 U18336 ( .ip1(n17400), .ip2(n17399), .ip3(n17398), .op(\ANSWER/N487 ) );
  buf_1 U18337 ( .ip(n17401), .op(n17533) );
  mux2_1 U18338 ( .ip1(\ANSWER/mem[0][0][2] ), .ip2(\ANSWER/mem[1][0][2] ), 
        .s(n17533), .op(n17403) );
  mux2_1 U18339 ( .ip1(\ANSWER/mem[2][0][2] ), .ip2(\ANSWER/mem[3][0][2] ), 
        .s(n17533), .op(n17402) );
  mux2_1 U18340 ( .ip1(n17403), .ip2(n17402), .s(n18112), .op(n17407) );
  mux2_1 U18341 ( .ip1(\ANSWER/mem[4][0][2] ), .ip2(\ANSWER/mem[5][0][2] ), 
        .s(n17533), .op(n17405) );
  mux2_1 U18342 ( .ip1(\ANSWER/mem[6][0][2] ), .ip2(\ANSWER/mem[7][0][2] ), 
        .s(n17533), .op(n17404) );
  mux2_1 U18343 ( .ip1(n17405), .ip2(n17404), .s(n18544), .op(n17406) );
  mux2_1 U18344 ( .ip1(n17407), .ip2(n17406), .s(n18906), .op(n17409) );
  mux2_1 U18345 ( .ip1(\ANSWER/mem[8][0][2] ), .ip2(\ANSWER/mem[9][0][2] ), 
        .s(n17533), .op(n17408) );
  mux2_1 U18346 ( .ip1(n17409), .ip2(n17408), .s(n18092), .op(n17410) );
  nand2_1 U18347 ( .ip1(n17410), .ip2(n18800), .op(n17482) );
  mux2_1 U18348 ( .ip1(\ANSWER/mem[0][6][2] ), .ip2(\ANSWER/mem[1][6][2] ), 
        .s(n17506), .op(n17412) );
  mux2_1 U18349 ( .ip1(\ANSWER/mem[2][6][2] ), .ip2(\ANSWER/mem[3][6][2] ), 
        .s(n17564), .op(n17411) );
  mux2_1 U18350 ( .ip1(n17412), .ip2(n17411), .s(n18354), .op(n17416) );
  mux2_1 U18351 ( .ip1(\ANSWER/mem[4][6][2] ), .ip2(\ANSWER/mem[5][6][2] ), 
        .s(n17506), .op(n17414) );
  mux2_1 U18352 ( .ip1(\ANSWER/mem[6][6][2] ), .ip2(\ANSWER/mem[7][6][2] ), 
        .s(n17506), .op(n17413) );
  mux2_1 U18353 ( .ip1(n17414), .ip2(n17413), .s(n15636), .op(n17415) );
  buf_1 U18354 ( .ip(n18859), .op(n18826) );
  mux2_1 U18355 ( .ip1(n17416), .ip2(n17415), .s(n18826), .op(n17418) );
  mux2_1 U18356 ( .ip1(\ANSWER/mem[8][6][2] ), .ip2(\ANSWER/mem[9][6][2] ), 
        .s(n17506), .op(n17417) );
  mux2_1 U18357 ( .ip1(n17418), .ip2(n17417), .s(n18252), .op(n17470) );
  mux2_1 U18358 ( .ip1(\ANSWER/mem[0][7][2] ), .ip2(\ANSWER/mem[1][7][2] ), 
        .s(n17506), .op(n17420) );
  mux2_1 U18359 ( .ip1(\ANSWER/mem[2][7][2] ), .ip2(\ANSWER/mem[3][7][2] ), 
        .s(n17506), .op(n17419) );
  mux2_1 U18360 ( .ip1(n17420), .ip2(n17419), .s(n17688), .op(n17424) );
  mux2_1 U18361 ( .ip1(\ANSWER/mem[4][7][2] ), .ip2(\ANSWER/mem[5][7][2] ), 
        .s(n17506), .op(n17422) );
  mux2_1 U18362 ( .ip1(\ANSWER/mem[6][7][2] ), .ip2(\ANSWER/mem[7][7][2] ), 
        .s(n17506), .op(n17421) );
  mux2_1 U18363 ( .ip1(n17422), .ip2(n17421), .s(n17605), .op(n17423) );
  mux2_1 U18364 ( .ip1(n17424), .ip2(n17423), .s(n18837), .op(n17426) );
  mux2_1 U18365 ( .ip1(\ANSWER/mem[8][7][2] ), .ip2(\ANSWER/mem[9][7][2] ), 
        .s(n17564), .op(n17425) );
  mux2_1 U18366 ( .ip1(n17426), .ip2(n17425), .s(n18252), .op(n17427) );
  and2_1 U18367 ( .ip1(n18865), .ip2(n17427), .op(n17469) );
  mux2_1 U18368 ( .ip1(\ANSWER/mem[0][3][2] ), .ip2(\ANSWER/mem[1][3][2] ), 
        .s(n17506), .op(n17429) );
  mux2_1 U18369 ( .ip1(\ANSWER/mem[2][3][2] ), .ip2(\ANSWER/mem[3][3][2] ), 
        .s(n17506), .op(n17428) );
  mux2_1 U18370 ( .ip1(n17429), .ip2(n17428), .s(n17581), .op(n17433) );
  mux2_1 U18371 ( .ip1(\ANSWER/mem[4][3][2] ), .ip2(\ANSWER/mem[5][3][2] ), 
        .s(n17506), .op(n17431) );
  mux2_1 U18372 ( .ip1(\ANSWER/mem[6][3][2] ), .ip2(\ANSWER/mem[7][3][2] ), 
        .s(n17506), .op(n17430) );
  mux2_1 U18373 ( .ip1(n17431), .ip2(n17430), .s(n17366), .op(n17432) );
  mux2_1 U18374 ( .ip1(n17433), .ip2(n17432), .s(n18815), .op(n17435) );
  mux2_1 U18375 ( .ip1(\ANSWER/mem[8][3][2] ), .ip2(\ANSWER/mem[9][3][2] ), 
        .s(n17506), .op(n17434) );
  mux2_1 U18376 ( .ip1(n17435), .ip2(n17434), .s(n18252), .op(n17436) );
  nand2_1 U18377 ( .ip1(n18854), .ip2(n17436), .op(n17467) );
  mux2_1 U18378 ( .ip1(\ANSWER/mem[0][5][2] ), .ip2(\ANSWER/mem[1][5][2] ), 
        .s(n17564), .op(n17438) );
  mux2_1 U18379 ( .ip1(\ANSWER/mem[2][5][2] ), .ip2(\ANSWER/mem[3][5][2] ), 
        .s(n17506), .op(n17437) );
  mux2_1 U18380 ( .ip1(n17438), .ip2(n17437), .s(n17990), .op(n17442) );
  mux2_1 U18381 ( .ip1(\ANSWER/mem[4][5][2] ), .ip2(\ANSWER/mem[5][5][2] ), 
        .s(n17506), .op(n17440) );
  mux2_1 U18382 ( .ip1(\ANSWER/mem[6][5][2] ), .ip2(\ANSWER/mem[7][5][2] ), 
        .s(n17506), .op(n17439) );
  mux2_1 U18383 ( .ip1(n17440), .ip2(n17439), .s(n17794), .op(n17441) );
  buf_1 U18384 ( .ip(n18878), .op(n18848) );
  mux2_1 U18385 ( .ip1(n17442), .ip2(n17441), .s(n18848), .op(n17444) );
  mux2_1 U18386 ( .ip1(\ANSWER/mem[8][5][2] ), .ip2(\ANSWER/mem[9][5][2] ), 
        .s(n17506), .op(n17443) );
  mux2_1 U18387 ( .ip1(n17444), .ip2(n17443), .s(n18252), .op(n17445) );
  nand2_1 U18388 ( .ip1(n18832), .ip2(n17445), .op(n17466) );
  mux2_1 U18389 ( .ip1(\ANSWER/mem[0][1][2] ), .ip2(\ANSWER/mem[1][1][2] ), 
        .s(n17533), .op(n17447) );
  mux2_1 U18390 ( .ip1(\ANSWER/mem[2][1][2] ), .ip2(\ANSWER/mem[3][1][2] ), 
        .s(n17533), .op(n17446) );
  mux2_1 U18391 ( .ip1(n17447), .ip2(n17446), .s(n17688), .op(n17451) );
  mux2_1 U18392 ( .ip1(\ANSWER/mem[4][1][2] ), .ip2(\ANSWER/mem[5][1][2] ), 
        .s(n17533), .op(n17449) );
  mux2_1 U18393 ( .ip1(\ANSWER/mem[6][1][2] ), .ip2(\ANSWER/mem[7][1][2] ), 
        .s(n17533), .op(n17448) );
  mux2_1 U18394 ( .ip1(n17449), .ip2(n17448), .s(n17605), .op(n17450) );
  buf_1 U18395 ( .ip(n18878), .op(n18806) );
  mux2_1 U18396 ( .ip1(n17451), .ip2(n17450), .s(n18806), .op(n17453) );
  mux2_1 U18397 ( .ip1(\ANSWER/mem[8][1][2] ), .ip2(\ANSWER/mem[9][1][2] ), 
        .s(n17533), .op(n17452) );
  mux2_1 U18398 ( .ip1(n17453), .ip2(n17452), .s(n18252), .op(n17454) );
  nand2_1 U18399 ( .ip1(n18872), .ip2(n17454), .op(n17465) );
  mux2_1 U18400 ( .ip1(\ANSWER/mem[0][2][2] ), .ip2(\ANSWER/mem[1][2][2] ), 
        .s(n17533), .op(n17456) );
  mux2_1 U18401 ( .ip1(\ANSWER/mem[2][2][2] ), .ip2(\ANSWER/mem[3][2][2] ), 
        .s(n17533), .op(n17455) );
  mux2_1 U18402 ( .ip1(n17456), .ip2(n17455), .s(n17581), .op(n17460) );
  mux2_1 U18403 ( .ip1(\ANSWER/mem[4][2][2] ), .ip2(\ANSWER/mem[5][2][2] ), 
        .s(n17533), .op(n17458) );
  mux2_1 U18404 ( .ip1(\ANSWER/mem[6][2][2] ), .ip2(\ANSWER/mem[7][2][2] ), 
        .s(n17506), .op(n17457) );
  mux2_1 U18405 ( .ip1(n17458), .ip2(n17457), .s(n4456), .op(n17459) );
  mux2_1 U18406 ( .ip1(n17460), .ip2(n17459), .s(n18848), .op(n17462) );
  mux2_1 U18407 ( .ip1(\ANSWER/mem[8][2][2] ), .ip2(\ANSWER/mem[9][2][2] ), 
        .s(n17506), .op(n17461) );
  mux2_1 U18408 ( .ip1(n17462), .ip2(n17461), .s(n18252), .op(n17463) );
  nand2_1 U18409 ( .ip1(n18884), .ip2(n17463), .op(n17464) );
  nand4_1 U18410 ( .ip1(n17467), .ip2(n17466), .ip3(n17465), .ip4(n17464), 
        .op(n17468) );
  not_ab_or_c_or_d U18411 ( .ip1(n17470), .ip2(n18821), .ip3(n17469), .ip4(
        n17468), .op(n17481) );
  mux2_1 U18412 ( .ip1(\ANSWER/mem[0][4][2] ), .ip2(\ANSWER/mem[1][4][2] ), 
        .s(n17506), .op(n17472) );
  mux2_1 U18413 ( .ip1(\ANSWER/mem[2][4][2] ), .ip2(\ANSWER/mem[3][4][2] ), 
        .s(n17506), .op(n17471) );
  mux2_1 U18414 ( .ip1(n17472), .ip2(n17471), .s(n18138), .op(n17476) );
  mux2_1 U18415 ( .ip1(\ANSWER/mem[4][4][2] ), .ip2(\ANSWER/mem[5][4][2] ), 
        .s(n17564), .op(n17474) );
  mux2_1 U18416 ( .ip1(\ANSWER/mem[6][4][2] ), .ip2(\ANSWER/mem[7][4][2] ), 
        .s(n17564), .op(n17473) );
  mux2_1 U18417 ( .ip1(n17474), .ip2(n17473), .s(n18330), .op(n17475) );
  buf_1 U18418 ( .ip(n18859), .op(n18906) );
  mux2_1 U18419 ( .ip1(n17476), .ip2(n17475), .s(n18906), .op(n17478) );
  mux2_1 U18420 ( .ip1(\ANSWER/mem[8][4][2] ), .ip2(\ANSWER/mem[9][4][2] ), 
        .s(n17564), .op(n17477) );
  mux2_1 U18421 ( .ip1(n17478), .ip2(n17477), .s(n18252), .op(n17479) );
  nand2_1 U18422 ( .ip1(n18843), .ip2(n17479), .op(n17480) );
  nand3_1 U18423 ( .ip1(n17482), .ip2(n17481), .ip3(n17480), .op(n17483) );
  nand2_1 U18424 ( .ip1(n17483), .ip2(n18888), .op(n17505) );
  mux2_1 U18425 ( .ip1(\ANSWER/mem[0][8][2] ), .ip2(\ANSWER/mem[1][8][2] ), 
        .s(n17564), .op(n17485) );
  mux2_1 U18426 ( .ip1(\ANSWER/mem[2][8][2] ), .ip2(\ANSWER/mem[3][8][2] ), 
        .s(n17564), .op(n17484) );
  mux2_1 U18427 ( .ip1(n17485), .ip2(n17484), .s(n17605), .op(n17490) );
  mux2_1 U18428 ( .ip1(\ANSWER/mem[4][8][2] ), .ip2(\ANSWER/mem[5][8][2] ), 
        .s(n17564), .op(n17487) );
  mux2_1 U18429 ( .ip1(\ANSWER/mem[6][8][2] ), .ip2(\ANSWER/mem[7][8][2] ), 
        .s(n17564), .op(n17486) );
  mux2_1 U18430 ( .ip1(n17487), .ip2(n17486), .s(n18354), .op(n17489) );
  mux2_1 U18431 ( .ip1(n17490), .ip2(n17489), .s(n18826), .op(n17492) );
  mux2_1 U18432 ( .ip1(\ANSWER/mem[8][8][2] ), .ip2(\ANSWER/mem[9][8][2] ), 
        .s(n17564), .op(n17491) );
  mux2_1 U18433 ( .ip1(n17492), .ip2(n17491), .s(n18092), .op(n17493) );
  nand2_1 U18434 ( .ip1(n18914), .ip2(n17493), .op(n17504) );
  mux2_1 U18435 ( .ip1(\ANSWER/mem[0][9][2] ), .ip2(\ANSWER/mem[1][9][2] ), 
        .s(n17564), .op(n17495) );
  mux2_1 U18436 ( .ip1(\ANSWER/mem[2][9][2] ), .ip2(\ANSWER/mem[3][9][2] ), 
        .s(n17564), .op(n17494) );
  mux2_1 U18437 ( .ip1(n17495), .ip2(n17494), .s(n17366), .op(n17499) );
  mux2_1 U18438 ( .ip1(\ANSWER/mem[4][9][2] ), .ip2(\ANSWER/mem[5][9][2] ), 
        .s(n17564), .op(n17497) );
  mux2_1 U18439 ( .ip1(\ANSWER/mem[6][9][2] ), .ip2(\ANSWER/mem[7][9][2] ), 
        .s(n17564), .op(n17496) );
  mux2_1 U18440 ( .ip1(n17497), .ip2(n17496), .s(n18544), .op(n17498) );
  mux2_1 U18441 ( .ip1(n17499), .ip2(n17498), .s(n18878), .op(n17501) );
  mux2_1 U18442 ( .ip1(\ANSWER/mem[8][9][2] ), .ip2(\ANSWER/mem[9][9][2] ), 
        .s(n17564), .op(n17500) );
  mux2_1 U18443 ( .ip1(n17501), .ip2(n17500), .s(n18092), .op(n17502) );
  nand2_1 U18444 ( .ip1(n18899), .ip2(n17502), .op(n17503) );
  nand3_1 U18445 ( .ip1(n17505), .ip2(n17504), .ip3(n17503), .op(\ANSWER/N485 ) );
  buf_1 U18446 ( .ip(n17506), .op(n17602) );
  mux2_1 U18447 ( .ip1(\ANSWER/mem[0][0][3] ), .ip2(\ANSWER/mem[1][0][3] ), 
        .s(n17602), .op(n17508) );
  mux2_1 U18448 ( .ip1(\ANSWER/mem[2][0][3] ), .ip2(\ANSWER/mem[3][0][3] ), 
        .s(n17602), .op(n17507) );
  inv_1 U18449 ( .ip(n4366), .op(n17581) );
  mux2_1 U18450 ( .ip1(n17508), .ip2(n17507), .s(n17581), .op(n17512) );
  mux2_1 U18451 ( .ip1(\ANSWER/mem[4][0][3] ), .ip2(\ANSWER/mem[5][0][3] ), 
        .s(n17602), .op(n17510) );
  mux2_1 U18452 ( .ip1(\ANSWER/mem[6][0][3] ), .ip2(\ANSWER/mem[7][0][3] ), 
        .s(n17602), .op(n17509) );
  mux2_1 U18453 ( .ip1(n17510), .ip2(n17509), .s(n17581), .op(n17511) );
  mux2_1 U18454 ( .ip1(n17512), .ip2(n17511), .s(n18806), .op(n17514) );
  mux2_1 U18455 ( .ip1(\ANSWER/mem[8][0][3] ), .ip2(\ANSWER/mem[9][0][3] ), 
        .s(n17602), .op(n17513) );
  mux2_1 U18456 ( .ip1(n17514), .ip2(n17513), .s(n18252), .op(n17515) );
  nand2_1 U18457 ( .ip1(n17515), .ip2(n18800), .op(n17591) );
  mux2_1 U18458 ( .ip1(\ANSWER/mem[0][1][3] ), .ip2(\ANSWER/mem[1][1][3] ), 
        .s(n17536), .op(n17517) );
  mux2_1 U18459 ( .ip1(\ANSWER/mem[2][1][3] ), .ip2(\ANSWER/mem[3][1][3] ), 
        .s(n17536), .op(n17516) );
  mux2_1 U18460 ( .ip1(n17517), .ip2(n17516), .s(n17581), .op(n17521) );
  mux2_1 U18461 ( .ip1(\ANSWER/mem[4][1][3] ), .ip2(\ANSWER/mem[5][1][3] ), 
        .s(n17533), .op(n17519) );
  mux2_1 U18462 ( .ip1(\ANSWER/mem[6][1][3] ), .ip2(\ANSWER/mem[7][1][3] ), 
        .s(n17536), .op(n17518) );
  mux2_1 U18463 ( .ip1(n17519), .ip2(n17518), .s(n17581), .op(n17520) );
  mux2_1 U18464 ( .ip1(n17521), .ip2(n17520), .s(n18848), .op(n17523) );
  mux2_1 U18465 ( .ip1(\ANSWER/mem[8][1][3] ), .ip2(\ANSWER/mem[9][1][3] ), 
        .s(n17602), .op(n17522) );
  mux2_1 U18466 ( .ip1(n17523), .ip2(n17522), .s(n18252), .op(n17578) );
  mux2_1 U18467 ( .ip1(\ANSWER/mem[0][7][3] ), .ip2(\ANSWER/mem[1][7][3] ), 
        .s(n17610), .op(n17525) );
  mux2_1 U18468 ( .ip1(\ANSWER/mem[2][7][3] ), .ip2(\ANSWER/mem[3][7][3] ), 
        .s(n17610), .op(n17524) );
  inv_1 U18469 ( .ip(n4366), .op(n17605) );
  mux2_1 U18470 ( .ip1(n17525), .ip2(n17524), .s(n17605), .op(n17529) );
  mux2_1 U18471 ( .ip1(\ANSWER/mem[4][7][3] ), .ip2(\ANSWER/mem[5][7][3] ), 
        .s(n17610), .op(n17527) );
  mux2_1 U18472 ( .ip1(\ANSWER/mem[6][7][3] ), .ip2(\ANSWER/mem[7][7][3] ), 
        .s(n17610), .op(n17526) );
  mux2_1 U18473 ( .ip1(n17527), .ip2(n17526), .s(n17605), .op(n17528) );
  mux2_1 U18474 ( .ip1(n17529), .ip2(n17528), .s(n18859), .op(n17531) );
  mux2_1 U18475 ( .ip1(\ANSWER/mem[8][7][3] ), .ip2(\ANSWER/mem[9][7][3] ), 
        .s(n17610), .op(n17530) );
  mux2_1 U18476 ( .ip1(n17531), .ip2(n17530), .s(n18252), .op(n17532) );
  and2_1 U18477 ( .ip1(n18865), .ip2(n17532), .op(n17577) );
  mux2_1 U18478 ( .ip1(\ANSWER/mem[0][2][3] ), .ip2(\ANSWER/mem[1][2][3] ), 
        .s(n17533), .op(n17535) );
  mux2_1 U18479 ( .ip1(\ANSWER/mem[2][2][3] ), .ip2(\ANSWER/mem[3][2][3] ), 
        .s(n17533), .op(n17534) );
  mux2_1 U18480 ( .ip1(n17535), .ip2(n17534), .s(n17581), .op(n17540) );
  mux2_1 U18481 ( .ip1(\ANSWER/mem[4][2][3] ), .ip2(\ANSWER/mem[5][2][3] ), 
        .s(n17536), .op(n17538) );
  mux2_1 U18482 ( .ip1(\ANSWER/mem[6][2][3] ), .ip2(\ANSWER/mem[7][2][3] ), 
        .s(n17602), .op(n17537) );
  mux2_1 U18483 ( .ip1(n17538), .ip2(n17537), .s(n17581), .op(n17539) );
  mux2_1 U18484 ( .ip1(n17540), .ip2(n17539), .s(n18815), .op(n17542) );
  mux2_1 U18485 ( .ip1(\ANSWER/mem[8][2][3] ), .ip2(\ANSWER/mem[9][2][3] ), 
        .s(n17602), .op(n17541) );
  mux2_1 U18486 ( .ip1(n17542), .ip2(n17541), .s(n18252), .op(n17543) );
  nand2_1 U18487 ( .ip1(n18884), .ip2(n17543), .op(n17575) );
  mux2_1 U18488 ( .ip1(\ANSWER/mem[0][3][3] ), .ip2(\ANSWER/mem[1][3][3] ), 
        .s(n17602), .op(n17545) );
  mux2_1 U18489 ( .ip1(\ANSWER/mem[2][3][3] ), .ip2(\ANSWER/mem[3][3][3] ), 
        .s(n17602), .op(n17544) );
  mux2_1 U18490 ( .ip1(n17545), .ip2(n17544), .s(n17581), .op(n17549) );
  mux2_1 U18491 ( .ip1(\ANSWER/mem[4][3][3] ), .ip2(\ANSWER/mem[5][3][3] ), 
        .s(n17602), .op(n17547) );
  mux2_1 U18492 ( .ip1(\ANSWER/mem[6][3][3] ), .ip2(\ANSWER/mem[7][3][3] ), 
        .s(n17602), .op(n17546) );
  mux2_1 U18493 ( .ip1(n17547), .ip2(n17546), .s(n17581), .op(n17548) );
  mux2_1 U18494 ( .ip1(n17549), .ip2(n17548), .s(n18859), .op(n17551) );
  mux2_1 U18495 ( .ip1(\ANSWER/mem[8][3][3] ), .ip2(\ANSWER/mem[9][3][3] ), 
        .s(n17602), .op(n17550) );
  mux2_1 U18496 ( .ip1(n17551), .ip2(n17550), .s(n18252), .op(n17552) );
  nand2_1 U18497 ( .ip1(n18854), .ip2(n17552), .op(n17574) );
  mux2_1 U18498 ( .ip1(\ANSWER/mem[0][6][3] ), .ip2(\ANSWER/mem[1][6][3] ), 
        .s(n17564), .op(n17554) );
  mux2_1 U18499 ( .ip1(\ANSWER/mem[2][6][3] ), .ip2(\ANSWER/mem[3][6][3] ), 
        .s(n17610), .op(n17553) );
  mux2_1 U18500 ( .ip1(n17554), .ip2(n17553), .s(n17581), .op(n17558) );
  mux2_1 U18501 ( .ip1(\ANSWER/mem[4][6][3] ), .ip2(\ANSWER/mem[5][6][3] ), 
        .s(n17610), .op(n17556) );
  mux2_1 U18502 ( .ip1(\ANSWER/mem[6][6][3] ), .ip2(\ANSWER/mem[7][6][3] ), 
        .s(n17610), .op(n17555) );
  mux2_1 U18503 ( .ip1(n17556), .ip2(n17555), .s(n17605), .op(n17557) );
  mux2_1 U18504 ( .ip1(n17558), .ip2(n17557), .s(n18859), .op(n17560) );
  mux2_1 U18505 ( .ip1(\ANSWER/mem[8][6][3] ), .ip2(\ANSWER/mem[9][6][3] ), 
        .s(n17610), .op(n17559) );
  mux2_1 U18506 ( .ip1(n17560), .ip2(n17559), .s(n18252), .op(n17561) );
  nand2_1 U18507 ( .ip1(n18821), .ip2(n17561), .op(n17573) );
  mux2_1 U18508 ( .ip1(\ANSWER/mem[0][5][3] ), .ip2(\ANSWER/mem[1][5][3] ), 
        .s(n17602), .op(n17563) );
  mux2_1 U18509 ( .ip1(\ANSWER/mem[2][5][3] ), .ip2(\ANSWER/mem[3][5][3] ), 
        .s(n17610), .op(n17562) );
  mux2_1 U18510 ( .ip1(n17563), .ip2(n17562), .s(n17581), .op(n17568) );
  mux2_1 U18511 ( .ip1(\ANSWER/mem[4][5][3] ), .ip2(\ANSWER/mem[5][5][3] ), 
        .s(n17564), .op(n17566) );
  mux2_1 U18512 ( .ip1(\ANSWER/mem[6][5][3] ), .ip2(\ANSWER/mem[7][5][3] ), 
        .s(n17610), .op(n17565) );
  mux2_1 U18513 ( .ip1(n17566), .ip2(n17565), .s(n17581), .op(n17567) );
  mux2_1 U18514 ( .ip1(n17568), .ip2(n17567), .s(n18837), .op(n17570) );
  mux2_1 U18515 ( .ip1(\ANSWER/mem[8][5][3] ), .ip2(\ANSWER/mem[9][5][3] ), 
        .s(n17610), .op(n17569) );
  mux2_1 U18516 ( .ip1(n17570), .ip2(n17569), .s(n18252), .op(n17571) );
  nand2_1 U18517 ( .ip1(n18832), .ip2(n17571), .op(n17572) );
  nand4_1 U18518 ( .ip1(n17575), .ip2(n17574), .ip3(n17573), .ip4(n17572), 
        .op(n17576) );
  not_ab_or_c_or_d U18519 ( .ip1(n18872), .ip2(n17578), .ip3(n17577), .ip4(
        n17576), .op(n17590) );
  mux2_1 U18520 ( .ip1(\ANSWER/mem[0][4][3] ), .ip2(\ANSWER/mem[1][4][3] ), 
        .s(n17602), .op(n17580) );
  mux2_1 U18521 ( .ip1(\ANSWER/mem[2][4][3] ), .ip2(\ANSWER/mem[3][4][3] ), 
        .s(n17602), .op(n17579) );
  mux2_1 U18522 ( .ip1(n17580), .ip2(n17579), .s(n17581), .op(n17585) );
  mux2_1 U18523 ( .ip1(\ANSWER/mem[4][4][3] ), .ip2(\ANSWER/mem[5][4][3] ), 
        .s(n17602), .op(n17583) );
  mux2_1 U18524 ( .ip1(\ANSWER/mem[6][4][3] ), .ip2(\ANSWER/mem[7][4][3] ), 
        .s(n17602), .op(n17582) );
  mux2_1 U18525 ( .ip1(n17583), .ip2(n17582), .s(n17581), .op(n17584) );
  mux2_1 U18526 ( .ip1(n17585), .ip2(n17584), .s(n18837), .op(n17587) );
  mux2_1 U18527 ( .ip1(\ANSWER/mem[8][4][3] ), .ip2(\ANSWER/mem[9][4][3] ), 
        .s(n17602), .op(n17586) );
  mux2_1 U18528 ( .ip1(n17587), .ip2(n17586), .s(n18252), .op(n17588) );
  nand2_1 U18529 ( .ip1(n18843), .ip2(n17588), .op(n17589) );
  nand3_1 U18530 ( .ip1(n17591), .ip2(n17590), .ip3(n17589), .op(n17592) );
  nand2_1 U18531 ( .ip1(n17592), .ip2(n18888), .op(n17616) );
  mux2_1 U18532 ( .ip1(\ANSWER/mem[0][9][3] ), .ip2(\ANSWER/mem[1][9][3] ), 
        .s(n17610), .op(n17594) );
  mux2_1 U18533 ( .ip1(\ANSWER/mem[2][9][3] ), .ip2(\ANSWER/mem[3][9][3] ), 
        .s(n17602), .op(n17593) );
  mux2_1 U18534 ( .ip1(n17594), .ip2(n17593), .s(n17605), .op(n17598) );
  mux2_1 U18535 ( .ip1(\ANSWER/mem[4][9][3] ), .ip2(\ANSWER/mem[5][9][3] ), 
        .s(n17610), .op(n17596) );
  mux2_1 U18536 ( .ip1(\ANSWER/mem[6][9][3] ), .ip2(\ANSWER/mem[7][9][3] ), 
        .s(n17610), .op(n17595) );
  mux2_1 U18537 ( .ip1(n17596), .ip2(n17595), .s(n17605), .op(n17597) );
  mux2_1 U18538 ( .ip1(n17598), .ip2(n17597), .s(n18906), .op(n17600) );
  mux2_1 U18539 ( .ip1(\ANSWER/mem[8][9][3] ), .ip2(\ANSWER/mem[9][9][3] ), 
        .s(n17610), .op(n17599) );
  mux2_1 U18540 ( .ip1(n17600), .ip2(n17599), .s(n18092), .op(n17601) );
  nand2_1 U18541 ( .ip1(n18899), .ip2(n17601), .op(n17615) );
  mux2_1 U18542 ( .ip1(\ANSWER/mem[0][8][3] ), .ip2(\ANSWER/mem[1][8][3] ), 
        .s(n17602), .op(n17604) );
  mux2_1 U18543 ( .ip1(\ANSWER/mem[2][8][3] ), .ip2(\ANSWER/mem[3][8][3] ), 
        .s(n17602), .op(n17603) );
  mux2_1 U18544 ( .ip1(n17604), .ip2(n17603), .s(n17605), .op(n17609) );
  mux2_1 U18545 ( .ip1(\ANSWER/mem[4][8][3] ), .ip2(\ANSWER/mem[5][8][3] ), 
        .s(n17610), .op(n17607) );
  mux2_1 U18546 ( .ip1(\ANSWER/mem[6][8][3] ), .ip2(\ANSWER/mem[7][8][3] ), 
        .s(n17610), .op(n17606) );
  mux2_1 U18547 ( .ip1(n17607), .ip2(n17606), .s(n17605), .op(n17608) );
  mux2_1 U18548 ( .ip1(n17609), .ip2(n17608), .s(n18815), .op(n17612) );
  mux2_1 U18549 ( .ip1(\ANSWER/mem[8][8][3] ), .ip2(\ANSWER/mem[9][8][3] ), 
        .s(n17610), .op(n17611) );
  mux2_1 U18550 ( .ip1(n17612), .ip2(n17611), .s(n18092), .op(n17613) );
  nand2_1 U18551 ( .ip1(n18914), .ip2(n17613), .op(n17614) );
  nand3_1 U18552 ( .ip1(n17616), .ip2(n17615), .ip3(n17614), .op(\ANSWER/N484 ) );
  mux2_1 U18553 ( .ip1(\ANSWER/mem[0][1][4] ), .ip2(\ANSWER/mem[1][1][4] ), 
        .s(n17711), .op(n17618) );
  mux2_1 U18554 ( .ip1(\ANSWER/mem[2][1][4] ), .ip2(\ANSWER/mem[3][1][4] ), 
        .s(n18780), .op(n17617) );
  inv_1 U18555 ( .ip(n4366), .op(n17688) );
  mux2_1 U18556 ( .ip1(n17618), .ip2(n17617), .s(n17688), .op(n17622) );
  mux2_1 U18557 ( .ip1(\ANSWER/mem[4][1][4] ), .ip2(\ANSWER/mem[5][1][4] ), 
        .s(n18458), .op(n17620) );
  mux2_1 U18558 ( .ip1(\ANSWER/mem[6][1][4] ), .ip2(\ANSWER/mem[7][1][4] ), 
        .s(n18565), .op(n17619) );
  mux2_1 U18559 ( .ip1(n17620), .ip2(n17619), .s(n17688), .op(n17621) );
  mux2_1 U18560 ( .ip1(n17622), .ip2(n17621), .s(n18826), .op(n17624) );
  mux2_1 U18561 ( .ip1(\ANSWER/mem[8][1][4] ), .ip2(\ANSWER/mem[9][1][4] ), 
        .s(n18671), .op(n17623) );
  inv_1 U18562 ( .ip(n18165), .op(n18174) );
  mux2_1 U18563 ( .ip1(n17624), .ip2(n17623), .s(n18174), .op(n17625) );
  nand2_1 U18564 ( .ip1(n18872), .ip2(n17625), .op(n17698) );
  inv_1 U18565 ( .ip(n4362), .op(n17716) );
  mux2_1 U18566 ( .ip1(\ANSWER/mem[0][3][4] ), .ip2(\ANSWER/mem[1][3][4] ), 
        .s(n17716), .op(n17627) );
  mux2_1 U18567 ( .ip1(\ANSWER/mem[2][3][4] ), .ip2(\ANSWER/mem[3][3][4] ), 
        .s(n17716), .op(n17626) );
  mux2_1 U18568 ( .ip1(n17627), .ip2(n17626), .s(n17688), .op(n17631) );
  mux2_1 U18569 ( .ip1(\ANSWER/mem[4][3][4] ), .ip2(\ANSWER/mem[5][3][4] ), 
        .s(n17716), .op(n17629) );
  mux2_1 U18570 ( .ip1(\ANSWER/mem[6][3][4] ), .ip2(\ANSWER/mem[7][3][4] ), 
        .s(n17716), .op(n17628) );
  mux2_1 U18571 ( .ip1(n17629), .ip2(n17628), .s(n17688), .op(n17630) );
  mux2_1 U18572 ( .ip1(n17631), .ip2(n17630), .s(n18826), .op(n17633) );
  mux2_1 U18573 ( .ip1(\ANSWER/mem[8][3][4] ), .ip2(\ANSWER/mem[9][3][4] ), 
        .s(n17716), .op(n17632) );
  mux2_1 U18574 ( .ip1(n17633), .ip2(n17632), .s(n18174), .op(n17685) );
  mux2_1 U18575 ( .ip1(\ANSWER/mem[0][4][4] ), .ip2(\ANSWER/mem[1][4][4] ), 
        .s(n17716), .op(n17635) );
  mux2_1 U18576 ( .ip1(\ANSWER/mem[2][4][4] ), .ip2(\ANSWER/mem[3][4][4] ), 
        .s(n17716), .op(n17634) );
  mux2_1 U18577 ( .ip1(n17635), .ip2(n17634), .s(n17688), .op(n17639) );
  mux2_1 U18578 ( .ip1(\ANSWER/mem[4][4][4] ), .ip2(\ANSWER/mem[5][4][4] ), 
        .s(n17716), .op(n17637) );
  mux2_1 U18579 ( .ip1(\ANSWER/mem[6][4][4] ), .ip2(\ANSWER/mem[7][4][4] ), 
        .s(n17716), .op(n17636) );
  mux2_1 U18580 ( .ip1(n17637), .ip2(n17636), .s(n17688), .op(n17638) );
  mux2_1 U18581 ( .ip1(n17639), .ip2(n17638), .s(n18826), .op(n17641) );
  mux2_1 U18582 ( .ip1(\ANSWER/mem[8][4][4] ), .ip2(\ANSWER/mem[9][4][4] ), 
        .s(n17716), .op(n17640) );
  mux2_1 U18583 ( .ip1(n17641), .ip2(n17640), .s(n18174), .op(n17642) );
  and2_1 U18584 ( .ip1(n18843), .ip2(n17642), .op(n17684) );
  mux2_1 U18585 ( .ip1(\ANSWER/mem[0][2][4] ), .ip2(\ANSWER/mem[1][2][4] ), 
        .s(n17711), .op(n17644) );
  mux2_1 U18586 ( .ip1(\ANSWER/mem[2][2][4] ), .ip2(\ANSWER/mem[3][2][4] ), 
        .s(n18565), .op(n17643) );
  mux2_1 U18587 ( .ip1(n17644), .ip2(n17643), .s(n17688), .op(n17648) );
  mux2_1 U18588 ( .ip1(\ANSWER/mem[4][2][4] ), .ip2(\ANSWER/mem[5][2][4] ), 
        .s(n18780), .op(n17646) );
  mux2_1 U18589 ( .ip1(\ANSWER/mem[6][2][4] ), .ip2(\ANSWER/mem[7][2][4] ), 
        .s(n17716), .op(n17645) );
  mux2_1 U18590 ( .ip1(n17646), .ip2(n17645), .s(n17688), .op(n17647) );
  mux2_1 U18591 ( .ip1(n17648), .ip2(n17647), .s(n18826), .op(n17650) );
  mux2_1 U18592 ( .ip1(\ANSWER/mem[8][2][4] ), .ip2(\ANSWER/mem[9][2][4] ), 
        .s(n17716), .op(n17649) );
  mux2_1 U18593 ( .ip1(n17650), .ip2(n17649), .s(n18174), .op(n17651) );
  nand2_1 U18594 ( .ip1(n18884), .ip2(n17651), .op(n17682) );
  mux2_1 U18595 ( .ip1(\ANSWER/mem[0][0][4] ), .ip2(\ANSWER/mem[1][0][4] ), 
        .s(n18137), .op(n17653) );
  mux2_1 U18596 ( .ip1(\ANSWER/mem[2][0][4] ), .ip2(\ANSWER/mem[3][0][4] ), 
        .s(n18458), .op(n17652) );
  mux2_1 U18597 ( .ip1(n17653), .ip2(n17652), .s(n17688), .op(n17657) );
  mux2_1 U18598 ( .ip1(\ANSWER/mem[4][0][4] ), .ip2(\ANSWER/mem[5][0][4] ), 
        .s(n18029), .op(n17655) );
  mux2_1 U18599 ( .ip1(\ANSWER/mem[6][0][4] ), .ip2(\ANSWER/mem[7][0][4] ), 
        .s(n18671), .op(n17654) );
  mux2_1 U18600 ( .ip1(n17655), .ip2(n17654), .s(n17688), .op(n17656) );
  mux2_1 U18601 ( .ip1(n17657), .ip2(n17656), .s(n18826), .op(n17659) );
  mux2_1 U18602 ( .ip1(\ANSWER/mem[8][0][4] ), .ip2(\ANSWER/mem[9][0][4] ), 
        .s(n18137), .op(n17658) );
  mux2_1 U18603 ( .ip1(n17659), .ip2(n17658), .s(n18174), .op(n17660) );
  nand2_1 U18604 ( .ip1(n18800), .ip2(n17660), .op(n17681) );
  buf_1 U18605 ( .ip(n17716), .op(n17711) );
  mux2_1 U18606 ( .ip1(\ANSWER/mem[0][6][4] ), .ip2(\ANSWER/mem[1][6][4] ), 
        .s(n17711), .op(n17662) );
  mux2_1 U18607 ( .ip1(\ANSWER/mem[2][6][4] ), .ip2(\ANSWER/mem[3][6][4] ), 
        .s(n17711), .op(n17661) );
  mux2_1 U18608 ( .ip1(n17662), .ip2(n17661), .s(n17688), .op(n17666) );
  mux2_1 U18609 ( .ip1(\ANSWER/mem[4][6][4] ), .ip2(\ANSWER/mem[5][6][4] ), 
        .s(n17711), .op(n17664) );
  mux2_1 U18610 ( .ip1(\ANSWER/mem[6][6][4] ), .ip2(\ANSWER/mem[7][6][4] ), 
        .s(n17711), .op(n17663) );
  mux2_1 U18611 ( .ip1(n17664), .ip2(n17663), .s(n17581), .op(n17665) );
  mux2_1 U18612 ( .ip1(n17666), .ip2(n17665), .s(n18826), .op(n17668) );
  mux2_1 U18613 ( .ip1(\ANSWER/mem[8][6][4] ), .ip2(\ANSWER/mem[9][6][4] ), 
        .s(n17711), .op(n17667) );
  mux2_1 U18614 ( .ip1(n17668), .ip2(n17667), .s(n18174), .op(n17669) );
  nand2_1 U18615 ( .ip1(n18821), .ip2(n17669), .op(n17680) );
  mux2_1 U18616 ( .ip1(\ANSWER/mem[0][7][4] ), .ip2(\ANSWER/mem[1][7][4] ), 
        .s(n17711), .op(n17671) );
  mux2_1 U18617 ( .ip1(\ANSWER/mem[2][7][4] ), .ip2(\ANSWER/mem[3][7][4] ), 
        .s(n17711), .op(n17670) );
  mux2_1 U18618 ( .ip1(n17671), .ip2(n17670), .s(n18112), .op(n17675) );
  mux2_1 U18619 ( .ip1(\ANSWER/mem[4][7][4] ), .ip2(\ANSWER/mem[5][7][4] ), 
        .s(n17711), .op(n17673) );
  mux2_1 U18620 ( .ip1(\ANSWER/mem[6][7][4] ), .ip2(\ANSWER/mem[7][7][4] ), 
        .s(n17711), .op(n17672) );
  mux2_1 U18621 ( .ip1(n17673), .ip2(n17672), .s(n17688), .op(n17674) );
  mux2_1 U18622 ( .ip1(n17675), .ip2(n17674), .s(n18826), .op(n17677) );
  mux2_1 U18623 ( .ip1(\ANSWER/mem[8][7][4] ), .ip2(\ANSWER/mem[9][7][4] ), 
        .s(n17716), .op(n17676) );
  mux2_1 U18624 ( .ip1(n17677), .ip2(n17676), .s(n18174), .op(n17678) );
  nand2_1 U18625 ( .ip1(n18865), .ip2(n17678), .op(n17679) );
  nand4_1 U18626 ( .ip1(n17682), .ip2(n17681), .ip3(n17680), .ip4(n17679), 
        .op(n17683) );
  not_ab_or_c_or_d U18627 ( .ip1(n18854), .ip2(n17685), .ip3(n17684), .ip4(
        n17683), .op(n17697) );
  mux2_1 U18628 ( .ip1(\ANSWER/mem[0][5][4] ), .ip2(\ANSWER/mem[1][5][4] ), 
        .s(n17716), .op(n17687) );
  mux2_1 U18629 ( .ip1(\ANSWER/mem[2][5][4] ), .ip2(\ANSWER/mem[3][5][4] ), 
        .s(n17711), .op(n17686) );
  mux2_1 U18630 ( .ip1(n17687), .ip2(n17686), .s(n17688), .op(n17692) );
  mux2_1 U18631 ( .ip1(\ANSWER/mem[4][5][4] ), .ip2(\ANSWER/mem[5][5][4] ), 
        .s(n17711), .op(n17690) );
  mux2_1 U18632 ( .ip1(\ANSWER/mem[6][5][4] ), .ip2(\ANSWER/mem[7][5][4] ), 
        .s(n17711), .op(n17689) );
  mux2_1 U18633 ( .ip1(n17690), .ip2(n17689), .s(n17688), .op(n17691) );
  mux2_1 U18634 ( .ip1(n17692), .ip2(n17691), .s(n18826), .op(n17694) );
  mux2_1 U18635 ( .ip1(\ANSWER/mem[8][5][4] ), .ip2(\ANSWER/mem[9][5][4] ), 
        .s(n17711), .op(n17693) );
  mux2_1 U18636 ( .ip1(n17694), .ip2(n17693), .s(n18174), .op(n17695) );
  nand2_1 U18637 ( .ip1(n18832), .ip2(n17695), .op(n17696) );
  nand3_1 U18638 ( .ip1(n17698), .ip2(n17697), .ip3(n17696), .op(n17699) );
  nand2_1 U18639 ( .ip1(n17699), .ip2(n18888), .op(n17722) );
  mux2_1 U18640 ( .ip1(\ANSWER/mem[0][9][4] ), .ip2(\ANSWER/mem[1][9][4] ), 
        .s(n17716), .op(n17701) );
  mux2_1 U18641 ( .ip1(\ANSWER/mem[2][9][4] ), .ip2(\ANSWER/mem[3][9][4] ), 
        .s(n17711), .op(n17700) );
  mux2_1 U18642 ( .ip1(n17701), .ip2(n17700), .s(n18138), .op(n17705) );
  mux2_1 U18643 ( .ip1(\ANSWER/mem[4][9][4] ), .ip2(\ANSWER/mem[5][9][4] ), 
        .s(n17716), .op(n17703) );
  mux2_1 U18644 ( .ip1(\ANSWER/mem[6][9][4] ), .ip2(\ANSWER/mem[7][9][4] ), 
        .s(n17716), .op(n17702) );
  mux2_1 U18645 ( .ip1(n17703), .ip2(n17702), .s(n17990), .op(n17704) );
  mux2_1 U18646 ( .ip1(n17705), .ip2(n17704), .s(n18826), .op(n17707) );
  mux2_1 U18647 ( .ip1(\ANSWER/mem[8][9][4] ), .ip2(\ANSWER/mem[9][9][4] ), 
        .s(n17716), .op(n17706) );
  mux2_1 U18648 ( .ip1(n17707), .ip2(n17706), .s(n18174), .op(n17708) );
  nand2_1 U18649 ( .ip1(n18899), .ip2(n17708), .op(n17721) );
  mux2_1 U18650 ( .ip1(\ANSWER/mem[0][8][4] ), .ip2(\ANSWER/mem[1][8][4] ), 
        .s(n17716), .op(n17710) );
  mux2_1 U18651 ( .ip1(\ANSWER/mem[2][8][4] ), .ip2(\ANSWER/mem[3][8][4] ), 
        .s(n17711), .op(n17709) );
  mux2_1 U18652 ( .ip1(n17710), .ip2(n17709), .s(n18354), .op(n17715) );
  mux2_1 U18653 ( .ip1(\ANSWER/mem[4][8][4] ), .ip2(\ANSWER/mem[5][8][4] ), 
        .s(n17716), .op(n17713) );
  mux2_1 U18654 ( .ip1(\ANSWER/mem[6][8][4] ), .ip2(\ANSWER/mem[7][8][4] ), 
        .s(n17711), .op(n17712) );
  mux2_1 U18655 ( .ip1(n17713), .ip2(n17712), .s(n18112), .op(n17714) );
  mux2_1 U18656 ( .ip1(n17715), .ip2(n17714), .s(n18826), .op(n17718) );
  mux2_1 U18657 ( .ip1(\ANSWER/mem[8][8][4] ), .ip2(\ANSWER/mem[9][8][4] ), 
        .s(n17716), .op(n17717) );
  mux2_1 U18658 ( .ip1(n17718), .ip2(n17717), .s(n18174), .op(n17719) );
  nand2_1 U18659 ( .ip1(n18914), .ip2(n17719), .op(n17720) );
  nand3_1 U18660 ( .ip1(n17722), .ip2(n17721), .ip3(n17720), .op(\ANSWER/N483 ) );
  inv_1 U18661 ( .ip(n4362), .op(n17822) );
  mux2_1 U18662 ( .ip1(\ANSWER/mem[0][3][5] ), .ip2(\ANSWER/mem[1][3][5] ), 
        .s(n17822), .op(n17724) );
  mux2_1 U18663 ( .ip1(\ANSWER/mem[2][3][5] ), .ip2(\ANSWER/mem[3][3][5] ), 
        .s(n17822), .op(n17723) );
  inv_1 U18664 ( .ip(n4366), .op(n17794) );
  mux2_1 U18665 ( .ip1(n17724), .ip2(n17723), .s(n17794), .op(n17728) );
  mux2_1 U18666 ( .ip1(\ANSWER/mem[4][3][5] ), .ip2(\ANSWER/mem[5][3][5] ), 
        .s(n17822), .op(n17726) );
  mux2_1 U18667 ( .ip1(\ANSWER/mem[6][3][5] ), .ip2(\ANSWER/mem[7][3][5] ), 
        .s(n17822), .op(n17725) );
  mux2_1 U18668 ( .ip1(n17726), .ip2(n17725), .s(n17794), .op(n17727) );
  mux2_1 U18669 ( .ip1(n17728), .ip2(n17727), .s(n18848), .op(n17730) );
  mux2_1 U18670 ( .ip1(\ANSWER/mem[8][3][5] ), .ip2(\ANSWER/mem[9][3][5] ), 
        .s(n17822), .op(n17729) );
  mux2_1 U18671 ( .ip1(n17730), .ip2(n17729), .s(n18174), .op(n17731) );
  nand2_1 U18672 ( .ip1(n17731), .ip2(n18854), .op(n17804) );
  mux2_1 U18673 ( .ip1(\ANSWER/mem[0][1][5] ), .ip2(\ANSWER/mem[1][1][5] ), 
        .s(n17817), .op(n17733) );
  mux2_1 U18674 ( .ip1(\ANSWER/mem[2][1][5] ), .ip2(\ANSWER/mem[3][1][5] ), 
        .s(n17533), .op(n17732) );
  mux2_1 U18675 ( .ip1(n17733), .ip2(n17732), .s(n17794), .op(n17737) );
  mux2_1 U18676 ( .ip1(\ANSWER/mem[4][1][5] ), .ip2(\ANSWER/mem[5][1][5] ), 
        .s(n17387), .op(n17735) );
  mux2_1 U18677 ( .ip1(\ANSWER/mem[6][1][5] ), .ip2(\ANSWER/mem[7][1][5] ), 
        .s(n17344), .op(n17734) );
  mux2_1 U18678 ( .ip1(n17735), .ip2(n17734), .s(n17794), .op(n17736) );
  mux2_1 U18679 ( .ip1(n17737), .ip2(n17736), .s(n18848), .op(n17739) );
  mux2_1 U18680 ( .ip1(\ANSWER/mem[8][1][5] ), .ip2(\ANSWER/mem[9][1][5] ), 
        .s(n18616), .op(n17738) );
  mux2_1 U18681 ( .ip1(n17739), .ip2(n17738), .s(n18174), .op(n17791) );
  mux2_1 U18682 ( .ip1(\ANSWER/mem[0][5][5] ), .ip2(\ANSWER/mem[1][5][5] ), 
        .s(n17822), .op(n17741) );
  buf_1 U18683 ( .ip(n17822), .op(n17817) );
  mux2_1 U18684 ( .ip1(\ANSWER/mem[2][5][5] ), .ip2(\ANSWER/mem[3][5][5] ), 
        .s(n17817), .op(n17740) );
  mux2_1 U18685 ( .ip1(n17741), .ip2(n17740), .s(n17794), .op(n17745) );
  mux2_1 U18686 ( .ip1(\ANSWER/mem[4][5][5] ), .ip2(\ANSWER/mem[5][5][5] ), 
        .s(n17817), .op(n17743) );
  mux2_1 U18687 ( .ip1(\ANSWER/mem[6][5][5] ), .ip2(\ANSWER/mem[7][5][5] ), 
        .s(n17817), .op(n17742) );
  mux2_1 U18688 ( .ip1(n17743), .ip2(n17742), .s(n17794), .op(n17744) );
  mux2_1 U18689 ( .ip1(n17745), .ip2(n17744), .s(n18848), .op(n17747) );
  mux2_1 U18690 ( .ip1(\ANSWER/mem[8][5][5] ), .ip2(\ANSWER/mem[9][5][5] ), 
        .s(n17817), .op(n17746) );
  mux2_1 U18691 ( .ip1(n17747), .ip2(n17746), .s(n18174), .op(n17748) );
  and2_1 U18692 ( .ip1(n18832), .ip2(n17748), .op(n17790) );
  mux2_1 U18693 ( .ip1(\ANSWER/mem[0][2][5] ), .ip2(\ANSWER/mem[1][2][5] ), 
        .s(n18029), .op(n17750) );
  mux2_1 U18694 ( .ip1(\ANSWER/mem[2][2][5] ), .ip2(\ANSWER/mem[3][2][5] ), 
        .s(n17884), .op(n17749) );
  mux2_1 U18695 ( .ip1(n17750), .ip2(n17749), .s(n17794), .op(n17754) );
  mux2_1 U18696 ( .ip1(\ANSWER/mem[4][2][5] ), .ip2(\ANSWER/mem[5][2][5] ), 
        .s(n18616), .op(n17752) );
  mux2_1 U18697 ( .ip1(\ANSWER/mem[6][2][5] ), .ip2(\ANSWER/mem[7][2][5] ), 
        .s(n17822), .op(n17751) );
  mux2_1 U18698 ( .ip1(n17752), .ip2(n17751), .s(n17794), .op(n17753) );
  mux2_1 U18699 ( .ip1(n17754), .ip2(n17753), .s(n18848), .op(n17756) );
  mux2_1 U18700 ( .ip1(\ANSWER/mem[8][2][5] ), .ip2(\ANSWER/mem[9][2][5] ), 
        .s(n17822), .op(n17755) );
  mux2_1 U18701 ( .ip1(n17756), .ip2(n17755), .s(n18174), .op(n17757) );
  nand2_1 U18702 ( .ip1(n18884), .ip2(n17757), .op(n17788) );
  mux2_1 U18703 ( .ip1(\ANSWER/mem[0][6][5] ), .ip2(\ANSWER/mem[1][6][5] ), 
        .s(n17817), .op(n17759) );
  mux2_1 U18704 ( .ip1(\ANSWER/mem[2][6][5] ), .ip2(\ANSWER/mem[3][6][5] ), 
        .s(n17817), .op(n17758) );
  mux2_1 U18705 ( .ip1(n17759), .ip2(n17758), .s(n17794), .op(n17763) );
  mux2_1 U18706 ( .ip1(\ANSWER/mem[4][6][5] ), .ip2(\ANSWER/mem[5][6][5] ), 
        .s(n17817), .op(n17761) );
  mux2_1 U18707 ( .ip1(\ANSWER/mem[6][6][5] ), .ip2(\ANSWER/mem[7][6][5] ), 
        .s(n17817), .op(n17760) );
  mux2_1 U18708 ( .ip1(n17761), .ip2(n17760), .s(n18330), .op(n17762) );
  mux2_1 U18709 ( .ip1(n17763), .ip2(n17762), .s(n18848), .op(n17765) );
  mux2_1 U18710 ( .ip1(\ANSWER/mem[8][6][5] ), .ip2(\ANSWER/mem[9][6][5] ), 
        .s(n17817), .op(n17764) );
  mux2_1 U18711 ( .ip1(n17765), .ip2(n17764), .s(n18174), .op(n17766) );
  nand2_1 U18712 ( .ip1(n18821), .ip2(n17766), .op(n17787) );
  mux2_1 U18713 ( .ip1(\ANSWER/mem[0][0][5] ), .ip2(\ANSWER/mem[1][0][5] ), 
        .s(n17817), .op(n17768) );
  mux2_1 U18714 ( .ip1(\ANSWER/mem[2][0][5] ), .ip2(\ANSWER/mem[3][0][5] ), 
        .s(n18741), .op(n17767) );
  mux2_1 U18715 ( .ip1(n17768), .ip2(n17767), .s(n17794), .op(n17772) );
  mux2_1 U18716 ( .ip1(\ANSWER/mem[4][0][5] ), .ip2(\ANSWER/mem[5][0][5] ), 
        .s(n17387), .op(n17770) );
  mux2_1 U18717 ( .ip1(\ANSWER/mem[6][0][5] ), .ip2(\ANSWER/mem[7][0][5] ), 
        .s(n17533), .op(n17769) );
  mux2_1 U18718 ( .ip1(n17770), .ip2(n17769), .s(n17794), .op(n17771) );
  mux2_1 U18719 ( .ip1(n17772), .ip2(n17771), .s(n18848), .op(n17774) );
  mux2_1 U18720 ( .ip1(\ANSWER/mem[8][0][5] ), .ip2(\ANSWER/mem[9][0][5] ), 
        .s(n18741), .op(n17773) );
  mux2_1 U18721 ( .ip1(n17774), .ip2(n17773), .s(n18174), .op(n17775) );
  nand2_1 U18722 ( .ip1(n18800), .ip2(n17775), .op(n17786) );
  mux2_1 U18723 ( .ip1(\ANSWER/mem[0][7][5] ), .ip2(\ANSWER/mem[1][7][5] ), 
        .s(n17817), .op(n17777) );
  mux2_1 U18724 ( .ip1(\ANSWER/mem[2][7][5] ), .ip2(\ANSWER/mem[3][7][5] ), 
        .s(n17817), .op(n17776) );
  mux2_1 U18725 ( .ip1(n17777), .ip2(n17776), .s(n17990), .op(n17781) );
  mux2_1 U18726 ( .ip1(\ANSWER/mem[4][7][5] ), .ip2(\ANSWER/mem[5][7][5] ), 
        .s(n17817), .op(n17779) );
  mux2_1 U18727 ( .ip1(\ANSWER/mem[6][7][5] ), .ip2(\ANSWER/mem[7][7][5] ), 
        .s(n17817), .op(n17778) );
  mux2_1 U18728 ( .ip1(n17779), .ip2(n17778), .s(n18138), .op(n17780) );
  mux2_1 U18729 ( .ip1(n17781), .ip2(n17780), .s(n18848), .op(n17783) );
  mux2_1 U18730 ( .ip1(\ANSWER/mem[8][7][5] ), .ip2(\ANSWER/mem[9][7][5] ), 
        .s(n17822), .op(n17782) );
  mux2_1 U18731 ( .ip1(n17783), .ip2(n17782), .s(n18174), .op(n17784) );
  nand2_1 U18732 ( .ip1(n18865), .ip2(n17784), .op(n17785) );
  nand4_1 U18733 ( .ip1(n17788), .ip2(n17787), .ip3(n17786), .ip4(n17785), 
        .op(n17789) );
  not_ab_or_c_or_d U18734 ( .ip1(n17791), .ip2(n18872), .ip3(n17790), .ip4(
        n17789), .op(n17803) );
  mux2_1 U18735 ( .ip1(\ANSWER/mem[0][4][5] ), .ip2(\ANSWER/mem[1][4][5] ), 
        .s(n17822), .op(n17793) );
  mux2_1 U18736 ( .ip1(\ANSWER/mem[2][4][5] ), .ip2(\ANSWER/mem[3][4][5] ), 
        .s(n17822), .op(n17792) );
  mux2_1 U18737 ( .ip1(n17793), .ip2(n17792), .s(n17794), .op(n17798) );
  mux2_1 U18738 ( .ip1(\ANSWER/mem[4][4][5] ), .ip2(\ANSWER/mem[5][4][5] ), 
        .s(n17822), .op(n17796) );
  mux2_1 U18739 ( .ip1(\ANSWER/mem[6][4][5] ), .ip2(\ANSWER/mem[7][4][5] ), 
        .s(n17822), .op(n17795) );
  mux2_1 U18740 ( .ip1(n17796), .ip2(n17795), .s(n17794), .op(n17797) );
  mux2_1 U18741 ( .ip1(n17798), .ip2(n17797), .s(n18848), .op(n17800) );
  mux2_1 U18742 ( .ip1(\ANSWER/mem[8][4][5] ), .ip2(\ANSWER/mem[9][4][5] ), 
        .s(n17822), .op(n17799) );
  mux2_1 U18743 ( .ip1(n17800), .ip2(n17799), .s(n18174), .op(n17801) );
  nand2_1 U18744 ( .ip1(n18843), .ip2(n17801), .op(n17802) );
  nand3_1 U18745 ( .ip1(n17804), .ip2(n17803), .ip3(n17802), .op(n17805) );
  nand2_1 U18746 ( .ip1(n17805), .ip2(n18888), .op(n17828) );
  mux2_1 U18747 ( .ip1(\ANSWER/mem[0][8][5] ), .ip2(\ANSWER/mem[1][8][5] ), 
        .s(n17822), .op(n17807) );
  mux2_1 U18748 ( .ip1(\ANSWER/mem[2][8][5] ), .ip2(\ANSWER/mem[3][8][5] ), 
        .s(n17817), .op(n17806) );
  mux2_1 U18749 ( .ip1(n17807), .ip2(n17806), .s(n18435), .op(n17811) );
  mux2_1 U18750 ( .ip1(\ANSWER/mem[4][8][5] ), .ip2(\ANSWER/mem[5][8][5] ), 
        .s(n17822), .op(n17809) );
  mux2_1 U18751 ( .ip1(\ANSWER/mem[6][8][5] ), .ip2(\ANSWER/mem[7][8][5] ), 
        .s(n17822), .op(n17808) );
  mux2_1 U18752 ( .ip1(n17809), .ip2(n17808), .s(n17688), .op(n17810) );
  mux2_1 U18753 ( .ip1(n17811), .ip2(n17810), .s(n18848), .op(n17813) );
  mux2_1 U18754 ( .ip1(\ANSWER/mem[8][8][5] ), .ip2(\ANSWER/mem[9][8][5] ), 
        .s(n17822), .op(n17812) );
  mux2_1 U18755 ( .ip1(n17813), .ip2(n17812), .s(n18174), .op(n17814) );
  nand2_1 U18756 ( .ip1(n18914), .ip2(n17814), .op(n17827) );
  mux2_1 U18757 ( .ip1(\ANSWER/mem[0][9][5] ), .ip2(\ANSWER/mem[1][9][5] ), 
        .s(n17822), .op(n17816) );
  mux2_1 U18758 ( .ip1(\ANSWER/mem[2][9][5] ), .ip2(\ANSWER/mem[3][9][5] ), 
        .s(n17817), .op(n17815) );
  mux2_1 U18759 ( .ip1(n17816), .ip2(n17815), .s(n18330), .op(n17821) );
  mux2_1 U18760 ( .ip1(\ANSWER/mem[4][9][5] ), .ip2(\ANSWER/mem[5][9][5] ), 
        .s(n17822), .op(n17819) );
  mux2_1 U18761 ( .ip1(\ANSWER/mem[6][9][5] ), .ip2(\ANSWER/mem[7][9][5] ), 
        .s(n17817), .op(n17818) );
  mux2_1 U18762 ( .ip1(n17819), .ip2(n17818), .s(n17990), .op(n17820) );
  mux2_1 U18763 ( .ip1(n17821), .ip2(n17820), .s(n18848), .op(n17824) );
  mux2_1 U18764 ( .ip1(\ANSWER/mem[8][9][5] ), .ip2(\ANSWER/mem[9][9][5] ), 
        .s(n17822), .op(n17823) );
  mux2_1 U18765 ( .ip1(n17824), .ip2(n17823), .s(n18174), .op(n17825) );
  nand2_1 U18766 ( .ip1(n18899), .ip2(n17825), .op(n17826) );
  nand3_1 U18767 ( .ip1(n17828), .ip2(n17827), .ip3(n17826), .op(\ANSWER/N482 ) );
  inv_1 U18768 ( .ip(n4362), .op(n17884) );
  mux2_1 U18769 ( .ip1(\ANSWER/mem[0][0][6] ), .ip2(\ANSWER/mem[1][0][6] ), 
        .s(n17884), .op(n17830) );
  mux2_1 U18770 ( .ip1(\ANSWER/mem[2][0][6] ), .ip2(\ANSWER/mem[3][0][6] ), 
        .s(n17884), .op(n17829) );
  mux2_1 U18771 ( .ip1(n17830), .ip2(n17829), .s(n18354), .op(n17834) );
  mux2_1 U18772 ( .ip1(\ANSWER/mem[4][0][6] ), .ip2(\ANSWER/mem[5][0][6] ), 
        .s(n17884), .op(n17832) );
  mux2_1 U18773 ( .ip1(\ANSWER/mem[6][0][6] ), .ip2(\ANSWER/mem[7][0][6] ), 
        .s(n17884), .op(n17831) );
  mux2_1 U18774 ( .ip1(n17832), .ip2(n17831), .s(n18330), .op(n17833) );
  mux2_1 U18775 ( .ip1(n17834), .ip2(n17833), .s(n18837), .op(n17836) );
  mux2_1 U18776 ( .ip1(\ANSWER/mem[8][0][6] ), .ip2(\ANSWER/mem[9][0][6] ), 
        .s(n17884), .op(n17835) );
  inv_1 U18777 ( .ip(n18165), .op(n18073) );
  mux2_1 U18778 ( .ip1(n17836), .ip2(n17835), .s(n18073), .op(n17837) );
  nand2_1 U18779 ( .ip1(n17837), .ip2(n18800), .op(n17910) );
  inv_1 U18780 ( .ip(n4362), .op(n17928) );
  buf_1 U18781 ( .ip(n17928), .op(n17921) );
  mux2_1 U18782 ( .ip1(\ANSWER/mem[0][5][6] ), .ip2(\ANSWER/mem[1][5][6] ), 
        .s(n17921), .op(n17839) );
  mux2_1 U18783 ( .ip1(\ANSWER/mem[2][5][6] ), .ip2(\ANSWER/mem[3][5][6] ), 
        .s(n17928), .op(n17838) );
  mux2_1 U18784 ( .ip1(n17839), .ip2(n17838), .s(n17794), .op(n17843) );
  mux2_1 U18785 ( .ip1(\ANSWER/mem[4][5][6] ), .ip2(\ANSWER/mem[5][5][6] ), 
        .s(n17928), .op(n17841) );
  mux2_1 U18786 ( .ip1(\ANSWER/mem[6][5][6] ), .ip2(\ANSWER/mem[7][5][6] ), 
        .s(n17928), .op(n17840) );
  mux2_1 U18787 ( .ip1(n17841), .ip2(n17840), .s(n17605), .op(n17842) );
  mux2_1 U18788 ( .ip1(n17843), .ip2(n17842), .s(n18859), .op(n17845) );
  mux2_1 U18789 ( .ip1(\ANSWER/mem[8][5][6] ), .ip2(\ANSWER/mem[9][5][6] ), 
        .s(n17928), .op(n17844) );
  mux2_1 U18790 ( .ip1(n17845), .ip2(n17844), .s(n18073), .op(n17898) );
  mux2_1 U18791 ( .ip1(\ANSWER/mem[0][7][6] ), .ip2(\ANSWER/mem[1][7][6] ), 
        .s(n17928), .op(n17847) );
  mux2_1 U18792 ( .ip1(\ANSWER/mem[2][7][6] ), .ip2(\ANSWER/mem[3][7][6] ), 
        .s(n17928), .op(n17846) );
  mux2_1 U18793 ( .ip1(n17847), .ip2(n17846), .s(n17581), .op(n17851) );
  mux2_1 U18794 ( .ip1(\ANSWER/mem[4][7][6] ), .ip2(\ANSWER/mem[5][7][6] ), 
        .s(n17928), .op(n17849) );
  mux2_1 U18795 ( .ip1(\ANSWER/mem[6][7][6] ), .ip2(\ANSWER/mem[7][7][6] ), 
        .s(n17928), .op(n17848) );
  mux2_1 U18796 ( .ip1(n17849), .ip2(n17848), .s(n18435), .op(n17850) );
  mux2_1 U18797 ( .ip1(n17851), .ip2(n17850), .s(n18837), .op(n17853) );
  mux2_1 U18798 ( .ip1(\ANSWER/mem[8][7][6] ), .ip2(\ANSWER/mem[9][7][6] ), 
        .s(n17928), .op(n17852) );
  mux2_1 U18799 ( .ip1(n17853), .ip2(n17852), .s(n18073), .op(n17854) );
  and2_1 U18800 ( .ip1(n18865), .ip2(n17854), .op(n17897) );
  mux2_1 U18801 ( .ip1(\ANSWER/mem[0][6][6] ), .ip2(\ANSWER/mem[1][6][6] ), 
        .s(n17928), .op(n17856) );
  mux2_1 U18802 ( .ip1(\ANSWER/mem[2][6][6] ), .ip2(\ANSWER/mem[3][6][6] ), 
        .s(n17928), .op(n17855) );
  mux2_1 U18803 ( .ip1(n17856), .ip2(n17855), .s(n17366), .op(n17860) );
  mux2_1 U18804 ( .ip1(\ANSWER/mem[4][6][6] ), .ip2(\ANSWER/mem[5][6][6] ), 
        .s(n17928), .op(n17858) );
  mux2_1 U18805 ( .ip1(\ANSWER/mem[6][6][6] ), .ip2(\ANSWER/mem[7][6][6] ), 
        .s(n17928), .op(n17857) );
  mux2_1 U18806 ( .ip1(n17858), .ip2(n17857), .s(n18138), .op(n17859) );
  mux2_1 U18807 ( .ip1(n17860), .ip2(n17859), .s(n18848), .op(n17862) );
  mux2_1 U18808 ( .ip1(\ANSWER/mem[8][6][6] ), .ip2(\ANSWER/mem[9][6][6] ), 
        .s(n17928), .op(n17861) );
  mux2_1 U18809 ( .ip1(n17862), .ip2(n17861), .s(n18073), .op(n17863) );
  nand2_1 U18810 ( .ip1(n18821), .ip2(n17863), .op(n17895) );
  mux2_1 U18811 ( .ip1(\ANSWER/mem[0][4][6] ), .ip2(\ANSWER/mem[1][4][6] ), 
        .s(n17921), .op(n17865) );
  mux2_1 U18812 ( .ip1(\ANSWER/mem[2][4][6] ), .ip2(\ANSWER/mem[3][4][6] ), 
        .s(n17921), .op(n17864) );
  mux2_1 U18813 ( .ip1(n17865), .ip2(n17864), .s(n18435), .op(n17869) );
  mux2_1 U18814 ( .ip1(\ANSWER/mem[4][4][6] ), .ip2(\ANSWER/mem[5][4][6] ), 
        .s(n17921), .op(n17867) );
  mux2_1 U18815 ( .ip1(\ANSWER/mem[6][4][6] ), .ip2(\ANSWER/mem[7][4][6] ), 
        .s(n17921), .op(n17866) );
  mux2_1 U18816 ( .ip1(n17867), .ip2(n17866), .s(n17688), .op(n17868) );
  mux2_1 U18817 ( .ip1(n17869), .ip2(n17868), .s(n18859), .op(n17871) );
  mux2_1 U18818 ( .ip1(\ANSWER/mem[8][4][6] ), .ip2(\ANSWER/mem[9][4][6] ), 
        .s(n17921), .op(n17870) );
  mux2_1 U18819 ( .ip1(n17871), .ip2(n17870), .s(n18073), .op(n17872) );
  nand2_1 U18820 ( .ip1(n18843), .ip2(n17872), .op(n17894) );
  mux2_1 U18821 ( .ip1(\ANSWER/mem[0][1][6] ), .ip2(\ANSWER/mem[1][1][6] ), 
        .s(n17884), .op(n17874) );
  mux2_1 U18822 ( .ip1(\ANSWER/mem[2][1][6] ), .ip2(\ANSWER/mem[3][1][6] ), 
        .s(n17884), .op(n17873) );
  mux2_1 U18823 ( .ip1(n17874), .ip2(n17873), .s(n18435), .op(n17878) );
  mux2_1 U18824 ( .ip1(\ANSWER/mem[4][1][6] ), .ip2(\ANSWER/mem[5][1][6] ), 
        .s(n17884), .op(n17876) );
  mux2_1 U18825 ( .ip1(\ANSWER/mem[6][1][6] ), .ip2(\ANSWER/mem[7][1][6] ), 
        .s(n17884), .op(n17875) );
  mux2_1 U18826 ( .ip1(n17876), .ip2(n17875), .s(n4456), .op(n17877) );
  mux2_1 U18827 ( .ip1(n17878), .ip2(n17877), .s(n18859), .op(n17880) );
  mux2_1 U18828 ( .ip1(\ANSWER/mem[8][1][6] ), .ip2(\ANSWER/mem[9][1][6] ), 
        .s(n17884), .op(n17879) );
  mux2_1 U18829 ( .ip1(n17880), .ip2(n17879), .s(n18073), .op(n17881) );
  nand2_1 U18830 ( .ip1(n18872), .ip2(n17881), .op(n17893) );
  mux2_1 U18831 ( .ip1(\ANSWER/mem[0][2][6] ), .ip2(\ANSWER/mem[1][2][6] ), 
        .s(n17884), .op(n17883) );
  mux2_1 U18832 ( .ip1(\ANSWER/mem[2][2][6] ), .ip2(\ANSWER/mem[3][2][6] ), 
        .s(n17884), .op(n17882) );
  mux2_1 U18833 ( .ip1(n17883), .ip2(n17882), .s(n18354), .op(n17888) );
  mux2_1 U18834 ( .ip1(\ANSWER/mem[4][2][6] ), .ip2(\ANSWER/mem[5][2][6] ), 
        .s(n17884), .op(n17886) );
  mux2_1 U18835 ( .ip1(\ANSWER/mem[6][2][6] ), .ip2(\ANSWER/mem[7][2][6] ), 
        .s(n17921), .op(n17885) );
  mux2_1 U18836 ( .ip1(n17886), .ip2(n17885), .s(n17581), .op(n17887) );
  mux2_1 U18837 ( .ip1(n17888), .ip2(n17887), .s(n18837), .op(n17890) );
  mux2_1 U18838 ( .ip1(\ANSWER/mem[8][2][6] ), .ip2(\ANSWER/mem[9][2][6] ), 
        .s(n17921), .op(n17889) );
  mux2_1 U18839 ( .ip1(n17890), .ip2(n17889), .s(n18073), .op(n17891) );
  nand2_1 U18840 ( .ip1(n18884), .ip2(n17891), .op(n17892) );
  nand4_1 U18841 ( .ip1(n17895), .ip2(n17894), .ip3(n17893), .ip4(n17892), 
        .op(n17896) );
  not_ab_or_c_or_d U18842 ( .ip1(n18832), .ip2(n17898), .ip3(n17897), .ip4(
        n17896), .op(n17909) );
  mux2_1 U18843 ( .ip1(\ANSWER/mem[0][3][6] ), .ip2(\ANSWER/mem[1][3][6] ), 
        .s(n17921), .op(n17900) );
  mux2_1 U18844 ( .ip1(\ANSWER/mem[2][3][6] ), .ip2(\ANSWER/mem[3][3][6] ), 
        .s(n17921), .op(n17899) );
  mux2_1 U18845 ( .ip1(n17900), .ip2(n17899), .s(n15636), .op(n17904) );
  mux2_1 U18846 ( .ip1(\ANSWER/mem[4][3][6] ), .ip2(\ANSWER/mem[5][3][6] ), 
        .s(n17921), .op(n17902) );
  mux2_1 U18847 ( .ip1(\ANSWER/mem[6][3][6] ), .ip2(\ANSWER/mem[7][3][6] ), 
        .s(n17921), .op(n17901) );
  mux2_1 U18848 ( .ip1(n17902), .ip2(n17901), .s(n18138), .op(n17903) );
  mux2_1 U18849 ( .ip1(n17904), .ip2(n17903), .s(n18848), .op(n17906) );
  mux2_1 U18850 ( .ip1(\ANSWER/mem[8][3][6] ), .ip2(\ANSWER/mem[9][3][6] ), 
        .s(n17921), .op(n17905) );
  mux2_1 U18851 ( .ip1(n17906), .ip2(n17905), .s(n18073), .op(n17907) );
  nand2_1 U18852 ( .ip1(n18854), .ip2(n17907), .op(n17908) );
  nand3_1 U18853 ( .ip1(n17910), .ip2(n17909), .ip3(n17908), .op(n17911) );
  nand2_1 U18854 ( .ip1(n17911), .ip2(n18888), .op(n17934) );
  mux2_1 U18855 ( .ip1(\ANSWER/mem[0][8][6] ), .ip2(\ANSWER/mem[1][8][6] ), 
        .s(n17928), .op(n17913) );
  mux2_1 U18856 ( .ip1(\ANSWER/mem[2][8][6] ), .ip2(\ANSWER/mem[3][8][6] ), 
        .s(n17921), .op(n17912) );
  mux2_1 U18857 ( .ip1(n17913), .ip2(n17912), .s(n18354), .op(n17917) );
  mux2_1 U18858 ( .ip1(\ANSWER/mem[4][8][6] ), .ip2(\ANSWER/mem[5][8][6] ), 
        .s(n17928), .op(n17915) );
  mux2_1 U18859 ( .ip1(\ANSWER/mem[6][8][6] ), .ip2(\ANSWER/mem[7][8][6] ), 
        .s(n17928), .op(n17914) );
  mux2_1 U18860 ( .ip1(n17915), .ip2(n17914), .s(n18138), .op(n17916) );
  mux2_1 U18861 ( .ip1(n17917), .ip2(n17916), .s(n18848), .op(n17919) );
  mux2_1 U18862 ( .ip1(\ANSWER/mem[8][8][6] ), .ip2(\ANSWER/mem[9][8][6] ), 
        .s(n17928), .op(n17918) );
  mux2_1 U18863 ( .ip1(n17919), .ip2(n17918), .s(n18073), .op(n17920) );
  nand2_1 U18864 ( .ip1(n18914), .ip2(n17920), .op(n17933) );
  mux2_1 U18865 ( .ip1(\ANSWER/mem[0][9][6] ), .ip2(\ANSWER/mem[1][9][6] ), 
        .s(n17921), .op(n17923) );
  mux2_1 U18866 ( .ip1(\ANSWER/mem[2][9][6] ), .ip2(\ANSWER/mem[3][9][6] ), 
        .s(n17921), .op(n17922) );
  mux2_1 U18867 ( .ip1(n17923), .ip2(n17922), .s(n17605), .op(n17927) );
  mux2_1 U18868 ( .ip1(\ANSWER/mem[4][9][6] ), .ip2(\ANSWER/mem[5][9][6] ), 
        .s(n17928), .op(n17925) );
  mux2_1 U18869 ( .ip1(\ANSWER/mem[6][9][6] ), .ip2(\ANSWER/mem[7][9][6] ), 
        .s(n17928), .op(n17924) );
  mux2_1 U18870 ( .ip1(n17925), .ip2(n17924), .s(n18330), .op(n17926) );
  mux2_1 U18871 ( .ip1(n17927), .ip2(n17926), .s(n18859), .op(n17930) );
  mux2_1 U18872 ( .ip1(\ANSWER/mem[8][9][6] ), .ip2(\ANSWER/mem[9][9][6] ), 
        .s(n17928), .op(n17929) );
  mux2_1 U18873 ( .ip1(n17930), .ip2(n17929), .s(n18073), .op(n17931) );
  nand2_1 U18874 ( .ip1(n18899), .ip2(n17931), .op(n17932) );
  nand3_1 U18875 ( .ip1(n17934), .ip2(n17933), .ip3(n17932), .op(\ANSWER/N481 ) );
  mux2_1 U18876 ( .ip1(\ANSWER/mem[0][0][7] ), .ip2(\ANSWER/mem[1][0][7] ), 
        .s(n18351), .op(n17936) );
  mux2_1 U18877 ( .ip1(\ANSWER/mem[2][0][7] ), .ip2(\ANSWER/mem[3][0][7] ), 
        .s(n18458), .op(n17935) );
  inv_1 U18878 ( .ip(n4366), .op(n17990) );
  mux2_1 U18879 ( .ip1(n17936), .ip2(n17935), .s(n17990), .op(n17940) );
  mux2_1 U18880 ( .ip1(\ANSWER/mem[4][0][7] ), .ip2(\ANSWER/mem[5][0][7] ), 
        .s(n18029), .op(n17938) );
  mux2_1 U18881 ( .ip1(\ANSWER/mem[6][0][7] ), .ip2(\ANSWER/mem[7][0][7] ), 
        .s(n17921), .op(n17937) );
  mux2_1 U18882 ( .ip1(n17938), .ip2(n17937), .s(n17990), .op(n17939) );
  mux2_1 U18883 ( .ip1(n17940), .ip2(n17939), .s(n18806), .op(n17942) );
  mux2_1 U18884 ( .ip1(\ANSWER/mem[8][0][7] ), .ip2(\ANSWER/mem[9][0][7] ), 
        .s(n15643), .op(n17941) );
  mux2_1 U18885 ( .ip1(n17942), .ip2(n17941), .s(n18073), .op(n17943) );
  nand2_1 U18886 ( .ip1(n17943), .ip2(n18800), .op(n18016) );
  inv_1 U18887 ( .ip(n4362), .op(n18034) );
  buf_1 U18888 ( .ip(n18034), .op(n18029) );
  mux2_1 U18889 ( .ip1(\ANSWER/mem[0][3][7] ), .ip2(\ANSWER/mem[1][3][7] ), 
        .s(n18029), .op(n17945) );
  mux2_1 U18890 ( .ip1(\ANSWER/mem[2][3][7] ), .ip2(\ANSWER/mem[3][3][7] ), 
        .s(n18029), .op(n17944) );
  mux2_1 U18891 ( .ip1(n17945), .ip2(n17944), .s(n17990), .op(n17949) );
  mux2_1 U18892 ( .ip1(\ANSWER/mem[4][3][7] ), .ip2(\ANSWER/mem[5][3][7] ), 
        .s(n18029), .op(n17947) );
  mux2_1 U18893 ( .ip1(\ANSWER/mem[6][3][7] ), .ip2(\ANSWER/mem[7][3][7] ), 
        .s(n18029), .op(n17946) );
  mux2_1 U18894 ( .ip1(n17947), .ip2(n17946), .s(n17990), .op(n17948) );
  mux2_1 U18895 ( .ip1(n17949), .ip2(n17948), .s(n18806), .op(n17951) );
  mux2_1 U18896 ( .ip1(\ANSWER/mem[8][3][7] ), .ip2(\ANSWER/mem[9][3][7] ), 
        .s(n18029), .op(n17950) );
  mux2_1 U18897 ( .ip1(n17951), .ip2(n17950), .s(n18073), .op(n18004) );
  mux2_1 U18898 ( .ip1(\ANSWER/mem[0][4][7] ), .ip2(\ANSWER/mem[1][4][7] ), 
        .s(n18029), .op(n17953) );
  mux2_1 U18899 ( .ip1(\ANSWER/mem[2][4][7] ), .ip2(\ANSWER/mem[3][4][7] ), 
        .s(n18029), .op(n17952) );
  mux2_1 U18900 ( .ip1(n17953), .ip2(n17952), .s(n17990), .op(n17957) );
  mux2_1 U18901 ( .ip1(\ANSWER/mem[4][4][7] ), .ip2(\ANSWER/mem[5][4][7] ), 
        .s(n18029), .op(n17955) );
  mux2_1 U18902 ( .ip1(\ANSWER/mem[6][4][7] ), .ip2(\ANSWER/mem[7][4][7] ), 
        .s(n18029), .op(n17954) );
  mux2_1 U18903 ( .ip1(n17955), .ip2(n17954), .s(n17990), .op(n17956) );
  mux2_1 U18904 ( .ip1(n17957), .ip2(n17956), .s(n18806), .op(n17959) );
  mux2_1 U18905 ( .ip1(\ANSWER/mem[8][4][7] ), .ip2(\ANSWER/mem[9][4][7] ), 
        .s(n18029), .op(n17958) );
  mux2_1 U18906 ( .ip1(n17959), .ip2(n17958), .s(n18073), .op(n17960) );
  and2_1 U18907 ( .ip1(n18843), .ip2(n17960), .op(n18003) );
  mux2_1 U18908 ( .ip1(\ANSWER/mem[0][6][7] ), .ip2(\ANSWER/mem[1][6][7] ), 
        .s(n18034), .op(n17962) );
  mux2_1 U18909 ( .ip1(\ANSWER/mem[2][6][7] ), .ip2(\ANSWER/mem[3][6][7] ), 
        .s(n18034), .op(n17961) );
  mux2_1 U18910 ( .ip1(n17962), .ip2(n17961), .s(n17990), .op(n17966) );
  mux2_1 U18911 ( .ip1(\ANSWER/mem[4][6][7] ), .ip2(\ANSWER/mem[5][6][7] ), 
        .s(n18034), .op(n17964) );
  mux2_1 U18912 ( .ip1(\ANSWER/mem[6][6][7] ), .ip2(\ANSWER/mem[7][6][7] ), 
        .s(n18034), .op(n17963) );
  mux2_1 U18913 ( .ip1(n17964), .ip2(n17963), .s(n18138), .op(n17965) );
  mux2_1 U18914 ( .ip1(n17966), .ip2(n17965), .s(n18806), .op(n17968) );
  mux2_1 U18915 ( .ip1(\ANSWER/mem[8][6][7] ), .ip2(\ANSWER/mem[9][6][7] ), 
        .s(n18034), .op(n17967) );
  mux2_1 U18916 ( .ip1(n17968), .ip2(n17967), .s(n18073), .op(n17969) );
  nand2_1 U18917 ( .ip1(n18821), .ip2(n17969), .op(n18001) );
  mux2_1 U18918 ( .ip1(\ANSWER/mem[0][5][7] ), .ip2(\ANSWER/mem[1][5][7] ), 
        .s(n18029), .op(n17971) );
  mux2_1 U18919 ( .ip1(\ANSWER/mem[2][5][7] ), .ip2(\ANSWER/mem[3][5][7] ), 
        .s(n18034), .op(n17970) );
  mux2_1 U18920 ( .ip1(n17971), .ip2(n17970), .s(n17990), .op(n17975) );
  mux2_1 U18921 ( .ip1(\ANSWER/mem[4][5][7] ), .ip2(\ANSWER/mem[5][5][7] ), 
        .s(n18034), .op(n17973) );
  mux2_1 U18922 ( .ip1(\ANSWER/mem[6][5][7] ), .ip2(\ANSWER/mem[7][5][7] ), 
        .s(n18034), .op(n17972) );
  mux2_1 U18923 ( .ip1(n17973), .ip2(n17972), .s(n17990), .op(n17974) );
  mux2_1 U18924 ( .ip1(n17975), .ip2(n17974), .s(n18806), .op(n17977) );
  mux2_1 U18925 ( .ip1(\ANSWER/mem[8][5][7] ), .ip2(\ANSWER/mem[9][5][7] ), 
        .s(n18034), .op(n17976) );
  mux2_1 U18926 ( .ip1(n17977), .ip2(n17976), .s(n18073), .op(n17978) );
  nand2_1 U18927 ( .ip1(n18832), .ip2(n17978), .op(n18000) );
  mux2_1 U18928 ( .ip1(\ANSWER/mem[0][2][7] ), .ip2(\ANSWER/mem[1][2][7] ), 
        .s(n18351), .op(n17980) );
  mux2_1 U18929 ( .ip1(\ANSWER/mem[2][2][7] ), .ip2(\ANSWER/mem[3][2][7] ), 
        .s(n18780), .op(n17979) );
  mux2_1 U18930 ( .ip1(n17980), .ip2(n17979), .s(n17990), .op(n17984) );
  mux2_1 U18931 ( .ip1(\ANSWER/mem[4][2][7] ), .ip2(\ANSWER/mem[5][2][7] ), 
        .s(n18458), .op(n17982) );
  mux2_1 U18932 ( .ip1(\ANSWER/mem[6][2][7] ), .ip2(\ANSWER/mem[7][2][7] ), 
        .s(n18029), .op(n17981) );
  mux2_1 U18933 ( .ip1(n17982), .ip2(n17981), .s(n17990), .op(n17983) );
  mux2_1 U18934 ( .ip1(n17984), .ip2(n17983), .s(n18806), .op(n17986) );
  mux2_1 U18935 ( .ip1(\ANSWER/mem[8][2][7] ), .ip2(\ANSWER/mem[9][2][7] ), 
        .s(n18029), .op(n17985) );
  mux2_1 U18936 ( .ip1(n17986), .ip2(n17985), .s(n18073), .op(n17987) );
  nand2_1 U18937 ( .ip1(n18884), .ip2(n17987), .op(n17999) );
  mux2_1 U18938 ( .ip1(\ANSWER/mem[0][1][7] ), .ip2(\ANSWER/mem[1][1][7] ), 
        .s(n17711), .op(n17989) );
  mux2_1 U18939 ( .ip1(\ANSWER/mem[2][1][7] ), .ip2(\ANSWER/mem[3][1][7] ), 
        .s(n17921), .op(n17988) );
  mux2_1 U18940 ( .ip1(n17989), .ip2(n17988), .s(n17990), .op(n17994) );
  mux2_1 U18941 ( .ip1(\ANSWER/mem[4][1][7] ), .ip2(\ANSWER/mem[5][1][7] ), 
        .s(n18565), .op(n17992) );
  mux2_1 U18942 ( .ip1(\ANSWER/mem[6][1][7] ), .ip2(\ANSWER/mem[7][1][7] ), 
        .s(n18671), .op(n17991) );
  mux2_1 U18943 ( .ip1(n17992), .ip2(n17991), .s(n17990), .op(n17993) );
  mux2_1 U18944 ( .ip1(n17994), .ip2(n17993), .s(n18806), .op(n17996) );
  mux2_1 U18945 ( .ip1(\ANSWER/mem[8][1][7] ), .ip2(\ANSWER/mem[9][1][7] ), 
        .s(n18137), .op(n17995) );
  mux2_1 U18946 ( .ip1(n17996), .ip2(n17995), .s(n18073), .op(n17997) );
  nand2_1 U18947 ( .ip1(n18872), .ip2(n17997), .op(n17998) );
  nand4_1 U18948 ( .ip1(n18001), .ip2(n18000), .ip3(n17999), .ip4(n17998), 
        .op(n18002) );
  not_ab_or_c_or_d U18949 ( .ip1(n18854), .ip2(n18004), .ip3(n18003), .ip4(
        n18002), .op(n18015) );
  mux2_1 U18950 ( .ip1(\ANSWER/mem[0][7][7] ), .ip2(\ANSWER/mem[1][7][7] ), 
        .s(n18034), .op(n18006) );
  mux2_1 U18951 ( .ip1(\ANSWER/mem[2][7][7] ), .ip2(\ANSWER/mem[3][7][7] ), 
        .s(n18034), .op(n18005) );
  mux2_1 U18952 ( .ip1(n18006), .ip2(n18005), .s(n17794), .op(n18010) );
  mux2_1 U18953 ( .ip1(\ANSWER/mem[4][7][7] ), .ip2(\ANSWER/mem[5][7][7] ), 
        .s(n18034), .op(n18008) );
  mux2_1 U18954 ( .ip1(\ANSWER/mem[6][7][7] ), .ip2(\ANSWER/mem[7][7][7] ), 
        .s(n18034), .op(n18007) );
  mux2_1 U18955 ( .ip1(n18008), .ip2(n18007), .s(n17688), .op(n18009) );
  mux2_1 U18956 ( .ip1(n18010), .ip2(n18009), .s(n18806), .op(n18012) );
  mux2_1 U18957 ( .ip1(\ANSWER/mem[8][7][7] ), .ip2(\ANSWER/mem[9][7][7] ), 
        .s(n18034), .op(n18011) );
  mux2_1 U18958 ( .ip1(n18012), .ip2(n18011), .s(n18073), .op(n18013) );
  nand2_1 U18959 ( .ip1(n18865), .ip2(n18013), .op(n18014) );
  nand3_1 U18960 ( .ip1(n18016), .ip2(n18015), .ip3(n18014), .op(n18017) );
  nand2_1 U18961 ( .ip1(n18017), .ip2(n18888), .op(n18040) );
  mux2_1 U18962 ( .ip1(\ANSWER/mem[0][9][7] ), .ip2(\ANSWER/mem[1][9][7] ), 
        .s(n18029), .op(n18019) );
  mux2_1 U18963 ( .ip1(\ANSWER/mem[2][9][7] ), .ip2(\ANSWER/mem[3][9][7] ), 
        .s(n18034), .op(n18018) );
  mux2_1 U18964 ( .ip1(n18019), .ip2(n18018), .s(n18112), .op(n18023) );
  mux2_1 U18965 ( .ip1(\ANSWER/mem[4][9][7] ), .ip2(\ANSWER/mem[5][9][7] ), 
        .s(n18029), .op(n18021) );
  mux2_1 U18966 ( .ip1(\ANSWER/mem[6][9][7] ), .ip2(\ANSWER/mem[7][9][7] ), 
        .s(n18034), .op(n18020) );
  mux2_1 U18967 ( .ip1(n18021), .ip2(n18020), .s(n18354), .op(n18022) );
  mux2_1 U18968 ( .ip1(n18023), .ip2(n18022), .s(n18806), .op(n18025) );
  mux2_1 U18969 ( .ip1(\ANSWER/mem[8][9][7] ), .ip2(\ANSWER/mem[9][9][7] ), 
        .s(n18034), .op(n18024) );
  mux2_1 U18970 ( .ip1(n18025), .ip2(n18024), .s(n18073), .op(n18026) );
  nand2_1 U18971 ( .ip1(n18899), .ip2(n18026), .op(n18039) );
  mux2_1 U18972 ( .ip1(\ANSWER/mem[0][8][7] ), .ip2(\ANSWER/mem[1][8][7] ), 
        .s(n18034), .op(n18028) );
  mux2_1 U18973 ( .ip1(\ANSWER/mem[2][8][7] ), .ip2(\ANSWER/mem[3][8][7] ), 
        .s(n18034), .op(n18027) );
  mux2_1 U18974 ( .ip1(n18028), .ip2(n18027), .s(n18138), .op(n18033) );
  mux2_1 U18975 ( .ip1(\ANSWER/mem[4][8][7] ), .ip2(\ANSWER/mem[5][8][7] ), 
        .s(n18029), .op(n18031) );
  mux2_1 U18976 ( .ip1(\ANSWER/mem[6][8][7] ), .ip2(\ANSWER/mem[7][8][7] ), 
        .s(n18034), .op(n18030) );
  mux2_1 U18977 ( .ip1(n18031), .ip2(n18030), .s(n17605), .op(n18032) );
  mux2_1 U18978 ( .ip1(n18033), .ip2(n18032), .s(n18806), .op(n18036) );
  mux2_1 U18979 ( .ip1(\ANSWER/mem[8][8][7] ), .ip2(\ANSWER/mem[9][8][7] ), 
        .s(n18034), .op(n18035) );
  mux2_1 U18980 ( .ip1(n18036), .ip2(n18035), .s(n18073), .op(n18037) );
  nand2_1 U18981 ( .ip1(n18914), .ip2(n18037), .op(n18038) );
  nand3_1 U18982 ( .ip1(n18040), .ip2(n18039), .ip3(n18038), .op(\ANSWER/N480 ) );
  inv_1 U18983 ( .ip(n4362), .op(n18143) );
  buf_1 U18984 ( .ip(n18143), .op(n18137) );
  mux2_1 U18985 ( .ip1(\ANSWER/mem[0][4][8] ), .ip2(\ANSWER/mem[1][4][8] ), 
        .s(n18137), .op(n18042) );
  mux2_1 U18986 ( .ip1(\ANSWER/mem[2][4][8] ), .ip2(\ANSWER/mem[3][4][8] ), 
        .s(n18137), .op(n18041) );
  inv_1 U18987 ( .ip(n4366), .op(n18112) );
  mux2_1 U18988 ( .ip1(n18042), .ip2(n18041), .s(n18112), .op(n18046) );
  mux2_1 U18989 ( .ip1(\ANSWER/mem[4][4][8] ), .ip2(\ANSWER/mem[5][4][8] ), 
        .s(n18137), .op(n18044) );
  mux2_1 U18990 ( .ip1(\ANSWER/mem[6][4][8] ), .ip2(\ANSWER/mem[7][4][8] ), 
        .s(n18137), .op(n18043) );
  mux2_1 U18991 ( .ip1(n18044), .ip2(n18043), .s(n18112), .op(n18045) );
  mux2_1 U18992 ( .ip1(n18046), .ip2(n18045), .s(n18837), .op(n18048) );
  mux2_1 U18993 ( .ip1(\ANSWER/mem[8][4][8] ), .ip2(\ANSWER/mem[9][4][8] ), 
        .s(n18137), .op(n18047) );
  mux2_1 U18994 ( .ip1(n18048), .ip2(n18047), .s(n18092), .op(n18049) );
  nand2_1 U18995 ( .ip1(n18049), .ip2(n18843), .op(n18124) );
  mux2_1 U18996 ( .ip1(\ANSWER/mem[0][1][8] ), .ip2(\ANSWER/mem[1][1][8] ), 
        .s(n18671), .op(n18051) );
  mux2_1 U18997 ( .ip1(\ANSWER/mem[2][1][8] ), .ip2(\ANSWER/mem[3][1][8] ), 
        .s(n17610), .op(n18050) );
  mux2_1 U18998 ( .ip1(n18051), .ip2(n18050), .s(n18112), .op(n18055) );
  mux2_1 U18999 ( .ip1(\ANSWER/mem[4][1][8] ), .ip2(\ANSWER/mem[5][1][8] ), 
        .s(n17564), .op(n18053) );
  mux2_1 U19000 ( .ip1(\ANSWER/mem[6][1][8] ), .ip2(\ANSWER/mem[7][1][8] ), 
        .s(n15643), .op(n18052) );
  mux2_1 U19001 ( .ip1(n18053), .ip2(n18052), .s(n18112), .op(n18054) );
  mux2_1 U19002 ( .ip1(n18055), .ip2(n18054), .s(n18815), .op(n18057) );
  mux2_1 U19003 ( .ip1(\ANSWER/mem[8][1][8] ), .ip2(\ANSWER/mem[9][1][8] ), 
        .s(n18137), .op(n18056) );
  mux2_1 U19004 ( .ip1(n18057), .ip2(n18056), .s(n18073), .op(n18111) );
  mux2_1 U19005 ( .ip1(\ANSWER/mem[0][2][8] ), .ip2(\ANSWER/mem[1][2][8] ), 
        .s(n18780), .op(n18059) );
  mux2_1 U19006 ( .ip1(\ANSWER/mem[2][2][8] ), .ip2(\ANSWER/mem[3][2][8] ), 
        .s(n15643), .op(n18058) );
  mux2_1 U19007 ( .ip1(n18059), .ip2(n18058), .s(n18112), .op(n18063) );
  mux2_1 U19008 ( .ip1(\ANSWER/mem[4][2][8] ), .ip2(\ANSWER/mem[5][2][8] ), 
        .s(n18565), .op(n18061) );
  mux2_1 U19009 ( .ip1(\ANSWER/mem[6][2][8] ), .ip2(\ANSWER/mem[7][2][8] ), 
        .s(n18137), .op(n18060) );
  mux2_1 U19010 ( .ip1(n18061), .ip2(n18060), .s(n18112), .op(n18062) );
  mux2_1 U19011 ( .ip1(n18063), .ip2(n18062), .s(n18848), .op(n18065) );
  mux2_1 U19012 ( .ip1(\ANSWER/mem[8][2][8] ), .ip2(\ANSWER/mem[9][2][8] ), 
        .s(n18137), .op(n18064) );
  mux2_1 U19013 ( .ip1(n18065), .ip2(n18064), .s(n18252), .op(n18066) );
  and2_1 U19014 ( .ip1(n18884), .ip2(n18066), .op(n18110) );
  mux2_1 U19015 ( .ip1(\ANSWER/mem[0][3][8] ), .ip2(\ANSWER/mem[1][3][8] ), 
        .s(n18137), .op(n18068) );
  mux2_1 U19016 ( .ip1(\ANSWER/mem[2][3][8] ), .ip2(\ANSWER/mem[3][3][8] ), 
        .s(n18137), .op(n18067) );
  mux2_1 U19017 ( .ip1(n18068), .ip2(n18067), .s(n18112), .op(n18072) );
  mux2_1 U19018 ( .ip1(\ANSWER/mem[4][3][8] ), .ip2(\ANSWER/mem[5][3][8] ), 
        .s(n18137), .op(n18070) );
  mux2_1 U19019 ( .ip1(\ANSWER/mem[6][3][8] ), .ip2(\ANSWER/mem[7][3][8] ), 
        .s(n18137), .op(n18069) );
  mux2_1 U19020 ( .ip1(n18070), .ip2(n18069), .s(n18112), .op(n18071) );
  mux2_1 U19021 ( .ip1(n18072), .ip2(n18071), .s(n18848), .op(n18075) );
  mux2_1 U19022 ( .ip1(\ANSWER/mem[8][3][8] ), .ip2(\ANSWER/mem[9][3][8] ), 
        .s(n18137), .op(n18074) );
  mux2_1 U19023 ( .ip1(n18075), .ip2(n18074), .s(n18073), .op(n18076) );
  nand2_1 U19024 ( .ip1(n18854), .ip2(n18076), .op(n18108) );
  mux2_1 U19025 ( .ip1(\ANSWER/mem[0][5][8] ), .ip2(\ANSWER/mem[1][5][8] ), 
        .s(n18137), .op(n18078) );
  mux2_1 U19026 ( .ip1(\ANSWER/mem[2][5][8] ), .ip2(\ANSWER/mem[3][5][8] ), 
        .s(n18143), .op(n18077) );
  mux2_1 U19027 ( .ip1(n18078), .ip2(n18077), .s(n18112), .op(n18082) );
  mux2_1 U19028 ( .ip1(\ANSWER/mem[4][5][8] ), .ip2(\ANSWER/mem[5][5][8] ), 
        .s(n18143), .op(n18080) );
  mux2_1 U19029 ( .ip1(\ANSWER/mem[6][5][8] ), .ip2(\ANSWER/mem[7][5][8] ), 
        .s(n18143), .op(n18079) );
  mux2_1 U19030 ( .ip1(n18080), .ip2(n18079), .s(n18112), .op(n18081) );
  mux2_1 U19031 ( .ip1(n18082), .ip2(n18081), .s(n18806), .op(n18084) );
  mux2_1 U19032 ( .ip1(\ANSWER/mem[8][5][8] ), .ip2(\ANSWER/mem[9][5][8] ), 
        .s(n18143), .op(n18083) );
  inv_1 U19033 ( .ip(n18165), .op(n18910) );
  mux2_1 U19034 ( .ip1(n18084), .ip2(n18083), .s(n18910), .op(n18085) );
  nand2_1 U19035 ( .ip1(n18832), .ip2(n18085), .op(n18107) );
  mux2_1 U19036 ( .ip1(\ANSWER/mem[0][7][8] ), .ip2(\ANSWER/mem[1][7][8] ), 
        .s(n18143), .op(n18087) );
  mux2_1 U19037 ( .ip1(\ANSWER/mem[2][7][8] ), .ip2(\ANSWER/mem[3][7][8] ), 
        .s(n18143), .op(n18086) );
  inv_1 U19038 ( .ip(n4366), .op(n18138) );
  mux2_1 U19039 ( .ip1(n18087), .ip2(n18086), .s(n18138), .op(n18091) );
  mux2_1 U19040 ( .ip1(\ANSWER/mem[4][7][8] ), .ip2(\ANSWER/mem[5][7][8] ), 
        .s(n18143), .op(n18089) );
  mux2_1 U19041 ( .ip1(\ANSWER/mem[6][7][8] ), .ip2(\ANSWER/mem[7][7][8] ), 
        .s(n18143), .op(n18088) );
  mux2_1 U19042 ( .ip1(n18089), .ip2(n18088), .s(n18138), .op(n18090) );
  mux2_1 U19043 ( .ip1(n18091), .ip2(n18090), .s(n18815), .op(n18094) );
  mux2_1 U19044 ( .ip1(\ANSWER/mem[8][7][8] ), .ip2(\ANSWER/mem[9][7][8] ), 
        .s(n18137), .op(n18093) );
  mux2_1 U19045 ( .ip1(n18094), .ip2(n18093), .s(n18092), .op(n18095) );
  nand2_1 U19046 ( .ip1(n18865), .ip2(n18095), .op(n18106) );
  mux2_1 U19047 ( .ip1(\ANSWER/mem[0][0][8] ), .ip2(\ANSWER/mem[1][0][8] ), 
        .s(n18137), .op(n18097) );
  mux2_1 U19048 ( .ip1(\ANSWER/mem[2][0][8] ), .ip2(\ANSWER/mem[3][0][8] ), 
        .s(n18900), .op(n18096) );
  mux2_1 U19049 ( .ip1(n18097), .ip2(n18096), .s(n18112), .op(n18101) );
  mux2_1 U19050 ( .ip1(\ANSWER/mem[4][0][8] ), .ip2(\ANSWER/mem[5][0][8] ), 
        .s(n18244), .op(n18099) );
  mux2_1 U19051 ( .ip1(\ANSWER/mem[6][0][8] ), .ip2(\ANSWER/mem[7][0][8] ), 
        .s(n18458), .op(n18098) );
  mux2_1 U19052 ( .ip1(n18099), .ip2(n18098), .s(n18112), .op(n18100) );
  mux2_1 U19053 ( .ip1(n18101), .ip2(n18100), .s(n18848), .op(n18103) );
  mux2_1 U19054 ( .ip1(\ANSWER/mem[8][0][8] ), .ip2(\ANSWER/mem[9][0][8] ), 
        .s(n17564), .op(n18102) );
  mux2_1 U19055 ( .ip1(n18103), .ip2(n18102), .s(n18174), .op(n18104) );
  nand2_1 U19056 ( .ip1(n18800), .ip2(n18104), .op(n18105) );
  nand4_1 U19057 ( .ip1(n18108), .ip2(n18107), .ip3(n18106), .ip4(n18105), 
        .op(n18109) );
  not_ab_or_c_or_d U19058 ( .ip1(n18872), .ip2(n18111), .ip3(n18110), .ip4(
        n18109), .op(n18123) );
  mux2_1 U19059 ( .ip1(\ANSWER/mem[0][6][8] ), .ip2(\ANSWER/mem[1][6][8] ), 
        .s(n18143), .op(n18114) );
  mux2_1 U19060 ( .ip1(\ANSWER/mem[2][6][8] ), .ip2(\ANSWER/mem[3][6][8] ), 
        .s(n18143), .op(n18113) );
  mux2_1 U19061 ( .ip1(n18114), .ip2(n18113), .s(n18112), .op(n18118) );
  mux2_1 U19062 ( .ip1(\ANSWER/mem[4][6][8] ), .ip2(\ANSWER/mem[5][6][8] ), 
        .s(n18143), .op(n18116) );
  mux2_1 U19063 ( .ip1(\ANSWER/mem[6][6][8] ), .ip2(\ANSWER/mem[7][6][8] ), 
        .s(n18143), .op(n18115) );
  mux2_1 U19064 ( .ip1(n18116), .ip2(n18115), .s(n18138), .op(n18117) );
  mux2_1 U19065 ( .ip1(n18118), .ip2(n18117), .s(n18848), .op(n18120) );
  mux2_1 U19066 ( .ip1(\ANSWER/mem[8][6][8] ), .ip2(\ANSWER/mem[9][6][8] ), 
        .s(n18143), .op(n18119) );
  inv_1 U19067 ( .ip(n18165), .op(n18679) );
  mux2_1 U19068 ( .ip1(n18120), .ip2(n18119), .s(n18679), .op(n18121) );
  nand2_1 U19069 ( .ip1(n18821), .ip2(n18121), .op(n18122) );
  nand3_1 U19070 ( .ip1(n18124), .ip2(n18123), .ip3(n18122), .op(n18125) );
  nand2_1 U19071 ( .ip1(n18125), .ip2(n18888), .op(n18149) );
  mux2_1 U19072 ( .ip1(\ANSWER/mem[0][9][8] ), .ip2(\ANSWER/mem[1][9][8] ), 
        .s(n18137), .op(n18127) );
  mux2_1 U19073 ( .ip1(\ANSWER/mem[2][9][8] ), .ip2(\ANSWER/mem[3][9][8] ), 
        .s(n18143), .op(n18126) );
  mux2_1 U19074 ( .ip1(n18127), .ip2(n18126), .s(n18138), .op(n18131) );
  mux2_1 U19075 ( .ip1(\ANSWER/mem[4][9][8] ), .ip2(\ANSWER/mem[5][9][8] ), 
        .s(n18143), .op(n18129) );
  mux2_1 U19076 ( .ip1(\ANSWER/mem[6][9][8] ), .ip2(\ANSWER/mem[7][9][8] ), 
        .s(n18143), .op(n18128) );
  mux2_1 U19077 ( .ip1(n18129), .ip2(n18128), .s(n18138), .op(n18130) );
  mux2_1 U19078 ( .ip1(n18131), .ip2(n18130), .s(n18837), .op(n18133) );
  mux2_1 U19079 ( .ip1(\ANSWER/mem[8][9][8] ), .ip2(\ANSWER/mem[9][9][8] ), 
        .s(n18143), .op(n18132) );
  mux2_1 U19080 ( .ip1(n18133), .ip2(n18132), .s(n18252), .op(n18134) );
  nand2_1 U19081 ( .ip1(n18899), .ip2(n18134), .op(n18148) );
  mux2_1 U19082 ( .ip1(\ANSWER/mem[0][8][8] ), .ip2(\ANSWER/mem[1][8][8] ), 
        .s(n18143), .op(n18136) );
  mux2_1 U19083 ( .ip1(\ANSWER/mem[2][8][8] ), .ip2(\ANSWER/mem[3][8][8] ), 
        .s(n18143), .op(n18135) );
  mux2_1 U19084 ( .ip1(n18136), .ip2(n18135), .s(n18138), .op(n18142) );
  mux2_1 U19085 ( .ip1(\ANSWER/mem[4][8][8] ), .ip2(\ANSWER/mem[5][8][8] ), 
        .s(n18137), .op(n18140) );
  mux2_1 U19086 ( .ip1(\ANSWER/mem[6][8][8] ), .ip2(\ANSWER/mem[7][8][8] ), 
        .s(n18143), .op(n18139) );
  mux2_1 U19087 ( .ip1(n18140), .ip2(n18139), .s(n18138), .op(n18141) );
  mux2_1 U19088 ( .ip1(n18142), .ip2(n18141), .s(n18815), .op(n18145) );
  mux2_1 U19089 ( .ip1(\ANSWER/mem[8][8][8] ), .ip2(\ANSWER/mem[9][8][8] ), 
        .s(n18143), .op(n18144) );
  mux2_1 U19090 ( .ip1(n18145), .ip2(n18144), .s(n18252), .op(n18146) );
  nand2_1 U19091 ( .ip1(n18914), .ip2(n18146), .op(n18147) );
  nand3_1 U19092 ( .ip1(n18149), .ip2(n18148), .ip3(n18147), .op(\ANSWER/N479 ) );
  mux2_1 U19093 ( .ip1(\ANSWER/mem[0][2][9] ), .ip2(\ANSWER/mem[1][2][9] ), 
        .s(n18616), .op(n18151) );
  mux2_1 U19094 ( .ip1(\ANSWER/mem[2][2][9] ), .ip2(\ANSWER/mem[3][2][9] ), 
        .s(n17711), .op(n18150) );
  mux2_1 U19095 ( .ip1(n18151), .ip2(n18150), .s(n15636), .op(n18155) );
  mux2_1 U19096 ( .ip1(\ANSWER/mem[4][2][9] ), .ip2(\ANSWER/mem[5][2][9] ), 
        .s(n17884), .op(n18153) );
  inv_1 U19097 ( .ip(n4362), .op(n18251) );
  buf_1 U19098 ( .ip(n18251), .op(n18244) );
  mux2_1 U19099 ( .ip1(\ANSWER/mem[6][2][9] ), .ip2(\ANSWER/mem[7][2][9] ), 
        .s(n18244), .op(n18152) );
  mux2_1 U19100 ( .ip1(n18153), .ip2(n18152), .s(n15636), .op(n18154) );
  mux2_1 U19101 ( .ip1(n18155), .ip2(n18154), .s(n18837), .op(n18157) );
  mux2_1 U19102 ( .ip1(\ANSWER/mem[8][2][9] ), .ip2(\ANSWER/mem[9][2][9] ), 
        .s(n18244), .op(n18156) );
  mux2_1 U19103 ( .ip1(n18157), .ip2(n18156), .s(n18252), .op(n18158) );
  nand2_1 U19104 ( .ip1(n18158), .ip2(n18884), .op(n18233) );
  mux2_1 U19105 ( .ip1(\ANSWER/mem[0][0][9] ), .ip2(\ANSWER/mem[1][0][9] ), 
        .s(n17921), .op(n18160) );
  mux2_1 U19106 ( .ip1(\ANSWER/mem[2][0][9] ), .ip2(\ANSWER/mem[3][0][9] ), 
        .s(n18244), .op(n18159) );
  mux2_1 U19107 ( .ip1(n18160), .ip2(n18159), .s(n15636), .op(n18164) );
  mux2_1 U19108 ( .ip1(\ANSWER/mem[4][0][9] ), .ip2(\ANSWER/mem[5][0][9] ), 
        .s(n17344), .op(n18162) );
  mux2_1 U19109 ( .ip1(\ANSWER/mem[6][0][9] ), .ip2(\ANSWER/mem[7][0][9] ), 
        .s(n18741), .op(n18161) );
  mux2_1 U19110 ( .ip1(n18162), .ip2(n18161), .s(n15636), .op(n18163) );
  mux2_1 U19111 ( .ip1(n18164), .ip2(n18163), .s(n18837), .op(n18167) );
  mux2_1 U19112 ( .ip1(\ANSWER/mem[8][0][9] ), .ip2(\ANSWER/mem[9][0][9] ), 
        .s(n17884), .op(n18166) );
  inv_1 U19113 ( .ip(n18165), .op(n18466) );
  mux2_1 U19114 ( .ip1(n18167), .ip2(n18166), .s(n18466), .op(n18220) );
  mux2_1 U19115 ( .ip1(\ANSWER/mem[0][6][9] ), .ip2(\ANSWER/mem[1][6][9] ), 
        .s(n18251), .op(n18169) );
  mux2_1 U19116 ( .ip1(\ANSWER/mem[2][6][9] ), .ip2(\ANSWER/mem[3][6][9] ), 
        .s(n18251), .op(n18168) );
  mux2_1 U19117 ( .ip1(n18169), .ip2(n18168), .s(n17581), .op(n18173) );
  mux2_1 U19118 ( .ip1(\ANSWER/mem[4][6][9] ), .ip2(\ANSWER/mem[5][6][9] ), 
        .s(n18251), .op(n18171) );
  mux2_1 U19119 ( .ip1(\ANSWER/mem[6][6][9] ), .ip2(\ANSWER/mem[7][6][9] ), 
        .s(n18251), .op(n18170) );
  mux2_1 U19120 ( .ip1(n18171), .ip2(n18170), .s(n17990), .op(n18172) );
  mux2_1 U19121 ( .ip1(n18173), .ip2(n18172), .s(n18837), .op(n18176) );
  mux2_1 U19122 ( .ip1(\ANSWER/mem[8][6][9] ), .ip2(\ANSWER/mem[9][6][9] ), 
        .s(n18251), .op(n18175) );
  mux2_1 U19123 ( .ip1(n18176), .ip2(n18175), .s(n18174), .op(n18177) );
  and2_1 U19124 ( .ip1(n18821), .ip2(n18177), .op(n18219) );
  mux2_1 U19125 ( .ip1(\ANSWER/mem[0][7][9] ), .ip2(\ANSWER/mem[1][7][9] ), 
        .s(n18251), .op(n18179) );
  mux2_1 U19126 ( .ip1(\ANSWER/mem[2][7][9] ), .ip2(\ANSWER/mem[3][7][9] ), 
        .s(n18251), .op(n18178) );
  mux2_1 U19127 ( .ip1(n18179), .ip2(n18178), .s(n18330), .op(n18183) );
  mux2_1 U19128 ( .ip1(\ANSWER/mem[4][7][9] ), .ip2(\ANSWER/mem[5][7][9] ), 
        .s(n18251), .op(n18181) );
  mux2_1 U19129 ( .ip1(\ANSWER/mem[6][7][9] ), .ip2(\ANSWER/mem[7][7][9] ), 
        .s(n18251), .op(n18180) );
  mux2_1 U19130 ( .ip1(n18181), .ip2(n18180), .s(n17990), .op(n18182) );
  mux2_1 U19131 ( .ip1(n18183), .ip2(n18182), .s(n18837), .op(n18185) );
  mux2_1 U19132 ( .ip1(\ANSWER/mem[8][7][9] ), .ip2(\ANSWER/mem[9][7][9] ), 
        .s(n18251), .op(n18184) );
  mux2_1 U19133 ( .ip1(n18185), .ip2(n18184), .s(n18679), .op(n18186) );
  nand2_1 U19134 ( .ip1(n18865), .ip2(n18186), .op(n18217) );
  mux2_1 U19135 ( .ip1(\ANSWER/mem[0][1][9] ), .ip2(\ANSWER/mem[1][1][9] ), 
        .s(n17344), .op(n18188) );
  mux2_1 U19136 ( .ip1(\ANSWER/mem[2][1][9] ), .ip2(\ANSWER/mem[3][1][9] ), 
        .s(n17533), .op(n18187) );
  mux2_1 U19137 ( .ip1(n18188), .ip2(n18187), .s(n18112), .op(n18192) );
  mux2_1 U19138 ( .ip1(\ANSWER/mem[4][1][9] ), .ip2(\ANSWER/mem[5][1][9] ), 
        .s(n18029), .op(n18190) );
  mux2_1 U19139 ( .ip1(\ANSWER/mem[6][1][9] ), .ip2(\ANSWER/mem[7][1][9] ), 
        .s(n17817), .op(n18189) );
  mux2_1 U19140 ( .ip1(n18190), .ip2(n18189), .s(n18544), .op(n18191) );
  mux2_1 U19141 ( .ip1(n18192), .ip2(n18191), .s(n18837), .op(n18194) );
  mux2_1 U19142 ( .ip1(\ANSWER/mem[8][1][9] ), .ip2(\ANSWER/mem[9][1][9] ), 
        .s(n18616), .op(n18193) );
  mux2_1 U19143 ( .ip1(n18194), .ip2(n18193), .s(n18910), .op(n18195) );
  nand2_1 U19144 ( .ip1(n18872), .ip2(n18195), .op(n18216) );
  mux2_1 U19145 ( .ip1(\ANSWER/mem[0][3][9] ), .ip2(\ANSWER/mem[1][3][9] ), 
        .s(n18244), .op(n18197) );
  mux2_1 U19146 ( .ip1(\ANSWER/mem[2][3][9] ), .ip2(\ANSWER/mem[3][3][9] ), 
        .s(n18244), .op(n18196) );
  mux2_1 U19147 ( .ip1(n18197), .ip2(n18196), .s(n18330), .op(n18201) );
  mux2_1 U19148 ( .ip1(\ANSWER/mem[4][3][9] ), .ip2(\ANSWER/mem[5][3][9] ), 
        .s(n18244), .op(n18199) );
  mux2_1 U19149 ( .ip1(\ANSWER/mem[6][3][9] ), .ip2(\ANSWER/mem[7][3][9] ), 
        .s(n18244), .op(n18198) );
  mux2_1 U19150 ( .ip1(n18199), .ip2(n18198), .s(n18435), .op(n18200) );
  mux2_1 U19151 ( .ip1(n18201), .ip2(n18200), .s(n18837), .op(n18203) );
  mux2_1 U19152 ( .ip1(\ANSWER/mem[8][3][9] ), .ip2(\ANSWER/mem[9][3][9] ), 
        .s(n18244), .op(n18202) );
  mux2_1 U19153 ( .ip1(n18203), .ip2(n18202), .s(n18227), .op(n18204) );
  nand2_1 U19154 ( .ip1(n18854), .ip2(n18204), .op(n18215) );
  mux2_1 U19155 ( .ip1(\ANSWER/mem[0][4][9] ), .ip2(\ANSWER/mem[1][4][9] ), 
        .s(n18244), .op(n18206) );
  mux2_1 U19156 ( .ip1(\ANSWER/mem[2][4][9] ), .ip2(\ANSWER/mem[3][4][9] ), 
        .s(n18244), .op(n18205) );
  mux2_1 U19157 ( .ip1(n18206), .ip2(n18205), .s(n18138), .op(n18210) );
  mux2_1 U19158 ( .ip1(\ANSWER/mem[4][4][9] ), .ip2(\ANSWER/mem[5][4][9] ), 
        .s(n18244), .op(n18208) );
  mux2_1 U19159 ( .ip1(\ANSWER/mem[6][4][9] ), .ip2(\ANSWER/mem[7][4][9] ), 
        .s(n18244), .op(n18207) );
  mux2_1 U19160 ( .ip1(n18208), .ip2(n18207), .s(n18354), .op(n18209) );
  mux2_1 U19161 ( .ip1(n18210), .ip2(n18209), .s(n18837), .op(n18212) );
  mux2_1 U19162 ( .ip1(\ANSWER/mem[8][4][9] ), .ip2(\ANSWER/mem[9][4][9] ), 
        .s(n18244), .op(n18211) );
  mux2_1 U19163 ( .ip1(n18212), .ip2(n18211), .s(n18466), .op(n18213) );
  nand2_1 U19164 ( .ip1(n18843), .ip2(n18213), .op(n18214) );
  nand4_1 U19165 ( .ip1(n18217), .ip2(n18216), .ip3(n18215), .ip4(n18214), 
        .op(n18218) );
  not_ab_or_c_or_d U19166 ( .ip1(n18220), .ip2(n18800), .ip3(n18219), .ip4(
        n18218), .op(n18232) );
  mux2_1 U19167 ( .ip1(\ANSWER/mem[0][5][9] ), .ip2(\ANSWER/mem[1][5][9] ), 
        .s(n18244), .op(n18222) );
  mux2_1 U19168 ( .ip1(\ANSWER/mem[2][5][9] ), .ip2(\ANSWER/mem[3][5][9] ), 
        .s(n18251), .op(n18221) );
  mux2_1 U19169 ( .ip1(n18222), .ip2(n18221), .s(n15636), .op(n18226) );
  mux2_1 U19170 ( .ip1(\ANSWER/mem[4][5][9] ), .ip2(\ANSWER/mem[5][5][9] ), 
        .s(n18251), .op(n18224) );
  mux2_1 U19171 ( .ip1(\ANSWER/mem[6][5][9] ), .ip2(\ANSWER/mem[7][5][9] ), 
        .s(n18251), .op(n18223) );
  mux2_1 U19172 ( .ip1(n18224), .ip2(n18223), .s(n15636), .op(n18225) );
  mux2_1 U19173 ( .ip1(n18226), .ip2(n18225), .s(n18837), .op(n18229) );
  mux2_1 U19174 ( .ip1(\ANSWER/mem[8][5][9] ), .ip2(\ANSWER/mem[9][5][9] ), 
        .s(n18251), .op(n18228) );
  mux2_1 U19175 ( .ip1(n18229), .ip2(n18228), .s(n18227), .op(n18230) );
  nand2_1 U19176 ( .ip1(n18832), .ip2(n18230), .op(n18231) );
  nand3_1 U19177 ( .ip1(n18233), .ip2(n18232), .ip3(n18231), .op(n18234) );
  nand2_1 U19178 ( .ip1(n18234), .ip2(n18888), .op(n18258) );
  mux2_1 U19179 ( .ip1(\ANSWER/mem[0][9][9] ), .ip2(\ANSWER/mem[1][9][9] ), 
        .s(n18251), .op(n18236) );
  mux2_1 U19180 ( .ip1(\ANSWER/mem[2][9][9] ), .ip2(\ANSWER/mem[3][9][9] ), 
        .s(n18244), .op(n18235) );
  mux2_1 U19181 ( .ip1(n18236), .ip2(n18235), .s(n17366), .op(n18240) );
  mux2_1 U19182 ( .ip1(\ANSWER/mem[4][9][9] ), .ip2(\ANSWER/mem[5][9][9] ), 
        .s(n18251), .op(n18238) );
  mux2_1 U19183 ( .ip1(\ANSWER/mem[6][9][9] ), .ip2(\ANSWER/mem[7][9][9] ), 
        .s(n18251), .op(n18237) );
  mux2_1 U19184 ( .ip1(n18238), .ip2(n18237), .s(n17605), .op(n18239) );
  mux2_1 U19185 ( .ip1(n18240), .ip2(n18239), .s(n18837), .op(n18242) );
  mux2_1 U19186 ( .ip1(\ANSWER/mem[8][9][9] ), .ip2(\ANSWER/mem[9][9][9] ), 
        .s(n18251), .op(n18241) );
  mux2_1 U19187 ( .ip1(n18242), .ip2(n18241), .s(n18252), .op(n18243) );
  nand2_1 U19188 ( .ip1(n18899), .ip2(n18243), .op(n18257) );
  mux2_1 U19189 ( .ip1(\ANSWER/mem[0][8][9] ), .ip2(\ANSWER/mem[1][8][9] ), 
        .s(n18244), .op(n18246) );
  mux2_1 U19190 ( .ip1(\ANSWER/mem[2][8][9] ), .ip2(\ANSWER/mem[3][8][9] ), 
        .s(n18244), .op(n18245) );
  mux2_1 U19191 ( .ip1(n18246), .ip2(n18245), .s(n18112), .op(n18250) );
  mux2_1 U19192 ( .ip1(\ANSWER/mem[4][8][9] ), .ip2(\ANSWER/mem[5][8][9] ), 
        .s(n18251), .op(n18248) );
  mux2_1 U19193 ( .ip1(\ANSWER/mem[6][8][9] ), .ip2(\ANSWER/mem[7][8][9] ), 
        .s(n18251), .op(n18247) );
  mux2_1 U19194 ( .ip1(n18248), .ip2(n18247), .s(n15636), .op(n18249) );
  mux2_1 U19195 ( .ip1(n18250), .ip2(n18249), .s(n18837), .op(n18254) );
  mux2_1 U19196 ( .ip1(\ANSWER/mem[8][8][9] ), .ip2(\ANSWER/mem[9][8][9] ), 
        .s(n18251), .op(n18253) );
  mux2_1 U19197 ( .ip1(n18254), .ip2(n18253), .s(n18252), .op(n18255) );
  nand2_1 U19198 ( .ip1(n18914), .ip2(n18255), .op(n18256) );
  nand3_1 U19199 ( .ip1(n18258), .ip2(n18257), .ip3(n18256), .op(\ANSWER/N478 ) );
  mux2_1 U19200 ( .ip1(\ANSWER/mem[0][0][10] ), .ip2(\ANSWER/mem[1][0][10] ), 
        .s(n18741), .op(n18260) );
  mux2_1 U19201 ( .ip1(\ANSWER/mem[2][0][10] ), .ip2(\ANSWER/mem[3][0][10] ), 
        .s(n18900), .op(n18259) );
  inv_1 U19202 ( .ip(n4366), .op(n18330) );
  mux2_1 U19203 ( .ip1(n18260), .ip2(n18259), .s(n18330), .op(n18264) );
  mux2_1 U19204 ( .ip1(\ANSWER/mem[4][0][10] ), .ip2(\ANSWER/mem[5][0][10] ), 
        .s(n18029), .op(n18262) );
  mux2_1 U19205 ( .ip1(\ANSWER/mem[6][0][10] ), .ip2(\ANSWER/mem[7][0][10] ), 
        .s(n17344), .op(n18261) );
  mux2_1 U19206 ( .ip1(n18262), .ip2(n18261), .s(n18330), .op(n18263) );
  mux2_1 U19207 ( .ip1(n18264), .ip2(n18263), .s(n18806), .op(n18266) );
  mux2_1 U19208 ( .ip1(\ANSWER/mem[8][0][10] ), .ip2(\ANSWER/mem[9][0][10] ), 
        .s(n18741), .op(n18265) );
  mux2_1 U19209 ( .ip1(n18266), .ip2(n18265), .s(n18466), .op(n18267) );
  nand2_1 U19210 ( .ip1(n18267), .ip2(n18800), .op(n18340) );
  inv_1 U19211 ( .ip(n4362), .op(n18359) );
  mux2_1 U19212 ( .ip1(\ANSWER/mem[0][5][10] ), .ip2(\ANSWER/mem[1][5][10] ), 
        .s(n18359), .op(n18269) );
  buf_1 U19213 ( .ip(n18359), .op(n18351) );
  mux2_1 U19214 ( .ip1(\ANSWER/mem[2][5][10] ), .ip2(\ANSWER/mem[3][5][10] ), 
        .s(n18351), .op(n18268) );
  mux2_1 U19215 ( .ip1(n18269), .ip2(n18268), .s(n18330), .op(n18273) );
  mux2_1 U19216 ( .ip1(\ANSWER/mem[4][5][10] ), .ip2(\ANSWER/mem[5][5][10] ), 
        .s(n18351), .op(n18271) );
  mux2_1 U19217 ( .ip1(\ANSWER/mem[6][5][10] ), .ip2(\ANSWER/mem[7][5][10] ), 
        .s(n18351), .op(n18270) );
  mux2_1 U19218 ( .ip1(n18271), .ip2(n18270), .s(n18330), .op(n18272) );
  mux2_1 U19219 ( .ip1(n18273), .ip2(n18272), .s(n18806), .op(n18275) );
  mux2_1 U19220 ( .ip1(\ANSWER/mem[8][5][10] ), .ip2(\ANSWER/mem[9][5][10] ), 
        .s(n18351), .op(n18274) );
  mux2_1 U19221 ( .ip1(n18275), .ip2(n18274), .s(n18466), .op(n18327) );
  mux2_1 U19222 ( .ip1(\ANSWER/mem[0][6][10] ), .ip2(\ANSWER/mem[1][6][10] ), 
        .s(n18351), .op(n18277) );
  mux2_1 U19223 ( .ip1(\ANSWER/mem[2][6][10] ), .ip2(\ANSWER/mem[3][6][10] ), 
        .s(n18351), .op(n18276) );
  mux2_1 U19224 ( .ip1(n18277), .ip2(n18276), .s(n18330), .op(n18281) );
  mux2_1 U19225 ( .ip1(\ANSWER/mem[4][6][10] ), .ip2(\ANSWER/mem[5][6][10] ), 
        .s(n18351), .op(n18279) );
  mux2_1 U19226 ( .ip1(\ANSWER/mem[6][6][10] ), .ip2(\ANSWER/mem[7][6][10] ), 
        .s(n18351), .op(n18278) );
  inv_1 U19227 ( .ip(n4366), .op(n18354) );
  mux2_1 U19228 ( .ip1(n18279), .ip2(n18278), .s(n18354), .op(n18280) );
  mux2_1 U19229 ( .ip1(n18281), .ip2(n18280), .s(n18806), .op(n18283) );
  mux2_1 U19230 ( .ip1(\ANSWER/mem[8][6][10] ), .ip2(\ANSWER/mem[9][6][10] ), 
        .s(n18351), .op(n18282) );
  mux2_1 U19231 ( .ip1(n18283), .ip2(n18282), .s(n18466), .op(n18284) );
  and2_1 U19232 ( .ip1(n18821), .ip2(n18284), .op(n18326) );
  mux2_1 U19233 ( .ip1(\ANSWER/mem[0][3][10] ), .ip2(\ANSWER/mem[1][3][10] ), 
        .s(n18359), .op(n18286) );
  mux2_1 U19234 ( .ip1(\ANSWER/mem[2][3][10] ), .ip2(\ANSWER/mem[3][3][10] ), 
        .s(n18359), .op(n18285) );
  mux2_1 U19235 ( .ip1(n18286), .ip2(n18285), .s(n18330), .op(n18290) );
  mux2_1 U19236 ( .ip1(\ANSWER/mem[4][3][10] ), .ip2(\ANSWER/mem[5][3][10] ), 
        .s(n18359), .op(n18288) );
  mux2_1 U19237 ( .ip1(\ANSWER/mem[6][3][10] ), .ip2(\ANSWER/mem[7][3][10] ), 
        .s(n18359), .op(n18287) );
  mux2_1 U19238 ( .ip1(n18288), .ip2(n18287), .s(n18330), .op(n18289) );
  mux2_1 U19239 ( .ip1(n18290), .ip2(n18289), .s(n18837), .op(n18292) );
  mux2_1 U19240 ( .ip1(\ANSWER/mem[8][3][10] ), .ip2(\ANSWER/mem[9][3][10] ), 
        .s(n18359), .op(n18291) );
  mux2_1 U19241 ( .ip1(n18292), .ip2(n18291), .s(n18466), .op(n18293) );
  nand2_1 U19242 ( .ip1(n18854), .ip2(n18293), .op(n18324) );
  mux2_1 U19243 ( .ip1(\ANSWER/mem[0][2][10] ), .ip2(\ANSWER/mem[1][2][10] ), 
        .s(n17884), .op(n18295) );
  mux2_1 U19244 ( .ip1(\ANSWER/mem[2][2][10] ), .ip2(\ANSWER/mem[3][2][10] ), 
        .s(n17387), .op(n18294) );
  mux2_1 U19245 ( .ip1(n18295), .ip2(n18294), .s(n18330), .op(n18299) );
  mux2_1 U19246 ( .ip1(\ANSWER/mem[4][2][10] ), .ip2(\ANSWER/mem[5][2][10] ), 
        .s(n17711), .op(n18297) );
  mux2_1 U19247 ( .ip1(\ANSWER/mem[6][2][10] ), .ip2(\ANSWER/mem[7][2][10] ), 
        .s(n18359), .op(n18296) );
  mux2_1 U19248 ( .ip1(n18297), .ip2(n18296), .s(n18330), .op(n18298) );
  mux2_1 U19249 ( .ip1(n18299), .ip2(n18298), .s(n18906), .op(n18301) );
  mux2_1 U19250 ( .ip1(\ANSWER/mem[8][2][10] ), .ip2(\ANSWER/mem[9][2][10] ), 
        .s(n18359), .op(n18300) );
  mux2_1 U19251 ( .ip1(n18301), .ip2(n18300), .s(n18466), .op(n18302) );
  nand2_1 U19252 ( .ip1(n18884), .ip2(n18302), .op(n18323) );
  mux2_1 U19253 ( .ip1(\ANSWER/mem[0][4][10] ), .ip2(\ANSWER/mem[1][4][10] ), 
        .s(n18359), .op(n18304) );
  mux2_1 U19254 ( .ip1(\ANSWER/mem[2][4][10] ), .ip2(\ANSWER/mem[3][4][10] ), 
        .s(n18359), .op(n18303) );
  mux2_1 U19255 ( .ip1(n18304), .ip2(n18303), .s(n18330), .op(n18308) );
  mux2_1 U19256 ( .ip1(\ANSWER/mem[4][4][10] ), .ip2(\ANSWER/mem[5][4][10] ), 
        .s(n18359), .op(n18306) );
  mux2_1 U19257 ( .ip1(\ANSWER/mem[6][4][10] ), .ip2(\ANSWER/mem[7][4][10] ), 
        .s(n18359), .op(n18305) );
  mux2_1 U19258 ( .ip1(n18306), .ip2(n18305), .s(n18330), .op(n18307) );
  mux2_1 U19259 ( .ip1(n18308), .ip2(n18307), .s(n18806), .op(n18310) );
  mux2_1 U19260 ( .ip1(\ANSWER/mem[8][4][10] ), .ip2(\ANSWER/mem[9][4][10] ), 
        .s(n18359), .op(n18309) );
  mux2_1 U19261 ( .ip1(n18310), .ip2(n18309), .s(n18466), .op(n18311) );
  nand2_1 U19262 ( .ip1(n18843), .ip2(n18311), .op(n18322) );
  mux2_1 U19263 ( .ip1(\ANSWER/mem[0][7][10] ), .ip2(\ANSWER/mem[1][7][10] ), 
        .s(n18351), .op(n18313) );
  mux2_1 U19264 ( .ip1(\ANSWER/mem[2][7][10] ), .ip2(\ANSWER/mem[3][7][10] ), 
        .s(n18351), .op(n18312) );
  mux2_1 U19265 ( .ip1(n18313), .ip2(n18312), .s(n18354), .op(n18317) );
  mux2_1 U19266 ( .ip1(\ANSWER/mem[4][7][10] ), .ip2(\ANSWER/mem[5][7][10] ), 
        .s(n18351), .op(n18315) );
  mux2_1 U19267 ( .ip1(\ANSWER/mem[6][7][10] ), .ip2(\ANSWER/mem[7][7][10] ), 
        .s(n18351), .op(n18314) );
  mux2_1 U19268 ( .ip1(n18315), .ip2(n18314), .s(n18354), .op(n18316) );
  mux2_1 U19269 ( .ip1(n18317), .ip2(n18316), .s(n18837), .op(n18319) );
  mux2_1 U19270 ( .ip1(\ANSWER/mem[8][7][10] ), .ip2(\ANSWER/mem[9][7][10] ), 
        .s(n18359), .op(n18318) );
  mux2_1 U19271 ( .ip1(n18319), .ip2(n18318), .s(n18466), .op(n18320) );
  nand2_1 U19272 ( .ip1(n18865), .ip2(n18320), .op(n18321) );
  nand4_1 U19273 ( .ip1(n18324), .ip2(n18323), .ip3(n18322), .ip4(n18321), 
        .op(n18325) );
  not_ab_or_c_or_d U19274 ( .ip1(n18327), .ip2(n18832), .ip3(n18326), .ip4(
        n18325), .op(n18339) );
  mux2_1 U19275 ( .ip1(\ANSWER/mem[0][1][10] ), .ip2(\ANSWER/mem[1][1][10] ), 
        .s(n18900), .op(n18329) );
  mux2_1 U19276 ( .ip1(\ANSWER/mem[2][1][10] ), .ip2(\ANSWER/mem[3][1][10] ), 
        .s(n17344), .op(n18328) );
  mux2_1 U19277 ( .ip1(n18329), .ip2(n18328), .s(n18330), .op(n18334) );
  mux2_1 U19278 ( .ip1(\ANSWER/mem[4][1][10] ), .ip2(\ANSWER/mem[5][1][10] ), 
        .s(n17884), .op(n18332) );
  mux2_1 U19279 ( .ip1(\ANSWER/mem[6][1][10] ), .ip2(\ANSWER/mem[7][1][10] ), 
        .s(n18244), .op(n18331) );
  mux2_1 U19280 ( .ip1(n18332), .ip2(n18331), .s(n18330), .op(n18333) );
  mux2_1 U19281 ( .ip1(n18334), .ip2(n18333), .s(n18859), .op(n18336) );
  mux2_1 U19282 ( .ip1(\ANSWER/mem[8][1][10] ), .ip2(\ANSWER/mem[9][1][10] ), 
        .s(n17387), .op(n18335) );
  mux2_1 U19283 ( .ip1(n18336), .ip2(n18335), .s(n18466), .op(n18337) );
  nand2_1 U19284 ( .ip1(n18872), .ip2(n18337), .op(n18338) );
  nand3_1 U19285 ( .ip1(n18340), .ip2(n18339), .ip3(n18338), .op(n18341) );
  nand2_1 U19286 ( .ip1(n18341), .ip2(n18888), .op(n18365) );
  mux2_1 U19287 ( .ip1(\ANSWER/mem[0][9][10] ), .ip2(\ANSWER/mem[1][9][10] ), 
        .s(n18359), .op(n18343) );
  mux2_1 U19288 ( .ip1(\ANSWER/mem[2][9][10] ), .ip2(\ANSWER/mem[3][9][10] ), 
        .s(n18351), .op(n18342) );
  mux2_1 U19289 ( .ip1(n18343), .ip2(n18342), .s(n18354), .op(n18347) );
  mux2_1 U19290 ( .ip1(\ANSWER/mem[4][9][10] ), .ip2(\ANSWER/mem[5][9][10] ), 
        .s(n18359), .op(n18345) );
  mux2_1 U19291 ( .ip1(\ANSWER/mem[6][9][10] ), .ip2(\ANSWER/mem[7][9][10] ), 
        .s(n18359), .op(n18344) );
  mux2_1 U19292 ( .ip1(n18345), .ip2(n18344), .s(n18354), .op(n18346) );
  mux2_1 U19293 ( .ip1(n18347), .ip2(n18346), .s(n18848), .op(n18349) );
  mux2_1 U19294 ( .ip1(\ANSWER/mem[8][9][10] ), .ip2(\ANSWER/mem[9][9][10] ), 
        .s(n18359), .op(n18348) );
  mux2_1 U19295 ( .ip1(n18349), .ip2(n18348), .s(n18466), .op(n18350) );
  nand2_1 U19296 ( .ip1(n18899), .ip2(n18350), .op(n18364) );
  mux2_1 U19297 ( .ip1(\ANSWER/mem[0][8][10] ), .ip2(\ANSWER/mem[1][8][10] ), 
        .s(n18351), .op(n18353) );
  mux2_1 U19298 ( .ip1(\ANSWER/mem[2][8][10] ), .ip2(\ANSWER/mem[3][8][10] ), 
        .s(n18351), .op(n18352) );
  mux2_1 U19299 ( .ip1(n18353), .ip2(n18352), .s(n18354), .op(n18358) );
  mux2_1 U19300 ( .ip1(\ANSWER/mem[4][8][10] ), .ip2(\ANSWER/mem[5][8][10] ), 
        .s(n18359), .op(n18356) );
  mux2_1 U19301 ( .ip1(\ANSWER/mem[6][8][10] ), .ip2(\ANSWER/mem[7][8][10] ), 
        .s(n18359), .op(n18355) );
  mux2_1 U19302 ( .ip1(n18356), .ip2(n18355), .s(n18354), .op(n18357) );
  mux2_1 U19303 ( .ip1(n18358), .ip2(n18357), .s(n18878), .op(n18361) );
  mux2_1 U19304 ( .ip1(\ANSWER/mem[8][8][10] ), .ip2(\ANSWER/mem[9][8][10] ), 
        .s(n18359), .op(n18360) );
  mux2_1 U19305 ( .ip1(n18361), .ip2(n18360), .s(n18466), .op(n18362) );
  nand2_1 U19306 ( .ip1(n18914), .ip2(n18362), .op(n18363) );
  nand3_1 U19307 ( .ip1(n18365), .ip2(n18364), .ip3(n18363), .op(\ANSWER/N477 ) );
  mux2_1 U19308 ( .ip1(\ANSWER/mem[0][0][11] ), .ip2(\ANSWER/mem[1][0][11] ), 
        .s(n17817), .op(n18367) );
  mux2_1 U19309 ( .ip1(\ANSWER/mem[2][0][11] ), .ip2(\ANSWER/mem[3][0][11] ), 
        .s(n18741), .op(n18366) );
  inv_1 U19310 ( .ip(n4366), .op(n18435) );
  mux2_1 U19311 ( .ip1(n18367), .ip2(n18366), .s(n18435), .op(n18371) );
  mux2_1 U19312 ( .ip1(\ANSWER/mem[4][0][11] ), .ip2(\ANSWER/mem[5][0][11] ), 
        .s(n18565), .op(n18369) );
  mux2_1 U19313 ( .ip1(\ANSWER/mem[6][0][11] ), .ip2(\ANSWER/mem[7][0][11] ), 
        .s(n18616), .op(n18368) );
  mux2_1 U19314 ( .ip1(n18369), .ip2(n18368), .s(n18435), .op(n18370) );
  mux2_1 U19315 ( .ip1(n18371), .ip2(n18370), .s(n18906), .op(n18373) );
  mux2_1 U19316 ( .ip1(\ANSWER/mem[8][0][11] ), .ip2(\ANSWER/mem[9][0][11] ), 
        .s(n17921), .op(n18372) );
  mux2_1 U19317 ( .ip1(n18373), .ip2(n18372), .s(n18466), .op(n18374) );
  nand2_1 U19318 ( .ip1(n18800), .ip2(n18374), .op(n18447) );
  mux2_1 U19319 ( .ip1(\ANSWER/mem[0][2][11] ), .ip2(\ANSWER/mem[1][2][11] ), 
        .s(n18741), .op(n18376) );
  mux2_1 U19320 ( .ip1(\ANSWER/mem[2][2][11] ), .ip2(\ANSWER/mem[3][2][11] ), 
        .s(n18244), .op(n18375) );
  mux2_1 U19321 ( .ip1(n18376), .ip2(n18375), .s(n18435), .op(n18380) );
  mux2_1 U19322 ( .ip1(\ANSWER/mem[4][2][11] ), .ip2(\ANSWER/mem[5][2][11] ), 
        .s(n17884), .op(n18378) );
  inv_1 U19323 ( .ip(n4362), .op(n18465) );
  mux2_1 U19324 ( .ip1(\ANSWER/mem[6][2][11] ), .ip2(\ANSWER/mem[7][2][11] ), 
        .s(n18465), .op(n18377) );
  mux2_1 U19325 ( .ip1(n18378), .ip2(n18377), .s(n18435), .op(n18379) );
  mux2_1 U19326 ( .ip1(n18380), .ip2(n18379), .s(n18906), .op(n18382) );
  mux2_1 U19327 ( .ip1(\ANSWER/mem[8][2][11] ), .ip2(\ANSWER/mem[9][2][11] ), 
        .s(n18465), .op(n18381) );
  mux2_1 U19328 ( .ip1(n18382), .ip2(n18381), .s(n18466), .op(n18434) );
  mux2_1 U19329 ( .ip1(\ANSWER/mem[0][4][11] ), .ip2(\ANSWER/mem[1][4][11] ), 
        .s(n18465), .op(n18384) );
  mux2_1 U19330 ( .ip1(\ANSWER/mem[2][4][11] ), .ip2(\ANSWER/mem[3][4][11] ), 
        .s(n18465), .op(n18383) );
  mux2_1 U19331 ( .ip1(n18384), .ip2(n18383), .s(n18435), .op(n18388) );
  mux2_1 U19332 ( .ip1(\ANSWER/mem[4][4][11] ), .ip2(\ANSWER/mem[5][4][11] ), 
        .s(n18465), .op(n18386) );
  mux2_1 U19333 ( .ip1(\ANSWER/mem[6][4][11] ), .ip2(\ANSWER/mem[7][4][11] ), 
        .s(n18465), .op(n18385) );
  mux2_1 U19334 ( .ip1(n18386), .ip2(n18385), .s(n18435), .op(n18387) );
  mux2_1 U19335 ( .ip1(n18388), .ip2(n18387), .s(n18906), .op(n18390) );
  mux2_1 U19336 ( .ip1(\ANSWER/mem[8][4][11] ), .ip2(\ANSWER/mem[9][4][11] ), 
        .s(n18465), .op(n18389) );
  mux2_1 U19337 ( .ip1(n18390), .ip2(n18389), .s(n18466), .op(n18391) );
  and2_1 U19338 ( .ip1(n18843), .ip2(n18391), .op(n18433) );
  mux2_1 U19339 ( .ip1(\ANSWER/mem[0][1][11] ), .ip2(\ANSWER/mem[1][1][11] ), 
        .s(n18616), .op(n18393) );
  mux2_1 U19340 ( .ip1(\ANSWER/mem[2][1][11] ), .ip2(\ANSWER/mem[3][1][11] ), 
        .s(n17921), .op(n18392) );
  mux2_1 U19341 ( .ip1(n18393), .ip2(n18392), .s(n18435), .op(n18397) );
  mux2_1 U19342 ( .ip1(\ANSWER/mem[4][1][11] ), .ip2(\ANSWER/mem[5][1][11] ), 
        .s(n17884), .op(n18395) );
  mux2_1 U19343 ( .ip1(\ANSWER/mem[6][1][11] ), .ip2(\ANSWER/mem[7][1][11] ), 
        .s(n17344), .op(n18394) );
  mux2_1 U19344 ( .ip1(n18395), .ip2(n18394), .s(n18435), .op(n18396) );
  mux2_1 U19345 ( .ip1(n18397), .ip2(n18396), .s(n18906), .op(n18399) );
  mux2_1 U19346 ( .ip1(\ANSWER/mem[8][1][11] ), .ip2(\ANSWER/mem[9][1][11] ), 
        .s(n17817), .op(n18398) );
  mux2_1 U19347 ( .ip1(n18399), .ip2(n18398), .s(n18466), .op(n18400) );
  nand2_1 U19348 ( .ip1(n18872), .ip2(n18400), .op(n18431) );
  mux2_1 U19349 ( .ip1(\ANSWER/mem[0][5][11] ), .ip2(\ANSWER/mem[1][5][11] ), 
        .s(n18465), .op(n18402) );
  buf_1 U19350 ( .ip(n18465), .op(n18458) );
  mux2_1 U19351 ( .ip1(\ANSWER/mem[2][5][11] ), .ip2(\ANSWER/mem[3][5][11] ), 
        .s(n18458), .op(n18401) );
  mux2_1 U19352 ( .ip1(n18402), .ip2(n18401), .s(n18435), .op(n18406) );
  mux2_1 U19353 ( .ip1(\ANSWER/mem[4][5][11] ), .ip2(\ANSWER/mem[5][5][11] ), 
        .s(n18458), .op(n18404) );
  mux2_1 U19354 ( .ip1(\ANSWER/mem[6][5][11] ), .ip2(\ANSWER/mem[7][5][11] ), 
        .s(n18458), .op(n18403) );
  mux2_1 U19355 ( .ip1(n18404), .ip2(n18403), .s(n18435), .op(n18405) );
  mux2_1 U19356 ( .ip1(n18406), .ip2(n18405), .s(n18906), .op(n18408) );
  mux2_1 U19357 ( .ip1(\ANSWER/mem[8][5][11] ), .ip2(\ANSWER/mem[9][5][11] ), 
        .s(n18458), .op(n18407) );
  mux2_1 U19358 ( .ip1(n18408), .ip2(n18407), .s(n18466), .op(n18409) );
  nand2_1 U19359 ( .ip1(n18832), .ip2(n18409), .op(n18430) );
  mux2_1 U19360 ( .ip1(\ANSWER/mem[0][3][11] ), .ip2(\ANSWER/mem[1][3][11] ), 
        .s(n18465), .op(n18411) );
  mux2_1 U19361 ( .ip1(\ANSWER/mem[2][3][11] ), .ip2(\ANSWER/mem[3][3][11] ), 
        .s(n18465), .op(n18410) );
  mux2_1 U19362 ( .ip1(n18411), .ip2(n18410), .s(n18435), .op(n18415) );
  mux2_1 U19363 ( .ip1(\ANSWER/mem[4][3][11] ), .ip2(\ANSWER/mem[5][3][11] ), 
        .s(n18465), .op(n18413) );
  mux2_1 U19364 ( .ip1(\ANSWER/mem[6][3][11] ), .ip2(\ANSWER/mem[7][3][11] ), 
        .s(n18465), .op(n18412) );
  mux2_1 U19365 ( .ip1(n18413), .ip2(n18412), .s(n18435), .op(n18414) );
  mux2_1 U19366 ( .ip1(n18415), .ip2(n18414), .s(n18906), .op(n18417) );
  mux2_1 U19367 ( .ip1(\ANSWER/mem[8][3][11] ), .ip2(\ANSWER/mem[9][3][11] ), 
        .s(n18465), .op(n18416) );
  mux2_1 U19368 ( .ip1(n18417), .ip2(n18416), .s(n18466), .op(n18418) );
  nand2_1 U19369 ( .ip1(n18854), .ip2(n18418), .op(n18429) );
  mux2_1 U19370 ( .ip1(\ANSWER/mem[0][7][11] ), .ip2(\ANSWER/mem[1][7][11] ), 
        .s(n18458), .op(n18420) );
  mux2_1 U19371 ( .ip1(\ANSWER/mem[2][7][11] ), .ip2(\ANSWER/mem[3][7][11] ), 
        .s(n18458), .op(n18419) );
  mux2_1 U19372 ( .ip1(n18420), .ip2(n18419), .s(n17688), .op(n18424) );
  mux2_1 U19373 ( .ip1(\ANSWER/mem[4][7][11] ), .ip2(\ANSWER/mem[5][7][11] ), 
        .s(n18458), .op(n18422) );
  mux2_1 U19374 ( .ip1(\ANSWER/mem[6][7][11] ), .ip2(\ANSWER/mem[7][7][11] ), 
        .s(n18458), .op(n18421) );
  mux2_1 U19375 ( .ip1(n18422), .ip2(n18421), .s(n4456), .op(n18423) );
  mux2_1 U19376 ( .ip1(n18424), .ip2(n18423), .s(n18906), .op(n18426) );
  mux2_1 U19377 ( .ip1(\ANSWER/mem[8][7][11] ), .ip2(\ANSWER/mem[9][7][11] ), 
        .s(n18465), .op(n18425) );
  mux2_1 U19378 ( .ip1(n18426), .ip2(n18425), .s(n18466), .op(n18427) );
  nand2_1 U19379 ( .ip1(n18865), .ip2(n18427), .op(n18428) );
  nand4_1 U19380 ( .ip1(n18431), .ip2(n18430), .ip3(n18429), .ip4(n18428), 
        .op(n18432) );
  not_ab_or_c_or_d U19381 ( .ip1(n18884), .ip2(n18434), .ip3(n18433), .ip4(
        n18432), .op(n18446) );
  mux2_1 U19382 ( .ip1(\ANSWER/mem[0][6][11] ), .ip2(\ANSWER/mem[1][6][11] ), 
        .s(n18458), .op(n18437) );
  mux2_1 U19383 ( .ip1(\ANSWER/mem[2][6][11] ), .ip2(\ANSWER/mem[3][6][11] ), 
        .s(n18458), .op(n18436) );
  mux2_1 U19384 ( .ip1(n18437), .ip2(n18436), .s(n18435), .op(n18441) );
  mux2_1 U19385 ( .ip1(\ANSWER/mem[4][6][11] ), .ip2(\ANSWER/mem[5][6][11] ), 
        .s(n18458), .op(n18439) );
  mux2_1 U19386 ( .ip1(\ANSWER/mem[6][6][11] ), .ip2(\ANSWER/mem[7][6][11] ), 
        .s(n18458), .op(n18438) );
  mux2_1 U19387 ( .ip1(n18439), .ip2(n18438), .s(n18435), .op(n18440) );
  mux2_1 U19388 ( .ip1(n18441), .ip2(n18440), .s(n18906), .op(n18443) );
  mux2_1 U19389 ( .ip1(\ANSWER/mem[8][6][11] ), .ip2(\ANSWER/mem[9][6][11] ), 
        .s(n18458), .op(n18442) );
  mux2_1 U19390 ( .ip1(n18443), .ip2(n18442), .s(n18466), .op(n18444) );
  nand2_1 U19391 ( .ip1(n18821), .ip2(n18444), .op(n18445) );
  nand3_1 U19392 ( .ip1(n18447), .ip2(n18446), .ip3(n18445), .op(n18448) );
  nand2_1 U19393 ( .ip1(n18448), .ip2(n18888), .op(n18472) );
  mux2_1 U19394 ( .ip1(\ANSWER/mem[0][9][11] ), .ip2(\ANSWER/mem[1][9][11] ), 
        .s(n18465), .op(n18450) );
  mux2_1 U19395 ( .ip1(\ANSWER/mem[2][9][11] ), .ip2(\ANSWER/mem[3][9][11] ), 
        .s(n18458), .op(n18449) );
  mux2_1 U19396 ( .ip1(n18450), .ip2(n18449), .s(n4456), .op(n18454) );
  mux2_1 U19397 ( .ip1(\ANSWER/mem[4][9][11] ), .ip2(\ANSWER/mem[5][9][11] ), 
        .s(n18465), .op(n18452) );
  mux2_1 U19398 ( .ip1(\ANSWER/mem[6][9][11] ), .ip2(\ANSWER/mem[7][9][11] ), 
        .s(n18465), .op(n18451) );
  mux2_1 U19399 ( .ip1(n18452), .ip2(n18451), .s(n17605), .op(n18453) );
  mux2_1 U19400 ( .ip1(n18454), .ip2(n18453), .s(n18906), .op(n18456) );
  mux2_1 U19401 ( .ip1(\ANSWER/mem[8][9][11] ), .ip2(\ANSWER/mem[9][9][11] ), 
        .s(n18465), .op(n18455) );
  mux2_1 U19402 ( .ip1(n18456), .ip2(n18455), .s(n18466), .op(n18457) );
  nand2_1 U19403 ( .ip1(n18899), .ip2(n18457), .op(n18471) );
  mux2_1 U19404 ( .ip1(\ANSWER/mem[0][8][11] ), .ip2(\ANSWER/mem[1][8][11] ), 
        .s(n18458), .op(n18460) );
  mux2_1 U19405 ( .ip1(\ANSWER/mem[2][8][11] ), .ip2(\ANSWER/mem[3][8][11] ), 
        .s(n18458), .op(n18459) );
  mux2_1 U19406 ( .ip1(n18460), .ip2(n18459), .s(n17581), .op(n18464) );
  mux2_1 U19407 ( .ip1(\ANSWER/mem[4][8][11] ), .ip2(\ANSWER/mem[5][8][11] ), 
        .s(n18465), .op(n18462) );
  mux2_1 U19408 ( .ip1(\ANSWER/mem[6][8][11] ), .ip2(\ANSWER/mem[7][8][11] ), 
        .s(n18465), .op(n18461) );
  mux2_1 U19409 ( .ip1(n18462), .ip2(n18461), .s(n17794), .op(n18463) );
  mux2_1 U19410 ( .ip1(n18464), .ip2(n18463), .s(n18906), .op(n18468) );
  mux2_1 U19411 ( .ip1(\ANSWER/mem[8][8][11] ), .ip2(\ANSWER/mem[9][8][11] ), 
        .s(n18465), .op(n18467) );
  mux2_1 U19412 ( .ip1(n18468), .ip2(n18467), .s(n18466), .op(n18469) );
  nand2_1 U19413 ( .ip1(n18914), .ip2(n18469), .op(n18470) );
  nand3_1 U19414 ( .ip1(n18472), .ip2(n18471), .ip3(n18470), .op(\ANSWER/N476 ) );
  inv_1 U19415 ( .ip(n4362), .op(n18572) );
  mux2_1 U19416 ( .ip1(\ANSWER/mem[0][3][12] ), .ip2(\ANSWER/mem[1][3][12] ), 
        .s(n18572), .op(n18474) );
  mux2_1 U19417 ( .ip1(\ANSWER/mem[2][3][12] ), .ip2(\ANSWER/mem[3][3][12] ), 
        .s(n18572), .op(n18473) );
  inv_1 U19418 ( .ip(n4366), .op(n18544) );
  mux2_1 U19419 ( .ip1(n18474), .ip2(n18473), .s(n18544), .op(n18478) );
  mux2_1 U19420 ( .ip1(\ANSWER/mem[4][3][12] ), .ip2(\ANSWER/mem[5][3][12] ), 
        .s(n18572), .op(n18476) );
  mux2_1 U19421 ( .ip1(\ANSWER/mem[6][3][12] ), .ip2(\ANSWER/mem[7][3][12] ), 
        .s(n18572), .op(n18475) );
  mux2_1 U19422 ( .ip1(n18476), .ip2(n18475), .s(n18544), .op(n18477) );
  mux2_1 U19423 ( .ip1(n18478), .ip2(n18477), .s(n18826), .op(n18480) );
  mux2_1 U19424 ( .ip1(\ANSWER/mem[8][3][12] ), .ip2(\ANSWER/mem[9][3][12] ), 
        .s(n18572), .op(n18479) );
  mux2_1 U19425 ( .ip1(n18480), .ip2(n18479), .s(n18679), .op(n18481) );
  nand2_1 U19426 ( .ip1(n18854), .ip2(n18481), .op(n18554) );
  mux2_1 U19427 ( .ip1(\ANSWER/mem[0][0][12] ), .ip2(\ANSWER/mem[1][0][12] ), 
        .s(n17536), .op(n18483) );
  mux2_1 U19428 ( .ip1(\ANSWER/mem[2][0][12] ), .ip2(\ANSWER/mem[3][0][12] ), 
        .s(n17536), .op(n18482) );
  mux2_1 U19429 ( .ip1(n18483), .ip2(n18482), .s(n18544), .op(n18487) );
  mux2_1 U19430 ( .ip1(\ANSWER/mem[4][0][12] ), .ip2(\ANSWER/mem[5][0][12] ), 
        .s(n17533), .op(n18485) );
  mux2_1 U19431 ( .ip1(\ANSWER/mem[6][0][12] ), .ip2(\ANSWER/mem[7][0][12] ), 
        .s(n17533), .op(n18484) );
  mux2_1 U19432 ( .ip1(n18485), .ip2(n18484), .s(n18544), .op(n18486) );
  mux2_1 U19433 ( .ip1(n18487), .ip2(n18486), .s(n18826), .op(n18489) );
  mux2_1 U19434 ( .ip1(\ANSWER/mem[8][0][12] ), .ip2(\ANSWER/mem[9][0][12] ), 
        .s(n18900), .op(n18488) );
  mux2_1 U19435 ( .ip1(n18489), .ip2(n18488), .s(n18679), .op(n18541) );
  buf_1 U19436 ( .ip(n18572), .op(n18565) );
  mux2_1 U19437 ( .ip1(\ANSWER/mem[0][6][12] ), .ip2(\ANSWER/mem[1][6][12] ), 
        .s(n18565), .op(n18491) );
  mux2_1 U19438 ( .ip1(\ANSWER/mem[2][6][12] ), .ip2(\ANSWER/mem[3][6][12] ), 
        .s(n18565), .op(n18490) );
  mux2_1 U19439 ( .ip1(n18491), .ip2(n18490), .s(n18544), .op(n18495) );
  mux2_1 U19440 ( .ip1(\ANSWER/mem[4][6][12] ), .ip2(\ANSWER/mem[5][6][12] ), 
        .s(n18565), .op(n18493) );
  mux2_1 U19441 ( .ip1(\ANSWER/mem[6][6][12] ), .ip2(\ANSWER/mem[7][6][12] ), 
        .s(n18565), .op(n18492) );
  mux2_1 U19442 ( .ip1(n18493), .ip2(n18492), .s(n17605), .op(n18494) );
  mux2_1 U19443 ( .ip1(n18495), .ip2(n18494), .s(n18906), .op(n18497) );
  mux2_1 U19444 ( .ip1(\ANSWER/mem[8][6][12] ), .ip2(\ANSWER/mem[9][6][12] ), 
        .s(n18565), .op(n18496) );
  mux2_1 U19445 ( .ip1(n18497), .ip2(n18496), .s(n18679), .op(n18498) );
  and2_1 U19446 ( .ip1(n18821), .ip2(n18498), .op(n18540) );
  mux2_1 U19447 ( .ip1(\ANSWER/mem[0][1][12] ), .ip2(\ANSWER/mem[1][1][12] ), 
        .s(n17344), .op(n18500) );
  mux2_1 U19448 ( .ip1(\ANSWER/mem[2][1][12] ), .ip2(\ANSWER/mem[3][1][12] ), 
        .s(n17533), .op(n18499) );
  mux2_1 U19449 ( .ip1(n18500), .ip2(n18499), .s(n18544), .op(n18504) );
  mux2_1 U19450 ( .ip1(\ANSWER/mem[4][1][12] ), .ip2(\ANSWER/mem[5][1][12] ), 
        .s(n17884), .op(n18502) );
  mux2_1 U19451 ( .ip1(\ANSWER/mem[6][1][12] ), .ip2(\ANSWER/mem[7][1][12] ), 
        .s(n17536), .op(n18501) );
  mux2_1 U19452 ( .ip1(n18502), .ip2(n18501), .s(n18544), .op(n18503) );
  mux2_1 U19453 ( .ip1(n18504), .ip2(n18503), .s(n18826), .op(n18506) );
  mux2_1 U19454 ( .ip1(\ANSWER/mem[8][1][12] ), .ip2(\ANSWER/mem[9][1][12] ), 
        .s(n17536), .op(n18505) );
  mux2_1 U19455 ( .ip1(n18506), .ip2(n18505), .s(n18679), .op(n18507) );
  nand2_1 U19456 ( .ip1(n18872), .ip2(n18507), .op(n18538) );
  mux2_1 U19457 ( .ip1(\ANSWER/mem[0][2][12] ), .ip2(\ANSWER/mem[1][2][12] ), 
        .s(n18351), .op(n18509) );
  mux2_1 U19458 ( .ip1(\ANSWER/mem[2][2][12] ), .ip2(\ANSWER/mem[3][2][12] ), 
        .s(n18616), .op(n18508) );
  mux2_1 U19459 ( .ip1(n18509), .ip2(n18508), .s(n18544), .op(n18513) );
  mux2_1 U19460 ( .ip1(\ANSWER/mem[4][2][12] ), .ip2(\ANSWER/mem[5][2][12] ), 
        .s(n18741), .op(n18511) );
  mux2_1 U19461 ( .ip1(\ANSWER/mem[6][2][12] ), .ip2(\ANSWER/mem[7][2][12] ), 
        .s(n18572), .op(n18510) );
  mux2_1 U19462 ( .ip1(n18511), .ip2(n18510), .s(n18544), .op(n18512) );
  mux2_1 U19463 ( .ip1(n18513), .ip2(n18512), .s(n18906), .op(n18515) );
  mux2_1 U19464 ( .ip1(\ANSWER/mem[8][2][12] ), .ip2(\ANSWER/mem[9][2][12] ), 
        .s(n18572), .op(n18514) );
  mux2_1 U19465 ( .ip1(n18515), .ip2(n18514), .s(n18679), .op(n18516) );
  nand2_1 U19466 ( .ip1(n18884), .ip2(n18516), .op(n18537) );
  mux2_1 U19467 ( .ip1(\ANSWER/mem[0][4][12] ), .ip2(\ANSWER/mem[1][4][12] ), 
        .s(n18572), .op(n18518) );
  mux2_1 U19468 ( .ip1(\ANSWER/mem[2][4][12] ), .ip2(\ANSWER/mem[3][4][12] ), 
        .s(n18572), .op(n18517) );
  mux2_1 U19469 ( .ip1(n18518), .ip2(n18517), .s(n18544), .op(n18522) );
  mux2_1 U19470 ( .ip1(\ANSWER/mem[4][4][12] ), .ip2(\ANSWER/mem[5][4][12] ), 
        .s(n18572), .op(n18520) );
  mux2_1 U19471 ( .ip1(\ANSWER/mem[6][4][12] ), .ip2(\ANSWER/mem[7][4][12] ), 
        .s(n18572), .op(n18519) );
  mux2_1 U19472 ( .ip1(n18520), .ip2(n18519), .s(n18544), .op(n18521) );
  mux2_1 U19473 ( .ip1(n18522), .ip2(n18521), .s(n18826), .op(n18524) );
  mux2_1 U19474 ( .ip1(\ANSWER/mem[8][4][12] ), .ip2(\ANSWER/mem[9][4][12] ), 
        .s(n18572), .op(n18523) );
  mux2_1 U19475 ( .ip1(n18524), .ip2(n18523), .s(n18679), .op(n18525) );
  nand2_1 U19476 ( .ip1(n18843), .ip2(n18525), .op(n18536) );
  mux2_1 U19477 ( .ip1(\ANSWER/mem[0][7][12] ), .ip2(\ANSWER/mem[1][7][12] ), 
        .s(n18565), .op(n18527) );
  mux2_1 U19478 ( .ip1(\ANSWER/mem[2][7][12] ), .ip2(\ANSWER/mem[3][7][12] ), 
        .s(n18565), .op(n18526) );
  mux2_1 U19479 ( .ip1(n18527), .ip2(n18526), .s(n17366), .op(n18531) );
  mux2_1 U19480 ( .ip1(\ANSWER/mem[4][7][12] ), .ip2(\ANSWER/mem[5][7][12] ), 
        .s(n18565), .op(n18529) );
  mux2_1 U19481 ( .ip1(\ANSWER/mem[6][7][12] ), .ip2(\ANSWER/mem[7][7][12] ), 
        .s(n18565), .op(n18528) );
  mux2_1 U19482 ( .ip1(n18529), .ip2(n18528), .s(n17366), .op(n18530) );
  mux2_1 U19483 ( .ip1(n18531), .ip2(n18530), .s(n18906), .op(n18533) );
  mux2_1 U19484 ( .ip1(\ANSWER/mem[8][7][12] ), .ip2(\ANSWER/mem[9][7][12] ), 
        .s(n18572), .op(n18532) );
  mux2_1 U19485 ( .ip1(n18533), .ip2(n18532), .s(n18679), .op(n18534) );
  nand2_1 U19486 ( .ip1(n18865), .ip2(n18534), .op(n18535) );
  nand4_1 U19487 ( .ip1(n18538), .ip2(n18537), .ip3(n18536), .ip4(n18535), 
        .op(n18539) );
  not_ab_or_c_or_d U19488 ( .ip1(n18800), .ip2(n18541), .ip3(n18540), .ip4(
        n18539), .op(n18553) );
  mux2_1 U19489 ( .ip1(\ANSWER/mem[0][5][12] ), .ip2(\ANSWER/mem[1][5][12] ), 
        .s(n18572), .op(n18543) );
  mux2_1 U19490 ( .ip1(\ANSWER/mem[2][5][12] ), .ip2(\ANSWER/mem[3][5][12] ), 
        .s(n18565), .op(n18542) );
  mux2_1 U19491 ( .ip1(n18543), .ip2(n18542), .s(n18544), .op(n18548) );
  mux2_1 U19492 ( .ip1(\ANSWER/mem[4][5][12] ), .ip2(\ANSWER/mem[5][5][12] ), 
        .s(n18565), .op(n18546) );
  mux2_1 U19493 ( .ip1(\ANSWER/mem[6][5][12] ), .ip2(\ANSWER/mem[7][5][12] ), 
        .s(n18565), .op(n18545) );
  mux2_1 U19494 ( .ip1(n18546), .ip2(n18545), .s(n18544), .op(n18547) );
  mux2_1 U19495 ( .ip1(n18548), .ip2(n18547), .s(n18906), .op(n18550) );
  mux2_1 U19496 ( .ip1(\ANSWER/mem[8][5][12] ), .ip2(\ANSWER/mem[9][5][12] ), 
        .s(n18565), .op(n18549) );
  mux2_1 U19497 ( .ip1(n18550), .ip2(n18549), .s(n18679), .op(n18551) );
  nand2_1 U19498 ( .ip1(n18832), .ip2(n18551), .op(n18552) );
  nand3_1 U19499 ( .ip1(n18554), .ip2(n18553), .ip3(n18552), .op(n18555) );
  nand2_1 U19500 ( .ip1(n18555), .ip2(n18888), .op(n18578) );
  mux2_1 U19501 ( .ip1(\ANSWER/mem[0][9][12] ), .ip2(\ANSWER/mem[1][9][12] ), 
        .s(n18572), .op(n18557) );
  mux2_1 U19502 ( .ip1(\ANSWER/mem[2][9][12] ), .ip2(\ANSWER/mem[3][9][12] ), 
        .s(n18565), .op(n18556) );
  mux2_1 U19503 ( .ip1(n18557), .ip2(n18556), .s(n18330), .op(n18561) );
  mux2_1 U19504 ( .ip1(\ANSWER/mem[4][9][12] ), .ip2(\ANSWER/mem[5][9][12] ), 
        .s(n18572), .op(n18559) );
  mux2_1 U19505 ( .ip1(\ANSWER/mem[6][9][12] ), .ip2(\ANSWER/mem[7][9][12] ), 
        .s(n18572), .op(n18558) );
  mux2_1 U19506 ( .ip1(n18559), .ip2(n18558), .s(n18435), .op(n18560) );
  mux2_1 U19507 ( .ip1(n18561), .ip2(n18560), .s(n18906), .op(n18563) );
  mux2_1 U19508 ( .ip1(\ANSWER/mem[8][9][12] ), .ip2(\ANSWER/mem[9][9][12] ), 
        .s(n18572), .op(n18562) );
  mux2_1 U19509 ( .ip1(n18563), .ip2(n18562), .s(n18679), .op(n18564) );
  nand2_1 U19510 ( .ip1(n18899), .ip2(n18564), .op(n18577) );
  mux2_1 U19511 ( .ip1(\ANSWER/mem[0][8][12] ), .ip2(\ANSWER/mem[1][8][12] ), 
        .s(n18565), .op(n18567) );
  mux2_1 U19512 ( .ip1(\ANSWER/mem[2][8][12] ), .ip2(\ANSWER/mem[3][8][12] ), 
        .s(n18565), .op(n18566) );
  mux2_1 U19513 ( .ip1(n18567), .ip2(n18566), .s(n18354), .op(n18571) );
  mux2_1 U19514 ( .ip1(\ANSWER/mem[4][8][12] ), .ip2(\ANSWER/mem[5][8][12] ), 
        .s(n18572), .op(n18569) );
  mux2_1 U19515 ( .ip1(\ANSWER/mem[6][8][12] ), .ip2(\ANSWER/mem[7][8][12] ), 
        .s(n18572), .op(n18568) );
  mux2_1 U19516 ( .ip1(n18569), .ip2(n18568), .s(n18112), .op(n18570) );
  mux2_1 U19517 ( .ip1(n18571), .ip2(n18570), .s(n18826), .op(n18574) );
  mux2_1 U19518 ( .ip1(\ANSWER/mem[8][8][12] ), .ip2(\ANSWER/mem[9][8][12] ), 
        .s(n18572), .op(n18573) );
  mux2_1 U19519 ( .ip1(n18574), .ip2(n18573), .s(n18679), .op(n18575) );
  nand2_1 U19520 ( .ip1(n18914), .ip2(n18575), .op(n18576) );
  nand3_1 U19521 ( .ip1(n18578), .ip2(n18577), .ip3(n18576), .op(\ANSWER/N475 ) );
  inv_1 U19522 ( .ip(n4362), .op(n18616) );
  mux2_1 U19523 ( .ip1(\ANSWER/mem[0][1][13] ), .ip2(\ANSWER/mem[1][1][13] ), 
        .s(n18616), .op(n18580) );
  mux2_1 U19524 ( .ip1(\ANSWER/mem[2][1][13] ), .ip2(\ANSWER/mem[3][1][13] ), 
        .s(n18616), .op(n18579) );
  mux2_1 U19525 ( .ip1(n18580), .ip2(n18579), .s(n18544), .op(n18584) );
  mux2_1 U19526 ( .ip1(\ANSWER/mem[4][1][13] ), .ip2(\ANSWER/mem[5][1][13] ), 
        .s(n18616), .op(n18582) );
  mux2_1 U19527 ( .ip1(\ANSWER/mem[6][1][13] ), .ip2(\ANSWER/mem[7][1][13] ), 
        .s(n18616), .op(n18581) );
  mux2_1 U19528 ( .ip1(n18582), .ip2(n18581), .s(n18138), .op(n18583) );
  mux2_1 U19529 ( .ip1(n18584), .ip2(n18583), .s(n18859), .op(n18586) );
  mux2_1 U19530 ( .ip1(\ANSWER/mem[8][1][13] ), .ip2(\ANSWER/mem[9][1][13] ), 
        .s(n18616), .op(n18585) );
  mux2_1 U19531 ( .ip1(n18586), .ip2(n18585), .s(n18679), .op(n18587) );
  nand2_1 U19532 ( .ip1(n18872), .ip2(n18587), .op(n18660) );
  inv_1 U19533 ( .ip(n4362), .op(n18678) );
  mux2_1 U19534 ( .ip1(\ANSWER/mem[0][4][13] ), .ip2(\ANSWER/mem[1][4][13] ), 
        .s(n18678), .op(n18589) );
  mux2_1 U19535 ( .ip1(\ANSWER/mem[2][4][13] ), .ip2(\ANSWER/mem[3][4][13] ), 
        .s(n18678), .op(n18588) );
  mux2_1 U19536 ( .ip1(n18589), .ip2(n18588), .s(n15636), .op(n18593) );
  mux2_1 U19537 ( .ip1(\ANSWER/mem[4][4][13] ), .ip2(\ANSWER/mem[5][4][13] ), 
        .s(n18678), .op(n18591) );
  mux2_1 U19538 ( .ip1(\ANSWER/mem[6][4][13] ), .ip2(\ANSWER/mem[7][4][13] ), 
        .s(n18678), .op(n18590) );
  mux2_1 U19539 ( .ip1(n18591), .ip2(n18590), .s(n18112), .op(n18592) );
  mux2_1 U19540 ( .ip1(n18593), .ip2(n18592), .s(n18815), .op(n18595) );
  mux2_1 U19541 ( .ip1(\ANSWER/mem[8][4][13] ), .ip2(\ANSWER/mem[9][4][13] ), 
        .s(n18678), .op(n18594) );
  mux2_1 U19542 ( .ip1(n18595), .ip2(n18594), .s(n18679), .op(n18648) );
  buf_1 U19543 ( .ip(n18678), .op(n18671) );
  mux2_1 U19544 ( .ip1(\ANSWER/mem[0][6][13] ), .ip2(\ANSWER/mem[1][6][13] ), 
        .s(n18671), .op(n18597) );
  mux2_1 U19545 ( .ip1(\ANSWER/mem[2][6][13] ), .ip2(\ANSWER/mem[3][6][13] ), 
        .s(n18671), .op(n18596) );
  mux2_1 U19546 ( .ip1(n18597), .ip2(n18596), .s(n4456), .op(n18601) );
  mux2_1 U19547 ( .ip1(\ANSWER/mem[4][6][13] ), .ip2(\ANSWER/mem[5][6][13] ), 
        .s(n18671), .op(n18599) );
  mux2_1 U19548 ( .ip1(\ANSWER/mem[6][6][13] ), .ip2(\ANSWER/mem[7][6][13] ), 
        .s(n18671), .op(n18598) );
  mux2_1 U19549 ( .ip1(n18599), .ip2(n18598), .s(n4456), .op(n18600) );
  mux2_1 U19550 ( .ip1(n18601), .ip2(n18600), .s(n18806), .op(n18603) );
  mux2_1 U19551 ( .ip1(\ANSWER/mem[8][6][13] ), .ip2(\ANSWER/mem[9][6][13] ), 
        .s(n18671), .op(n18602) );
  mux2_1 U19552 ( .ip1(n18603), .ip2(n18602), .s(n18679), .op(n18604) );
  and2_1 U19553 ( .ip1(n18821), .ip2(n18604), .op(n18647) );
  mux2_1 U19554 ( .ip1(\ANSWER/mem[0][0][13] ), .ip2(\ANSWER/mem[1][0][13] ), 
        .s(n18616), .op(n18606) );
  mux2_1 U19555 ( .ip1(\ANSWER/mem[2][0][13] ), .ip2(\ANSWER/mem[3][0][13] ), 
        .s(n18616), .op(n18605) );
  mux2_1 U19556 ( .ip1(n18606), .ip2(n18605), .s(n18544), .op(n18610) );
  mux2_1 U19557 ( .ip1(\ANSWER/mem[4][0][13] ), .ip2(\ANSWER/mem[5][0][13] ), 
        .s(n18616), .op(n18608) );
  mux2_1 U19558 ( .ip1(\ANSWER/mem[6][0][13] ), .ip2(\ANSWER/mem[7][0][13] ), 
        .s(n18616), .op(n18607) );
  mux2_1 U19559 ( .ip1(n18608), .ip2(n18607), .s(n18138), .op(n18609) );
  mux2_1 U19560 ( .ip1(n18610), .ip2(n18609), .s(n18815), .op(n18612) );
  mux2_1 U19561 ( .ip1(\ANSWER/mem[8][0][13] ), .ip2(\ANSWER/mem[9][0][13] ), 
        .s(n18616), .op(n18611) );
  mux2_1 U19562 ( .ip1(n18612), .ip2(n18611), .s(n18679), .op(n18613) );
  nand2_1 U19563 ( .ip1(n18800), .ip2(n18613), .op(n18645) );
  mux2_1 U19564 ( .ip1(\ANSWER/mem[0][2][13] ), .ip2(\ANSWER/mem[1][2][13] ), 
        .s(n18616), .op(n18615) );
  mux2_1 U19565 ( .ip1(\ANSWER/mem[2][2][13] ), .ip2(\ANSWER/mem[3][2][13] ), 
        .s(n18616), .op(n18614) );
  mux2_1 U19566 ( .ip1(n18615), .ip2(n18614), .s(n17366), .op(n18620) );
  mux2_1 U19567 ( .ip1(\ANSWER/mem[4][2][13] ), .ip2(\ANSWER/mem[5][2][13] ), 
        .s(n18616), .op(n18618) );
  mux2_1 U19568 ( .ip1(\ANSWER/mem[6][2][13] ), .ip2(\ANSWER/mem[7][2][13] ), 
        .s(n18678), .op(n18617) );
  mux2_1 U19569 ( .ip1(n18618), .ip2(n18617), .s(n18354), .op(n18619) );
  mux2_1 U19570 ( .ip1(n18620), .ip2(n18619), .s(n18806), .op(n18622) );
  mux2_1 U19571 ( .ip1(\ANSWER/mem[8][2][13] ), .ip2(\ANSWER/mem[9][2][13] ), 
        .s(n18678), .op(n18621) );
  mux2_1 U19572 ( .ip1(n18622), .ip2(n18621), .s(n18679), .op(n18623) );
  nand2_1 U19573 ( .ip1(n18884), .ip2(n18623), .op(n18644) );
  mux2_1 U19574 ( .ip1(\ANSWER/mem[0][5][13] ), .ip2(\ANSWER/mem[1][5][13] ), 
        .s(n18678), .op(n18625) );
  mux2_1 U19575 ( .ip1(\ANSWER/mem[2][5][13] ), .ip2(\ANSWER/mem[3][5][13] ), 
        .s(n18671), .op(n18624) );
  mux2_1 U19576 ( .ip1(n18625), .ip2(n18624), .s(n18544), .op(n18629) );
  mux2_1 U19577 ( .ip1(\ANSWER/mem[4][5][13] ), .ip2(\ANSWER/mem[5][5][13] ), 
        .s(n18671), .op(n18627) );
  mux2_1 U19578 ( .ip1(\ANSWER/mem[6][5][13] ), .ip2(\ANSWER/mem[7][5][13] ), 
        .s(n18671), .op(n18626) );
  mux2_1 U19579 ( .ip1(n18627), .ip2(n18626), .s(n18544), .op(n18628) );
  mux2_1 U19580 ( .ip1(n18629), .ip2(n18628), .s(n18806), .op(n18631) );
  mux2_1 U19581 ( .ip1(\ANSWER/mem[8][5][13] ), .ip2(\ANSWER/mem[9][5][13] ), 
        .s(n18671), .op(n18630) );
  mux2_1 U19582 ( .ip1(n18631), .ip2(n18630), .s(n18679), .op(n18632) );
  nand2_1 U19583 ( .ip1(n18832), .ip2(n18632), .op(n18643) );
  mux2_1 U19584 ( .ip1(\ANSWER/mem[0][7][13] ), .ip2(\ANSWER/mem[1][7][13] ), 
        .s(n18671), .op(n18634) );
  mux2_1 U19585 ( .ip1(\ANSWER/mem[2][7][13] ), .ip2(\ANSWER/mem[3][7][13] ), 
        .s(n18671), .op(n18633) );
  mux2_1 U19586 ( .ip1(n18634), .ip2(n18633), .s(n17581), .op(n18638) );
  mux2_1 U19587 ( .ip1(\ANSWER/mem[4][7][13] ), .ip2(\ANSWER/mem[5][7][13] ), 
        .s(n18671), .op(n18636) );
  mux2_1 U19588 ( .ip1(\ANSWER/mem[6][7][13] ), .ip2(\ANSWER/mem[7][7][13] ), 
        .s(n18671), .op(n18635) );
  mux2_1 U19589 ( .ip1(n18636), .ip2(n18635), .s(n18435), .op(n18637) );
  mux2_1 U19590 ( .ip1(n18638), .ip2(n18637), .s(n18815), .op(n18640) );
  mux2_1 U19591 ( .ip1(\ANSWER/mem[8][7][13] ), .ip2(\ANSWER/mem[9][7][13] ), 
        .s(n18678), .op(n18639) );
  mux2_1 U19592 ( .ip1(n18640), .ip2(n18639), .s(n18679), .op(n18641) );
  nand2_1 U19593 ( .ip1(n18865), .ip2(n18641), .op(n18642) );
  nand4_1 U19594 ( .ip1(n18645), .ip2(n18644), .ip3(n18643), .ip4(n18642), 
        .op(n18646) );
  not_ab_or_c_or_d U19595 ( .ip1(n18843), .ip2(n18648), .ip3(n18647), .ip4(
        n18646), .op(n18659) );
  mux2_1 U19596 ( .ip1(\ANSWER/mem[0][3][13] ), .ip2(\ANSWER/mem[1][3][13] ), 
        .s(n18678), .op(n18650) );
  mux2_1 U19597 ( .ip1(\ANSWER/mem[2][3][13] ), .ip2(\ANSWER/mem[3][3][13] ), 
        .s(n18678), .op(n18649) );
  mux2_1 U19598 ( .ip1(n18650), .ip2(n18649), .s(n17605), .op(n18654) );
  mux2_1 U19599 ( .ip1(\ANSWER/mem[4][3][13] ), .ip2(\ANSWER/mem[5][3][13] ), 
        .s(n18678), .op(n18652) );
  mux2_1 U19600 ( .ip1(\ANSWER/mem[6][3][13] ), .ip2(\ANSWER/mem[7][3][13] ), 
        .s(n18678), .op(n18651) );
  mux2_1 U19601 ( .ip1(n18652), .ip2(n18651), .s(n17688), .op(n18653) );
  mux2_1 U19602 ( .ip1(n18654), .ip2(n18653), .s(n18815), .op(n18656) );
  mux2_1 U19603 ( .ip1(\ANSWER/mem[8][3][13] ), .ip2(\ANSWER/mem[9][3][13] ), 
        .s(n18678), .op(n18655) );
  mux2_1 U19604 ( .ip1(n18656), .ip2(n18655), .s(n18679), .op(n18657) );
  nand2_1 U19605 ( .ip1(n18854), .ip2(n18657), .op(n18658) );
  nand3_1 U19606 ( .ip1(n18660), .ip2(n18659), .ip3(n18658), .op(n18661) );
  nand2_1 U19607 ( .ip1(n18661), .ip2(n18888), .op(n18685) );
  mux2_1 U19608 ( .ip1(\ANSWER/mem[0][8][13] ), .ip2(\ANSWER/mem[1][8][13] ), 
        .s(n18678), .op(n18663) );
  mux2_1 U19609 ( .ip1(\ANSWER/mem[2][8][13] ), .ip2(\ANSWER/mem[3][8][13] ), 
        .s(n18671), .op(n18662) );
  mux2_1 U19610 ( .ip1(n18663), .ip2(n18662), .s(n18901), .op(n18667) );
  mux2_1 U19611 ( .ip1(\ANSWER/mem[4][8][13] ), .ip2(\ANSWER/mem[5][8][13] ), 
        .s(n18678), .op(n18665) );
  mux2_1 U19612 ( .ip1(\ANSWER/mem[6][8][13] ), .ip2(\ANSWER/mem[7][8][13] ), 
        .s(n18678), .op(n18664) );
  mux2_1 U19613 ( .ip1(n18665), .ip2(n18664), .s(n18901), .op(n18666) );
  mux2_1 U19614 ( .ip1(n18667), .ip2(n18666), .s(n18806), .op(n18669) );
  mux2_1 U19615 ( .ip1(\ANSWER/mem[8][8][13] ), .ip2(\ANSWER/mem[9][8][13] ), 
        .s(n18678), .op(n18668) );
  mux2_1 U19616 ( .ip1(n18669), .ip2(n18668), .s(n18679), .op(n18670) );
  nand2_1 U19617 ( .ip1(n18914), .ip2(n18670), .op(n18684) );
  mux2_1 U19618 ( .ip1(\ANSWER/mem[0][9][13] ), .ip2(\ANSWER/mem[1][9][13] ), 
        .s(n18671), .op(n18673) );
  mux2_1 U19619 ( .ip1(\ANSWER/mem[2][9][13] ), .ip2(\ANSWER/mem[3][9][13] ), 
        .s(n18671), .op(n18672) );
  mux2_1 U19620 ( .ip1(n18673), .ip2(n18672), .s(n18901), .op(n18677) );
  mux2_1 U19621 ( .ip1(\ANSWER/mem[4][9][13] ), .ip2(\ANSWER/mem[5][9][13] ), 
        .s(n18678), .op(n18675) );
  mux2_1 U19622 ( .ip1(\ANSWER/mem[6][9][13] ), .ip2(\ANSWER/mem[7][9][13] ), 
        .s(n18678), .op(n18674) );
  mux2_1 U19623 ( .ip1(n18675), .ip2(n18674), .s(n18901), .op(n18676) );
  mux2_1 U19624 ( .ip1(n18677), .ip2(n18676), .s(n18859), .op(n18681) );
  mux2_1 U19625 ( .ip1(\ANSWER/mem[8][9][13] ), .ip2(\ANSWER/mem[9][9][13] ), 
        .s(n18678), .op(n18680) );
  mux2_1 U19626 ( .ip1(n18681), .ip2(n18680), .s(n18679), .op(n18682) );
  nand2_1 U19627 ( .ip1(n18899), .ip2(n18682), .op(n18683) );
  nand3_1 U19628 ( .ip1(n18685), .ip2(n18684), .ip3(n18683), .op(\ANSWER/N474 ) );
  inv_1 U19629 ( .ip(n4362), .op(n18785) );
  mux2_1 U19630 ( .ip1(\ANSWER/mem[0][5][14] ), .ip2(\ANSWER/mem[1][5][14] ), 
        .s(n18785), .op(n18687) );
  buf_1 U19631 ( .ip(n18785), .op(n18780) );
  mux2_1 U19632 ( .ip1(\ANSWER/mem[2][5][14] ), .ip2(\ANSWER/mem[3][5][14] ), 
        .s(n18780), .op(n18686) );
  mux2_1 U19633 ( .ip1(n18687), .ip2(n18686), .s(n4456), .op(n18691) );
  mux2_1 U19634 ( .ip1(\ANSWER/mem[4][5][14] ), .ip2(\ANSWER/mem[5][5][14] ), 
        .s(n18780), .op(n18689) );
  mux2_1 U19635 ( .ip1(\ANSWER/mem[6][5][14] ), .ip2(\ANSWER/mem[7][5][14] ), 
        .s(n18780), .op(n18688) );
  mux2_1 U19636 ( .ip1(n18689), .ip2(n18688), .s(n17605), .op(n18690) );
  mux2_1 U19637 ( .ip1(n18691), .ip2(n18690), .s(n18878), .op(n18693) );
  mux2_1 U19638 ( .ip1(\ANSWER/mem[8][5][14] ), .ip2(\ANSWER/mem[9][5][14] ), 
        .s(n18780), .op(n18692) );
  mux2_1 U19639 ( .ip1(n18693), .ip2(n18692), .s(n18910), .op(n18694) );
  nand2_1 U19640 ( .ip1(n18832), .ip2(n18694), .op(n18767) );
  mux2_1 U19641 ( .ip1(\ANSWER/mem[0][3][14] ), .ip2(\ANSWER/mem[1][3][14] ), 
        .s(n18785), .op(n18696) );
  mux2_1 U19642 ( .ip1(\ANSWER/mem[2][3][14] ), .ip2(\ANSWER/mem[3][3][14] ), 
        .s(n18785), .op(n18695) );
  mux2_1 U19643 ( .ip1(n18696), .ip2(n18695), .s(n18544), .op(n18700) );
  mux2_1 U19644 ( .ip1(\ANSWER/mem[4][3][14] ), .ip2(\ANSWER/mem[5][3][14] ), 
        .s(n18785), .op(n18698) );
  mux2_1 U19645 ( .ip1(\ANSWER/mem[6][3][14] ), .ip2(\ANSWER/mem[7][3][14] ), 
        .s(n18785), .op(n18697) );
  mux2_1 U19646 ( .ip1(n18698), .ip2(n18697), .s(n18354), .op(n18699) );
  mux2_1 U19647 ( .ip1(n18700), .ip2(n18699), .s(n18878), .op(n18702) );
  mux2_1 U19648 ( .ip1(\ANSWER/mem[8][3][14] ), .ip2(\ANSWER/mem[9][3][14] ), 
        .s(n18785), .op(n18701) );
  mux2_1 U19649 ( .ip1(n18702), .ip2(n18701), .s(n18910), .op(n18755) );
  mux2_1 U19650 ( .ip1(\ANSWER/mem[0][4][14] ), .ip2(\ANSWER/mem[1][4][14] ), 
        .s(n18785), .op(n18704) );
  mux2_1 U19651 ( .ip1(\ANSWER/mem[2][4][14] ), .ip2(\ANSWER/mem[3][4][14] ), 
        .s(n18785), .op(n18703) );
  mux2_1 U19652 ( .ip1(n18704), .ip2(n18703), .s(n17366), .op(n18708) );
  mux2_1 U19653 ( .ip1(\ANSWER/mem[4][4][14] ), .ip2(\ANSWER/mem[5][4][14] ), 
        .s(n18785), .op(n18706) );
  mux2_1 U19654 ( .ip1(\ANSWER/mem[6][4][14] ), .ip2(\ANSWER/mem[7][4][14] ), 
        .s(n18785), .op(n18705) );
  mux2_1 U19655 ( .ip1(n18706), .ip2(n18705), .s(n17990), .op(n18707) );
  mux2_1 U19656 ( .ip1(n18708), .ip2(n18707), .s(n18878), .op(n18710) );
  mux2_1 U19657 ( .ip1(\ANSWER/mem[8][4][14] ), .ip2(\ANSWER/mem[9][4][14] ), 
        .s(n18785), .op(n18709) );
  mux2_1 U19658 ( .ip1(n18710), .ip2(n18709), .s(n18910), .op(n18711) );
  and2_1 U19659 ( .ip1(n18843), .ip2(n18711), .op(n18754) );
  inv_1 U19660 ( .ip(n4362), .op(n18741) );
  mux2_1 U19661 ( .ip1(\ANSWER/mem[0][0][14] ), .ip2(\ANSWER/mem[1][0][14] ), 
        .s(n18741), .op(n18713) );
  mux2_1 U19662 ( .ip1(\ANSWER/mem[2][0][14] ), .ip2(\ANSWER/mem[3][0][14] ), 
        .s(n18741), .op(n18712) );
  mux2_1 U19663 ( .ip1(n18713), .ip2(n18712), .s(n17366), .op(n18717) );
  mux2_1 U19664 ( .ip1(\ANSWER/mem[4][0][14] ), .ip2(\ANSWER/mem[5][0][14] ), 
        .s(n18741), .op(n18715) );
  mux2_1 U19665 ( .ip1(\ANSWER/mem[6][0][14] ), .ip2(\ANSWER/mem[7][0][14] ), 
        .s(n18741), .op(n18714) );
  mux2_1 U19666 ( .ip1(n18715), .ip2(n18714), .s(n4456), .op(n18716) );
  mux2_1 U19667 ( .ip1(n18717), .ip2(n18716), .s(n18878), .op(n18719) );
  mux2_1 U19668 ( .ip1(\ANSWER/mem[8][0][14] ), .ip2(\ANSWER/mem[9][0][14] ), 
        .s(n18741), .op(n18718) );
  mux2_1 U19669 ( .ip1(n18719), .ip2(n18718), .s(n18910), .op(n18720) );
  nand2_1 U19670 ( .ip1(n18800), .ip2(n18720), .op(n18752) );
  mux2_1 U19671 ( .ip1(\ANSWER/mem[0][6][14] ), .ip2(\ANSWER/mem[1][6][14] ), 
        .s(n18780), .op(n18722) );
  mux2_1 U19672 ( .ip1(\ANSWER/mem[2][6][14] ), .ip2(\ANSWER/mem[3][6][14] ), 
        .s(n18780), .op(n18721) );
  mux2_1 U19673 ( .ip1(n18722), .ip2(n18721), .s(n18138), .op(n18726) );
  mux2_1 U19674 ( .ip1(\ANSWER/mem[4][6][14] ), .ip2(\ANSWER/mem[5][6][14] ), 
        .s(n18780), .op(n18724) );
  mux2_1 U19675 ( .ip1(\ANSWER/mem[6][6][14] ), .ip2(\ANSWER/mem[7][6][14] ), 
        .s(n18780), .op(n18723) );
  mux2_1 U19676 ( .ip1(n18724), .ip2(n18723), .s(n17581), .op(n18725) );
  mux2_1 U19677 ( .ip1(n18726), .ip2(n18725), .s(n18878), .op(n18728) );
  mux2_1 U19678 ( .ip1(\ANSWER/mem[8][6][14] ), .ip2(\ANSWER/mem[9][6][14] ), 
        .s(n18780), .op(n18727) );
  mux2_1 U19679 ( .ip1(n18728), .ip2(n18727), .s(n18910), .op(n18729) );
  nand2_1 U19680 ( .ip1(n18821), .ip2(n18729), .op(n18751) );
  mux2_1 U19681 ( .ip1(\ANSWER/mem[0][1][14] ), .ip2(\ANSWER/mem[1][1][14] ), 
        .s(n18741), .op(n18731) );
  mux2_1 U19682 ( .ip1(\ANSWER/mem[2][1][14] ), .ip2(\ANSWER/mem[3][1][14] ), 
        .s(n18741), .op(n18730) );
  mux2_1 U19683 ( .ip1(n18731), .ip2(n18730), .s(n18138), .op(n18735) );
  mux2_1 U19684 ( .ip1(\ANSWER/mem[4][1][14] ), .ip2(\ANSWER/mem[5][1][14] ), 
        .s(n18741), .op(n18733) );
  mux2_1 U19685 ( .ip1(\ANSWER/mem[6][1][14] ), .ip2(\ANSWER/mem[7][1][14] ), 
        .s(n18741), .op(n18732) );
  mux2_1 U19686 ( .ip1(n18733), .ip2(n18732), .s(n17794), .op(n18734) );
  mux2_1 U19687 ( .ip1(n18735), .ip2(n18734), .s(n18878), .op(n18737) );
  mux2_1 U19688 ( .ip1(\ANSWER/mem[8][1][14] ), .ip2(\ANSWER/mem[9][1][14] ), 
        .s(n18741), .op(n18736) );
  mux2_1 U19689 ( .ip1(n18737), .ip2(n18736), .s(n18910), .op(n18738) );
  nand2_1 U19690 ( .ip1(n18872), .ip2(n18738), .op(n18750) );
  mux2_1 U19691 ( .ip1(\ANSWER/mem[0][2][14] ), .ip2(\ANSWER/mem[1][2][14] ), 
        .s(n18741), .op(n18740) );
  mux2_1 U19692 ( .ip1(\ANSWER/mem[2][2][14] ), .ip2(\ANSWER/mem[3][2][14] ), 
        .s(n18741), .op(n18739) );
  mux2_1 U19693 ( .ip1(n18740), .ip2(n18739), .s(n17990), .op(n18745) );
  mux2_1 U19694 ( .ip1(\ANSWER/mem[4][2][14] ), .ip2(\ANSWER/mem[5][2][14] ), 
        .s(n18741), .op(n18743) );
  mux2_1 U19695 ( .ip1(\ANSWER/mem[6][2][14] ), .ip2(\ANSWER/mem[7][2][14] ), 
        .s(n18785), .op(n18742) );
  mux2_1 U19696 ( .ip1(n18743), .ip2(n18742), .s(n17605), .op(n18744) );
  mux2_1 U19697 ( .ip1(n18745), .ip2(n18744), .s(n18878), .op(n18747) );
  mux2_1 U19698 ( .ip1(\ANSWER/mem[8][2][14] ), .ip2(\ANSWER/mem[9][2][14] ), 
        .s(n18785), .op(n18746) );
  mux2_1 U19699 ( .ip1(n18747), .ip2(n18746), .s(n18910), .op(n18748) );
  nand2_1 U19700 ( .ip1(n18884), .ip2(n18748), .op(n18749) );
  nand4_1 U19701 ( .ip1(n18752), .ip2(n18751), .ip3(n18750), .ip4(n18749), 
        .op(n18753) );
  not_ab_or_c_or_d U19702 ( .ip1(n18854), .ip2(n18755), .ip3(n18754), .ip4(
        n18753), .op(n18766) );
  mux2_1 U19703 ( .ip1(\ANSWER/mem[0][7][14] ), .ip2(\ANSWER/mem[1][7][14] ), 
        .s(n18780), .op(n18757) );
  mux2_1 U19704 ( .ip1(\ANSWER/mem[2][7][14] ), .ip2(\ANSWER/mem[3][7][14] ), 
        .s(n18780), .op(n18756) );
  mux2_1 U19705 ( .ip1(n18757), .ip2(n18756), .s(n18901), .op(n18761) );
  mux2_1 U19706 ( .ip1(\ANSWER/mem[4][7][14] ), .ip2(\ANSWER/mem[5][7][14] ), 
        .s(n18780), .op(n18759) );
  mux2_1 U19707 ( .ip1(\ANSWER/mem[6][7][14] ), .ip2(\ANSWER/mem[7][7][14] ), 
        .s(n18780), .op(n18758) );
  mux2_1 U19708 ( .ip1(n18759), .ip2(n18758), .s(n18901), .op(n18760) );
  mux2_1 U19709 ( .ip1(n18761), .ip2(n18760), .s(n18878), .op(n18763) );
  mux2_1 U19710 ( .ip1(\ANSWER/mem[8][7][14] ), .ip2(\ANSWER/mem[9][7][14] ), 
        .s(n18785), .op(n18762) );
  mux2_1 U19711 ( .ip1(n18763), .ip2(n18762), .s(n18910), .op(n18764) );
  nand2_1 U19712 ( .ip1(n18865), .ip2(n18764), .op(n18765) );
  nand3_1 U19713 ( .ip1(n18767), .ip2(n18766), .ip3(n18765), .op(n18768) );
  nand2_1 U19714 ( .ip1(n18768), .ip2(n18888), .op(n18791) );
  mux2_1 U19715 ( .ip1(\ANSWER/mem[0][9][14] ), .ip2(\ANSWER/mem[1][9][14] ), 
        .s(n18785), .op(n18770) );
  mux2_1 U19716 ( .ip1(\ANSWER/mem[2][9][14] ), .ip2(\ANSWER/mem[3][9][14] ), 
        .s(n18785), .op(n18769) );
  mux2_1 U19717 ( .ip1(n18770), .ip2(n18769), .s(n18901), .op(n18774) );
  mux2_1 U19718 ( .ip1(\ANSWER/mem[4][9][14] ), .ip2(\ANSWER/mem[5][9][14] ), 
        .s(n18780), .op(n18772) );
  mux2_1 U19719 ( .ip1(\ANSWER/mem[6][9][14] ), .ip2(\ANSWER/mem[7][9][14] ), 
        .s(n18780), .op(n18771) );
  mux2_1 U19720 ( .ip1(n18772), .ip2(n18771), .s(n18901), .op(n18773) );
  mux2_1 U19721 ( .ip1(n18774), .ip2(n18773), .s(n18878), .op(n18776) );
  mux2_1 U19722 ( .ip1(\ANSWER/mem[8][9][14] ), .ip2(\ANSWER/mem[9][9][14] ), 
        .s(n18785), .op(n18775) );
  mux2_1 U19723 ( .ip1(n18776), .ip2(n18775), .s(n18910), .op(n18777) );
  nand2_1 U19724 ( .ip1(n18899), .ip2(n18777), .op(n18790) );
  mux2_1 U19725 ( .ip1(\ANSWER/mem[0][8][14] ), .ip2(\ANSWER/mem[1][8][14] ), 
        .s(n18785), .op(n18779) );
  mux2_1 U19726 ( .ip1(\ANSWER/mem[2][8][14] ), .ip2(\ANSWER/mem[3][8][14] ), 
        .s(n18785), .op(n18778) );
  mux2_1 U19727 ( .ip1(n18779), .ip2(n18778), .s(n18901), .op(n18784) );
  mux2_1 U19728 ( .ip1(\ANSWER/mem[4][8][14] ), .ip2(\ANSWER/mem[5][8][14] ), 
        .s(n18780), .op(n18782) );
  mux2_1 U19729 ( .ip1(\ANSWER/mem[6][8][14] ), .ip2(\ANSWER/mem[7][8][14] ), 
        .s(n18785), .op(n18781) );
  mux2_1 U19730 ( .ip1(n18782), .ip2(n18781), .s(n18354), .op(n18783) );
  mux2_1 U19731 ( .ip1(n18784), .ip2(n18783), .s(n18878), .op(n18787) );
  mux2_1 U19732 ( .ip1(\ANSWER/mem[8][8][14] ), .ip2(\ANSWER/mem[9][8][14] ), 
        .s(n18785), .op(n18786) );
  mux2_1 U19733 ( .ip1(n18787), .ip2(n18786), .s(n18910), .op(n18788) );
  nand2_1 U19734 ( .ip1(n18914), .ip2(n18788), .op(n18789) );
  nand3_1 U19735 ( .ip1(n18791), .ip2(n18790), .ip3(n18789), .op(\ANSWER/N473 ) );
  mux2_1 U19736 ( .ip1(\ANSWER/mem[0][0][15] ), .ip2(\ANSWER/mem[1][0][15] ), 
        .s(n18244), .op(n18793) );
  mux2_1 U19737 ( .ip1(\ANSWER/mem[2][0][15] ), .ip2(\ANSWER/mem[3][0][15] ), 
        .s(n18780), .op(n18792) );
  mux2_1 U19738 ( .ip1(n18793), .ip2(n18792), .s(n18435), .op(n18797) );
  mux2_1 U19739 ( .ip1(\ANSWER/mem[4][0][15] ), .ip2(\ANSWER/mem[5][0][15] ), 
        .s(n18741), .op(n18795) );
  mux2_1 U19740 ( .ip1(\ANSWER/mem[6][0][15] ), .ip2(\ANSWER/mem[7][0][15] ), 
        .s(n18616), .op(n18794) );
  mux2_1 U19741 ( .ip1(n18795), .ip2(n18794), .s(n18901), .op(n18796) );
  mux2_1 U19742 ( .ip1(n18797), .ip2(n18796), .s(n18826), .op(n18799) );
  mux2_1 U19743 ( .ip1(\ANSWER/mem[8][0][15] ), .ip2(\ANSWER/mem[9][0][15] ), 
        .s(n17387), .op(n18798) );
  mux2_1 U19744 ( .ip1(n18799), .ip2(n18798), .s(n18910), .op(n18801) );
  nand2_1 U19745 ( .ip1(n18801), .ip2(n18800), .op(n18887) );
  mux2_1 U19746 ( .ip1(\ANSWER/mem[0][1][15] ), .ip2(\ANSWER/mem[1][1][15] ), 
        .s(n17536), .op(n18803) );
  mux2_1 U19747 ( .ip1(\ANSWER/mem[2][1][15] ), .ip2(\ANSWER/mem[3][1][15] ), 
        .s(n17344), .op(n18802) );
  mux2_1 U19748 ( .ip1(n18803), .ip2(n18802), .s(n18901), .op(n18808) );
  mux2_1 U19749 ( .ip1(\ANSWER/mem[4][1][15] ), .ip2(\ANSWER/mem[5][1][15] ), 
        .s(n18351), .op(n18805) );
  mux2_1 U19750 ( .ip1(\ANSWER/mem[6][1][15] ), .ip2(\ANSWER/mem[7][1][15] ), 
        .s(n18616), .op(n18804) );
  mux2_1 U19751 ( .ip1(n18805), .ip2(n18804), .s(n15636), .op(n18807) );
  mux2_1 U19752 ( .ip1(n18808), .ip2(n18807), .s(n18806), .op(n18810) );
  mux2_1 U19753 ( .ip1(\ANSWER/mem[8][1][15] ), .ip2(\ANSWER/mem[9][1][15] ), 
        .s(n17884), .op(n18809) );
  mux2_1 U19754 ( .ip1(n18810), .ip2(n18809), .s(n18910), .op(n18873) );
  inv_1 U19755 ( .ip(n4362), .op(n18909) );
  buf_1 U19756 ( .ip(n18909), .op(n18900) );
  mux2_1 U19757 ( .ip1(\ANSWER/mem[0][6][15] ), .ip2(\ANSWER/mem[1][6][15] ), 
        .s(n18900), .op(n18812) );
  mux2_1 U19758 ( .ip1(\ANSWER/mem[2][6][15] ), .ip2(\ANSWER/mem[3][6][15] ), 
        .s(n18900), .op(n18811) );
  mux2_1 U19759 ( .ip1(n18812), .ip2(n18811), .s(n17794), .op(n18817) );
  mux2_1 U19760 ( .ip1(\ANSWER/mem[4][6][15] ), .ip2(\ANSWER/mem[5][6][15] ), 
        .s(n18900), .op(n18814) );
  mux2_1 U19761 ( .ip1(\ANSWER/mem[6][6][15] ), .ip2(\ANSWER/mem[7][6][15] ), 
        .s(n18900), .op(n18813) );
  mux2_1 U19762 ( .ip1(n18814), .ip2(n18813), .s(n18901), .op(n18816) );
  mux2_1 U19763 ( .ip1(n18817), .ip2(n18816), .s(n18815), .op(n18819) );
  mux2_1 U19764 ( .ip1(\ANSWER/mem[8][6][15] ), .ip2(\ANSWER/mem[9][6][15] ), 
        .s(n18900), .op(n18818) );
  mux2_1 U19765 ( .ip1(n18819), .ip2(n18818), .s(n18910), .op(n18820) );
  and2_1 U19766 ( .ip1(n18821), .ip2(n18820), .op(n18871) );
  mux2_1 U19767 ( .ip1(\ANSWER/mem[0][5][15] ), .ip2(\ANSWER/mem[1][5][15] ), 
        .s(n18909), .op(n18823) );
  mux2_1 U19768 ( .ip1(\ANSWER/mem[2][5][15] ), .ip2(\ANSWER/mem[3][5][15] ), 
        .s(n18900), .op(n18822) );
  mux2_1 U19769 ( .ip1(n18823), .ip2(n18822), .s(n18354), .op(n18828) );
  mux2_1 U19770 ( .ip1(\ANSWER/mem[4][5][15] ), .ip2(\ANSWER/mem[5][5][15] ), 
        .s(n18900), .op(n18825) );
  mux2_1 U19771 ( .ip1(\ANSWER/mem[6][5][15] ), .ip2(\ANSWER/mem[7][5][15] ), 
        .s(n18900), .op(n18824) );
  mux2_1 U19772 ( .ip1(n18825), .ip2(n18824), .s(n18138), .op(n18827) );
  mux2_1 U19773 ( .ip1(n18828), .ip2(n18827), .s(n18826), .op(n18830) );
  mux2_1 U19774 ( .ip1(\ANSWER/mem[8][5][15] ), .ip2(\ANSWER/mem[9][5][15] ), 
        .s(n18900), .op(n18829) );
  mux2_1 U19775 ( .ip1(n18830), .ip2(n18829), .s(n18910), .op(n18831) );
  nand2_1 U19776 ( .ip1(n18832), .ip2(n18831), .op(n18869) );
  mux2_1 U19777 ( .ip1(\ANSWER/mem[0][4][15] ), .ip2(\ANSWER/mem[1][4][15] ), 
        .s(n18909), .op(n18834) );
  mux2_1 U19778 ( .ip1(\ANSWER/mem[2][4][15] ), .ip2(\ANSWER/mem[3][4][15] ), 
        .s(n18909), .op(n18833) );
  mux2_1 U19779 ( .ip1(n18834), .ip2(n18833), .s(n17605), .op(n18839) );
  mux2_1 U19780 ( .ip1(\ANSWER/mem[4][4][15] ), .ip2(\ANSWER/mem[5][4][15] ), 
        .s(n18909), .op(n18836) );
  mux2_1 U19781 ( .ip1(\ANSWER/mem[6][4][15] ), .ip2(\ANSWER/mem[7][4][15] ), 
        .s(n18909), .op(n18835) );
  mux2_1 U19782 ( .ip1(n18836), .ip2(n18835), .s(n18330), .op(n18838) );
  mux2_1 U19783 ( .ip1(n18839), .ip2(n18838), .s(n18837), .op(n18841) );
  mux2_1 U19784 ( .ip1(\ANSWER/mem[8][4][15] ), .ip2(\ANSWER/mem[9][4][15] ), 
        .s(n18909), .op(n18840) );
  mux2_1 U19785 ( .ip1(n18841), .ip2(n18840), .s(n18910), .op(n18842) );
  nand2_1 U19786 ( .ip1(n18843), .ip2(n18842), .op(n18868) );
  mux2_1 U19787 ( .ip1(\ANSWER/mem[0][3][15] ), .ip2(\ANSWER/mem[1][3][15] ), 
        .s(n18909), .op(n18845) );
  mux2_1 U19788 ( .ip1(\ANSWER/mem[2][3][15] ), .ip2(\ANSWER/mem[3][3][15] ), 
        .s(n18909), .op(n18844) );
  mux2_1 U19789 ( .ip1(n18845), .ip2(n18844), .s(n18544), .op(n18850) );
  mux2_1 U19790 ( .ip1(\ANSWER/mem[4][3][15] ), .ip2(\ANSWER/mem[5][3][15] ), 
        .s(n18909), .op(n18847) );
  mux2_1 U19791 ( .ip1(\ANSWER/mem[6][3][15] ), .ip2(\ANSWER/mem[7][3][15] ), 
        .s(n18909), .op(n18846) );
  mux2_1 U19792 ( .ip1(n18847), .ip2(n18846), .s(n17605), .op(n18849) );
  mux2_1 U19793 ( .ip1(n18850), .ip2(n18849), .s(n18848), .op(n18852) );
  mux2_1 U19794 ( .ip1(\ANSWER/mem[8][3][15] ), .ip2(\ANSWER/mem[9][3][15] ), 
        .s(n18909), .op(n18851) );
  mux2_1 U19795 ( .ip1(n18852), .ip2(n18851), .s(n18910), .op(n18853) );
  nand2_1 U19796 ( .ip1(n18854), .ip2(n18853), .op(n18867) );
  mux2_1 U19797 ( .ip1(\ANSWER/mem[0][7][15] ), .ip2(\ANSWER/mem[1][7][15] ), 
        .s(n18900), .op(n18856) );
  mux2_1 U19798 ( .ip1(\ANSWER/mem[2][7][15] ), .ip2(\ANSWER/mem[3][7][15] ), 
        .s(n18900), .op(n18855) );
  mux2_1 U19799 ( .ip1(n18856), .ip2(n18855), .s(n18354), .op(n18861) );
  mux2_1 U19800 ( .ip1(\ANSWER/mem[4][7][15] ), .ip2(\ANSWER/mem[5][7][15] ), 
        .s(n18900), .op(n18858) );
  mux2_1 U19801 ( .ip1(\ANSWER/mem[6][7][15] ), .ip2(\ANSWER/mem[7][7][15] ), 
        .s(n18900), .op(n18857) );
  mux2_1 U19802 ( .ip1(n18858), .ip2(n18857), .s(n17605), .op(n18860) );
  mux2_1 U19803 ( .ip1(n18861), .ip2(n18860), .s(n18859), .op(n18863) );
  mux2_1 U19804 ( .ip1(\ANSWER/mem[8][7][15] ), .ip2(\ANSWER/mem[9][7][15] ), 
        .s(n18909), .op(n18862) );
  mux2_1 U19805 ( .ip1(n18863), .ip2(n18862), .s(n18910), .op(n18864) );
  nand2_1 U19806 ( .ip1(n18865), .ip2(n18864), .op(n18866) );
  nand4_1 U19807 ( .ip1(n18869), .ip2(n18868), .ip3(n18867), .ip4(n18866), 
        .op(n18870) );
  not_ab_or_c_or_d U19808 ( .ip1(n18873), .ip2(n18872), .ip3(n18871), .ip4(
        n18870), .op(n18886) );
  mux2_1 U19809 ( .ip1(\ANSWER/mem[0][2][15] ), .ip2(\ANSWER/mem[1][2][15] ), 
        .s(n18900), .op(n18875) );
  mux2_1 U19810 ( .ip1(\ANSWER/mem[2][2][15] ), .ip2(\ANSWER/mem[3][2][15] ), 
        .s(n18351), .op(n18874) );
  mux2_1 U19811 ( .ip1(n18875), .ip2(n18874), .s(n17990), .op(n18880) );
  mux2_1 U19812 ( .ip1(\ANSWER/mem[4][2][15] ), .ip2(\ANSWER/mem[5][2][15] ), 
        .s(n17344), .op(n18877) );
  mux2_1 U19813 ( .ip1(\ANSWER/mem[6][2][15] ), .ip2(\ANSWER/mem[7][2][15] ), 
        .s(n18909), .op(n18876) );
  mux2_1 U19814 ( .ip1(n18877), .ip2(n18876), .s(n18901), .op(n18879) );
  mux2_1 U19815 ( .ip1(n18880), .ip2(n18879), .s(n18878), .op(n18882) );
  mux2_1 U19816 ( .ip1(\ANSWER/mem[8][2][15] ), .ip2(\ANSWER/mem[9][2][15] ), 
        .s(n18909), .op(n18881) );
  mux2_1 U19817 ( .ip1(n18882), .ip2(n18881), .s(n18910), .op(n18883) );
  nand2_1 U19818 ( .ip1(n18884), .ip2(n18883), .op(n18885) );
  nand3_1 U19819 ( .ip1(n18887), .ip2(n18886), .ip3(n18885), .op(n18889) );
  nand2_1 U19820 ( .ip1(n18889), .ip2(n18888), .op(n18917) );
  mux2_1 U19821 ( .ip1(\ANSWER/mem[0][9][15] ), .ip2(\ANSWER/mem[1][9][15] ), 
        .s(n18909), .op(n18891) );
  mux2_1 U19822 ( .ip1(\ANSWER/mem[2][9][15] ), .ip2(\ANSWER/mem[3][9][15] ), 
        .s(n18900), .op(n18890) );
  mux2_1 U19823 ( .ip1(n18891), .ip2(n18890), .s(n18901), .op(n18895) );
  mux2_1 U19824 ( .ip1(\ANSWER/mem[4][9][15] ), .ip2(\ANSWER/mem[5][9][15] ), 
        .s(n18909), .op(n18893) );
  mux2_1 U19825 ( .ip1(\ANSWER/mem[6][9][15] ), .ip2(\ANSWER/mem[7][9][15] ), 
        .s(n18909), .op(n18892) );
  mux2_1 U19826 ( .ip1(n18893), .ip2(n18892), .s(n18901), .op(n18894) );
  mux2_1 U19827 ( .ip1(n18895), .ip2(n18894), .s(n18826), .op(n18897) );
  mux2_1 U19828 ( .ip1(\ANSWER/mem[8][9][15] ), .ip2(\ANSWER/mem[9][9][15] ), 
        .s(n18909), .op(n18896) );
  mux2_1 U19829 ( .ip1(n18897), .ip2(n18896), .s(n18910), .op(n18898) );
  nand2_1 U19830 ( .ip1(n18899), .ip2(n18898), .op(n18916) );
  mux2_1 U19831 ( .ip1(\ANSWER/mem[0][8][15] ), .ip2(\ANSWER/mem[1][8][15] ), 
        .s(n18900), .op(n18903) );
  mux2_1 U19832 ( .ip1(\ANSWER/mem[2][8][15] ), .ip2(\ANSWER/mem[3][8][15] ), 
        .s(n18900), .op(n18902) );
  mux2_1 U19833 ( .ip1(n18903), .ip2(n18902), .s(n18901), .op(n18908) );
  mux2_1 U19834 ( .ip1(\ANSWER/mem[4][8][15] ), .ip2(\ANSWER/mem[5][8][15] ), 
        .s(n18909), .op(n18905) );
  mux2_1 U19835 ( .ip1(\ANSWER/mem[6][8][15] ), .ip2(\ANSWER/mem[7][8][15] ), 
        .s(n18909), .op(n18904) );
  mux2_1 U19836 ( .ip1(n18905), .ip2(n18904), .s(n18354), .op(n18907) );
  mux2_1 U19837 ( .ip1(n18908), .ip2(n18907), .s(n18906), .op(n18912) );
  mux2_1 U19838 ( .ip1(\ANSWER/mem[8][8][15] ), .ip2(\ANSWER/mem[9][8][15] ), 
        .s(n18909), .op(n18911) );
  mux2_1 U19839 ( .ip1(n18912), .ip2(n18911), .s(n18910), .op(n18913) );
  nand2_1 U19840 ( .ip1(n18914), .ip2(n18913), .op(n18915) );
  nand3_1 U19841 ( .ip1(n18917), .ip2(n18916), .ip3(n18915), .op(\ANSWER/N472 ) );
endmodule

